/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2021_07", key_method = "rsa", key_block
NtAd9OZUX95s/dSCRNODTF9HgTWl+h4DTOkNb9Y3Ju8T8NsGbsgq1H0S/UY/ncbohmCQIVToM89N
haVItze+LvwnwYWnQsvE2QE3wSn2vHQBgtpF75htH3YYukKxaf+OWkteqlivrrYC67CenOg2L+F2
eDqr7yjC6pMxu4Ko0VI7zbm7JD6T/YF2iCb7EOvSaTDEVWZY68mzTG9bIUY0qZtjz6l6XTv3Quxt
aEodQdzA5VK7AI0QwWxXrcBvzCCG0Z+LBrGFhpzsF4KSwOHU+jRAu6uIF9Mtk7xllqFcpU95pCXa
f9sqX/ti/taMnyqGQUTUL6eUBij3vlT7VnLfBQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="QVR4QZEDqi0w5f9eyB33tNffNvNEl48tInsLa5sl0gI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 52624)
`pragma protect data_block
Mffvdu9pcmgNJk6bmxz8vUs8YelIvq9EC/+tHH8nrcTSrePtbPtRpnHjxkbVFNUdJyPFprcNO0Hq
+T4PTEYTYhjiWPS2NE7z69cGLXhAs8CuGS5Qjlwo7tmpZmBf5WD367r0DAmnXOWhoFIO25mudT1v
jSkfBk4PgjWoQciwRICfncxklmMLg//NJ4Uk9cWBvATOAlJ9EF5UlkiaghSh3fpn771cWD5VW44v
LnytlHL2Q3ali4+2nG5o2gMOBXnoye87hXnYrQMdOx/vXjqQZjsCRMfsBL6MgWzdCz8xKDvjbNKX
jieffDfuEZKIu9R9miDXPPzM5AIZ0E3QLEok1TEBwDuNaxDMu2FvmJMExV01umNQ+ieo+GFm63qn
+KJmqV1odkko5HUdWbctm/11fn3moyjxkx4JmcCYxvfNiy5No37xdvQfchpH1k9u+AVB4DwoynBJ
CxCBXxRwSE5D5ekJK25DEkdcsGjIjNshYnbeSWWmO9pjfwFdToXktq8rovtj2o2VFv2U/3FFSNEc
1bzIZlVXEj8N+vrTuRqxaGWuLi0JhEbB50tg3FU9j2EM9dPfiQSbrBaiHi76g9V7in25WMTS9NxB
kipk/j3amFr1ZFcAxrn4UTLDcJtU+CmCh1LHa6V7jjnEtszL3Nfs4UR3QaDBGtOP07qT98W0idb2
bqRlTUGI2SNtTzKXxePETRAFSIuWPtWUCvgcAnqkVDQPxidGVkTh0VQpA9oRzMQmyKYhLIkLCSn4
Dlo6klnJS0hoS+Smw/WSJL1/1Ha20GUaCWjxxOD6n0R8dVMn1cP3P51k5zps//RFfaFRf8RXTADY
Tpl53Ks9JXhK5QOX1Wu6TS5DKINHfLoIVP+yB6fEhNfEpN0wm9/6MdiyGUwHpzeu9MZYUbkyJrde
P7lVaMGpGW9BkwG1WwH5rADsJ+6G5JZ6JcmwZxzV6DQ1IJLU/E/FP90fHtQDAVcN22PrhekzNojk
xB2hRAmpONJjr885Nwi3sP6Mj83t/wS1jKW2QXgJ9ywSYDj31RYHQH1Zh3Z2fwT3vZWJz9p3XUcc
Wa7Tidh1BhtGOVNHdvtwtMLcLqTFBHpYiosBOZknoMCI/LSYYQ84ZkaRftJJAwP+rBNfywlLUT4S
lpR0G7bik6hfm5xAEHeqjW08AjFCQIXznZFs2JuSjSIZrRTy8TwRDy7l/mjWjOF710HybjwSfI2t
EeanViadPJ/Pzkd54CJtAnObz+FEU1r/kNzkC5D0l7s7X4x8JwbcJPa180X/w9BThtlOf+F0ZWcY
dbIDpJXoSBLFe4rFGoqse3fdiMstUI8ijKc5aVA8zyeL7TR2BXNgBFfEGsP3633t7LmcBa7xKJ4E
KKDxu53+UTC++k7hp6UMO1flF6DNaIW7SVmGcCPjIrVCcrNPnhbbExZfHRHZMyMVubtVLhr+Q4h8
Nn8TpAoYJbtVWkOKkdGEvp8LlZmWYxID+0CovPgyevAq9OAzGtuLwRhmfUuzi5HEM052lq5GmYce
XDhlnw3R2sV8IE4f4Y068GYujTCDEn0AjbJ+PwVm2ovWX9qgcWSRkMmVq7w3YNHDPZOnYR49bnjC
hnzv0WYECJ0ydVAtHNb4tXLJ6Rfg9Q1W0aZRzIFxC0f3a0q19wqQVx+RFlF1ExpFfFCnGmpwMHJT
RT1OZu/sX5XyPtLCZ6Vtiay0/hqW0dwPJ+QOdiaYyFoDe6jVu6ENzDz38JiuzfHPANRnzzRG6URq
WRzqPAgP1xpN5m/o5PbbFljumiqiaj0/YgsjL03bDv+sUo+xc6MHqfwIO8W2gMcfDcPDFTYU7HZ2
Ub1j4G2e0N4esAAQkEmMYnf8mPZdblk82y6A2uBvspmiFPjizcvg8i6f8UfUonMKBiwawszgr6tt
fz16eYnFdEqMJUfEcfwAVKqB/cFB354NkFbiwbGrmO/CAVP2O6tQt7Kbf2yFou1bFdLKTtxe/AFn
rRKK0Ho0R+cQdTrBajo+jh90ez4qm8SC8hhIiouiSDDXg+1KQgnwr6SdzgAD1LGA8M/issCgzK2s
NuB2AsyfLq5r3Ud1c4IhQg/VQwHCJkAM2II81NQzkaQYbL/IaCboSkHa3l1tQuHesl7SNpQBKgg1
Cg1jh19XeEdK6mxhmKUY6nYq1bvLWCBqd11B05MjqA/Ga4KP1wryN5SoELivqlGBWgCfGo6Xnuy3
MDaI8PHj4xCxeEHP7gsYH0CDHhPxsOWpfAH9Z3TxNMIISig8/0aXiAQ0x6dFN1+J91iBl/J5JxFi
eE7zY61FkpH8mZA7wYgonxujBNkydVc6GdreAaULHexIx0ZTjw58dn/Lvxyvy5IXVOGBEIuMEiwE
FuNu2I38F1WRv5OzsbgSQ0Rv+oiHwyti1+QL+ETe4/OmmsmjhCyte4+LQInPQsIzRCOkxGI7Po1M
FB9aAVNnHOFUVqBREkRj3Owto+hveJ5J3wv5fAEPvNeCeCeio6Ele/HufeTW42PUK5woDTUlKG+x
pUuM5TiYcUxdkSmyF2mE6IXfAuhY/jtBK93iycR5mqPaI9hO4uM/VNf2wypronx2JcJNUAlHIuod
fK+HCJKoGCQ1oqQs4GY2vJ5LQECx3Gx4BstZ5hPYiMXZvK9rOXgLkh5C0i/Mp95x7thhrxIwWPBg
GDbmNWAkTb88xhsFh4QHg36ZV/iLm/McoD4eKouP2dbW1k77UKJxSfQ4SwtECYeuBH9Sq3JJeA9U
qswI5gWj4vLPRCKG977989BziQXfWy8/eOE57AEkWCt8bk6Ebx9jA+ccQlhaUcSy4KoJ1DnljqFh
cp/3R85ehGnSYZweLGM0HJqddu16/cg5ITr6iMnqWeg5pBGalcM8O68w5kfyDCXGBO1LGLhhhUIg
u6PCe/53mggEzzsipfyysrIyoIpZ2Miu2rTZduKt9hUCLYk0HPG2ptr0YqektITrfm6kUWvVRsZJ
4FPkLEpeTororMa9wMrwAnwS91cshhMjBLdu1a119XYNf8oF1Pfm0FDkGbp0KQBqBj7nb+EQOQSA
sb4OtEipEbJ3oqbifFb9PcIVk37BCXxgOlJUuYt4yvlEUtXQiUewxGpVqUa0o2HUE2Vrt9beWzM2
v27tkkYCD+Zup0GNojONdb2B6l+YFFwpt53IBrAQZQsC6dz5C3SS1iklD8XOYToSV8o4av/FkYcz
vSQ7sylmYF8ua8fs5K4MfP6BlbFaC9Lh+2b+yt4axxqqH8ncVdOSlNCUEOSTEtEpo90VZXd0AxGk
oJl8QP1eUVw+Xd+et0MakzwIs/IgmujGthWX/tqmyAuACXJFE4BMlf6kk44ImcS18X/xMFhWASpt
PyMq3ALu5f/cZznCsjAJADsKJCuYFFjKGIdU3MeePkES65ZiA9E/BTvQ0Glg6f7SENFpCVZaKJCj
mZbBzEyvoCH8bMtm3Zz9/y7KcWY25Zh64nGiWo87QIC0lc2IlyMMqzSKti41z8VLiRL32sxdOfK0
jScrCR4GFfofwh0fLZwxet4Cz55slRHF83KwhAKiek+QPCgRzqr6ALzaV6hx95BWK3C80ixYz8Bt
fVTKg298OJWg01G0S4Fh+3Doa+z22DZ/DASrE8ry2K1wq/GZYKJG5hHRP0mEWzu6C3z8waev251g
DMB+b/KMxHzvxO+84bpG38tdoQH/9wXSjYHsyYaSLN8ZT/6iMvP8AEC+1B9WrpfY2wqw2uaqWT2r
SyKjmBHl6wiA7mCqshKmJuLY2m2Bl7T9q/7EC9oo50OUs8XsEg7kGmaeQrsPHCqOPHi4W2/Yto1s
JvmVsFPUddcth+sms1EOGE26VD0u3j2Y1FEuT8TcHBsiNEORXMZL3m1uHHdy6chkJE6Yiw7qGN3i
Qf7ZyDEmnY8kgB/glkSQ/9etaSolGP9/pzw+Luc43uzdKbp4uQHcVuSjMhcp1F+HV9Q4ZQTVUkfM
jahIwokquJkbwDnjDaf3QtXy9X3QZyhkapJ9doWWpXiCU4LJ7Cq4NYD1a1n8klrexYFsD9b4SQuL
JWS4wN0MydhqOKOIAjHyNQ1G0zRItx9zx46medd7kcJjYJvWKiCLAiciQGj4jQjnIXNDGPWI6msS
cL9AMtx6E6q59KG41TlPkppXhdbeAXVD7tN0BswNYLfmlovwTdugOuK5eDVmADkj/eRvfSUJex4J
1/hULsQcaWqmstkJX0NsiO/E/UKxd+Sw06GH5MbK9cCzV9f1f0DJ+2UUlhsokhRMI8adPtA7tuXh
r4w0Y5t/bPPGsImmr+6M8gqoHDFb68WDFaZduiS/13q+pvBTaCFYRfm6GoNUH8ynHoGisblwhEsx
s8gV9BpQz0CDfvBa/PRBhVGe7tMUK98H2Q2s5CTijlps7oKUeminJkKpAecO3e62CjDlI4ItnQrX
1UfpGJ2Wyfj6p2xv+2JBBzUZBEnLLQh3hZLsjSg8Z3gg60wTpnYAIcUskDlk67Gnlg4HLq+46g1A
1tCfkdI7wIO1v1bpiQgrWNbb8ChX//8R7cQbjoQnjtmM83dqWBPNTLqjkSm/dLOW87vSrHFcL0pa
6QfQ7+Owz1XlgX+4QxeQphf2reN0S+33BCShk/mhRmoWegvkHuqe/1lPqxbgyPrYvlBYzJ53m4f6
H21xSwHXL2kYCn+Ndcwj7OUAPRwRrYuSPGDIiKDoWE/srEz2Qol4HAzVb2PTtqMvmYQ6QTDHMXB7
0qovG2FaQQ/mFMWYNo6jO6l22X95Uhy7oA+Kbg7Y+06vCn1Bib7gzri6hnTkN7qI11piCZumvw5x
oHTDYS/2zHEi8t5OpJueduEbc2efMF+zdgJ7+07kYqxPOFAai83ZPXPkgLx1osp/2Zy3RrJ6mFew
mciaeWtlE3pi9rWAu6Mpr8oAWdfhrhTXBxsQYHVVsErX76AqhJmsYc1AOW8dhJd7sxJWBPikRtjG
iIZ1dBh8YlmgTWKoSss4abh00KJPp+ZV0bnfxolZAmG34cRTu21pz3lQcqea9KGXcJaIGQBsoJai
wpq0BP9yJod4CUH46aPnxXyQnXfFVe6GMWCdETrSoKbsCblEXpsuG4t8StSL/pAYkmdutQBOrjhr
kA1bik+vBuABtHaE97ZQf4bnLHzYlJaVe7xneKeAyN44S0hCKYhzMR7fhpM/N7ccnxWkudRaqnKz
5e0jNCpB5kF7jr7j2zBWp6iccB4ZYmidnjldKh/6LO7/70fDApgKGOfsP+CFiQ8ofoVabPo2hOZl
pndg4jl3RQk+DqcHuwfCdaAuAIIz/5jDVl3bmb0d8stKEnpClfPrqWAK1vQMBKra4mD3HFoYvJ+3
8FUeIqBTNw68clYEAEn7uuiBlehXyf129++85H4hIsxOqp6SyepdmeRrWupMm7tdLNeMzYO6Gsnw
A5Xb+cyDX4uoeaUypl1rwJSyYO8agIgONTCI/m5BTBvjEMERuQ+HJ0leuAegnRTvZ+rKIKVOzzlP
zPLl37PqXsrcXkw2oTvUWXJJIEF3YU/6pNfjiqS8UNTEhSYphk8f9eI4HJEmchWxI9MZMC5Nro5l
G8pPZyRbAPARemniimtVnkML4Q4h4Yn891p796pLva3QAlYUwu5KBsSUC6D/2/xxvW3vWCNwcu3M
PGV4r8g2fsv6zWupt/ai/dSNSBVwAxhTWQ/DI/JbNECbmTtvf1SvDs/uDHkIRDM1rZywICWGAMmj
q87ZCjH/rP6IaHnX28Hkbc1p83kSuuSUH8lr+fFnEef/92BoMpGv73LR20dHmF5Jyfc9QDUuokHG
q6BYi56d7S8ASl75yTCby67OVLziFrBdO8eFIBYnijKATtvFm6jW30F7rMng41xir0Z5L056NK0v
/wo4LItLcOm4F5LgcyF7e8ye9DJtCowhdrHZ/gfmcEOxQsJ5yKqdaEJyJA3sp5+P9LPkPcPFnsJf
FOrUGwOftBqEGtvWl7dNpomODJvX1SpUgEn5185jr6KuWCoDb8KLv3/YiBj/J8yCfe/d5tjS38qR
ZKp7/ub/9D6F2JzrmuxVgzE2pffKOGVsCWZxosoMPUrovHRzxbdYmIFaTPB5X0POJeV+aJtU53V9
5rw97XCPgl1YiISxSZ+XIwCesMKLqJ2c3VKDUUSVCBCqsQ0ghQwXrYPEX1lc2W063d/uvBbHUmPM
1rHk+C6cEQN0uiTcLz3ZXYeQVL3RvraAMhQF6h0CAqiuO4id4zBK2zr1GvP76yUhOWercI01D9d3
B+9fVt38zt5tE6FmNPRyumbZQgUBeIYunPNbm6BonnJAU6CTnOz4oVwZzbg++E1lCEg03vqhlexs
XccWaBQddlElt3nJtQlPTpe2zT73tiMLQEg5vNF8xkCB52GMRwfKqQr+LM46SMn2BjwYluVx7XSH
mqBbXsbluMCMSGm5P+XAPKfXGfQ+vSrZElj3UdDViaoNpGXfuCwnpGkZwRhD3suDy4yPcDjyolbC
X/bA3d+PtBos0xkrf1l36fZSnddBc8S9DAYqkqabxM34O7GT2J1ES7NgLD2c72Ynq5cxgLR5GPo0
yY5INt/EOT/LH+8vP4avrYNnV5AyB5IgKkhewiqwi1N4J14NhSsK330gPZQZIjkNIP+5EspTRj9K
J9zvj0ejQcshe4EeebepLKcuCpcgYukPkaTFtVAOI4rufe3KUPAxVfOHddILly8t4Nc7kqjjT8rm
slaUYJ+2HDWfgy07Syky/OlT/MUowTvDfomy7f33Z3UWBWe3yiBxZqcr4mnSzpIofzaP70yQNuWT
e6fs1eDN3hlzctnzQ8Ksx7Ko+vyZF+Tb0tPSUO7moeq1iQA5YBDJDyP+IBpyjNUFzEpJsN3dSTX5
K8pZgGTq1RJm996aV5ELy+2J4Ry2RRf0MdWpnNUzJJo8SObLr+sy8eaJZyzszalrswDkl7wE4tIh
gqAqn+WkvOW3XWDEBwUQmNy7TwgN9OrKywdwR7JNwT5qVSSTP4nXza8vr+DduPtOYyYYgvFjHAoE
K9by8YA6D+5515aNMb96I2VZqCWqQ+6sYO3qzTy8/9Rks/0ldh7m0iBhtqYpwCkuxqQ9kvjf6IK1
pZEBVIz7pwuK+4YqIKP06NgXtnPGI77t/tNF75LrghTs0fEqIYg3OgEQb9sXI8FUzF2JHhLyUiDw
hHOAimKm2ptPwoPsvJUb9RtamSHyjPGxdkppgmY3R/BQAWqPAAjQv09cY5Se1b+MvLuXqIkhtmNO
7Fo1sx6cmgQUldYnVgJZl7i8sDdkH5hehXrc/TByx6eGn2kTGNNiWRRcx5fS54UcIdZksjZePIRb
CWKGQ76q7V2yBR8fA776ffCOdkdQnMbWJguMOyZIG90uV01l/67m2Jnz36jnZmER2T6MYWam58JO
gIMo2JCSE1UHosnHTBmffPzH2q8b5PT5+woEM5rSMGo4xT3faP9wH8Rs5AK4GFPdbbY0Da7hZj3Z
NME87OX8CO04jtAGluFUIIQw/DGnc3vZ7UyzngaMMEfMTyGLHwlbBFLxtD+7Uc+rebH1OXsmeHsE
1ger2Tm5w3qTMfeaVwA7qNJKZtbNHGdH3uL9+Cc0MuC1zu/8TlpxKWGtyWCmKbtW/ICirc9V9LKD
3OPj/UTOgR4WA/kFjh2Pc1woWcU5qqCuBZB2SIYdtqilIfYiqUaywb1AWERve3PfXSgRnynGE4li
5qjNVksJXXkNNhGHEESWI633aPjnT6S58fm27IqE9/4rW9vhylx5v0kclaO/xGCLOtasqz1ruZDz
EURK6M/Qob3eabNEWkCTuRd81tnLnZEHwwQlb5GVBzbr5/Le7p0dneK8pSnKJgEv9pAb9WY5duyS
ekjAYc4aymQdA9SWZL3OhyG9NN8IIeLhHYXUNmRgYWg+ocWfpcp+xJtgo+Beekb9/2UqfWTKX0P8
1RUz/hKWz6a/PEOrWBwd3Aoqym0RnfVbrm5MNE4Ecfqw5aCTB0VV0jTl6RgiR5/0NczZg0TPsdXI
yLn/dcy0sBQcgp1OLTgSzOeG+2doh3NqI28ftlrmhM9652Bw7STOmPwLRM4hRc6GgqpSlytxD2qE
KkE8Rt5ovG+I1kiA/wgMWWzu5O+PjpePrD1nswFZNESSwH3rqzVDXutKHs9H6ij8fpIzh0pVnopT
yYDC6EvwtTK68xPLtjwjZfyyGsJm/gUkdNhZQbvwoLnFkF/EfovTvedWdS2lfo4Z19J6fx16txOu
5BgAi/NUWVRLXwsY0EbmQI+psj916uBk0RbZZQZV+dVSy/nzo6w7/kR75Y5ZLbivJRlYSRe+Agr1
zv7AIvXqkWUCvBY9DbV8LZmmLd4hFdJvJC/dRENtS4KG5U+1M+B5rysWbkFKFMTRmmbx9Ip1BUHV
vxmny6tJZr04r3c3PQkErdNamfG7fBLRfSPRC70Vsag2O3c/YgVIM0x40ZKYmB6WJ3vJCwBazF78
5sbF4oEamtiXLBb9td1MX+knkwsa4QqtfXEpHGGXn1eH4FE6Uu+2jitlGYVu7Le2Dkqa7buVoFFD
BB5yOeuTEUwiVMVsICLfUY19jaAbj6eR6IRrtYNa1glz6xyJg0cGphLoCf2UlgXM/wXuDOSCdWrj
zUVneM2GlZh8ytGAdrk1yYYINJpKHPGrTIqgR1iY8SBDM7tBlGqxQUhE9UxIMandlS8vsxCXupB5
qelCEkfxj1axVKrwQJOp7LsH2a0BifuiWhKoFKJDAPSihJ4qPudZ5rkfLVBCwxF12uGnOmocMKLq
rsgwkB2zlrpGCZ74i0w+V0CKS3eAfZ1/dYHBzJsPGs/DXfGCsrO/5K8wRnxKkl8XGRns7jM5zkl9
FS0HkX/KMJCRX90PIs0jqf/Nu8ieNfM9Ae2bZT3s05GeiKP+xOsupT20LTzSiHs3CGtmSKYIYsFK
LRMDmxwgnxbq5tlBsqZTG1j4BilVAXXiKvLhPLRgOVuAl+YEYCIiBPbM2NFXNsNkLzF6p9fCv3fd
7XwdvMJxpkbwdGhVszwINKPEW+Snswjo/92C1aIFVih6hwxrjLM9F2d8dDcTmEFiSxNOHhUDGlUW
lQUSsjlYNgB0CirrjIawnhlK8UNogOI7UHRz/jnkB1vCp0HD7KrSTBD+CLHpa8Jsh/SBxfpSCc11
2cFDMy/IKtg9cwW5uZoN4pjQRl0Q4IxO6kfp+fE3l1BlcZdyDRGFf/RLzAwTRunKYHV95ME1MheZ
Ty52qBt6T5tL86g5iOWiqURME9GUH46XDKmh4JWjKxbCZcAA2pGf0VAH32rG+NfTLy8Ee5j5JSf2
uTVLgHxR4WZEj52MKK2ARAr4SiaH7BwZGlPzl0ydSHUMWMBdmjFgex/WVaaU78/Noj7v46aZZ4DI
exDXW9Ol2WZ87uuuayshe65UGmbC5ZcICYWmvtvJbUKIvK2dIGsxWJRBOoxbaM3eJL4OfVhZV17e
6Cck7YuJEEYObnFA/l4GxT7HiEI6z8/BgpNluJx/fXt+Uhm5gOfLhh2hOjVeVEcjQZK8ptyj7MhQ
8c6PEq2i5BWf46xADtbVXeW5fos1Qs8JkELCkbP4TnaS53exrjyhlumKJOxW+HbnA0B0ZnHZ0IyO
3qYcgqbFBgDwGTFhqFPUxCcwrNUjVOUW1ZqokSqQAffqBEXya4id+ligokgqc18slkF5iqOd5aku
w6KwNVbjYJvSUDUJcV4G6SbX85AvfJ/9LwhmAutRqzDMMe4YAhn0ZdcYf2PXONJJEc/GlRmzxDN+
HvVPRxzho4UpJO8mKyHxWrdrnIoXIqDteDmCwhWSFagGuFpfxulXrDjb+TmHFyTuwmrPlrZ5VI3l
4gJO0Gd2GeJZ1E06ESLcUupxqB/p4sAcjHwmhiFw27ObB8Sg8mBoEkfLUNOUEtwN7rJQLsOxmHtc
g/Xhe6dzVQCOIv+WKwFtSb0znLWSWh2wFhMmTULI076eVZ4iqqCKax+8E/7HO6wpVto4LW5zGpXF
7CcGxiQ3ojeTIuGcucX/GjqX4TU6tectWd4RoJscTE4bAOHyzBaSiz2mpOIvNPEpuG6GDDv4I3in
ycVIz3uEfN5Z0F4upFcV7Tx8FnwgiT9pGRXI4wP8x2CTFRt+gq96aTvVFWLBCR91JqoG8txSmfJz
8fbLDLxaEJlg4OGXkUdTSfpLWxzVUWJWwp8CC+lw7cDKEvDZxVFS8axejyn4ynI6ysTacDCi/Cy3
Ij3oGrM7cFGBVqAoYqNHAP7m8zmg1XpQEPo1t1C+jK1vgtXj2HJbk2TKJipZkkRoAPbLzcuF0MHv
bufgqV1jP6ekQIiTbNJzeN7bmgwgybrHLY4XS1Bs8lyv8/CHFDkA8QFKnNYDBQkecdkZzjWcBHaz
ASLTWsh5gKsydPplMiM8LPcXfWEXS9/DCdHvi75JRaX8LnKVo84/K6uvARXoRgsNfWdpT6RnAqaC
f6bYsIBB2QTH4p1n079YdV247uRFEuaIZszgEpWFRJ+hmECEG8EDs9UcNOrObSXxW4ifkgChTpJm
d3TOaKnQ5ZaBqqns2Sq4tCFkCfjS6pijf2g3pEfqFe1727riiecKMHeG/YIm3JIuCxURhnEgnLh1
mTX2LGcNOg9DpASkCeC1/Z8ackp83ixmDRDOKkL0DFY8g2Wk9sgUO3CJvdNgUlrSZNLTZfpGY5so
lLh1Xbp+MDXqmVUzIkwv4O1m4+E+w3ah3WHRcIuVBAIRVbCPaXqYCQceCEVLIUQ4Tim2XPVyb6iL
UpkaquaIQR95cIgtxP5Sa0eJ/Ye8bN0X76zY9OTvwIHYhJcFvkQCVXRXhM7QzhCQNhpEWja81w8q
QU1MgyhTVFzwa2GsNv3zdJT2FO/zNyW36jGpeoDSJlt0e7iXEPQe2ZeboEZJRZlpb1QRzyk7RGqM
4mEvvItxOetPpzif8FwqL4gcOl+uT7o6BqNthCNrXUFuJQm2Sb3VtuR8jJorwuKs4pW23BJnfgxW
sbqKWGtdhOOCMV5PR7/bi840gVDIX2ipvZ6Xxhhb5DMtJj0DTtI8m+01hygFx6DzRhpXEb8rbYt+
sSG0BAmpl0+rxpQr+u13mP7bLBNZ/q7sndiwX8QhS8CFKkMFZ/AcbtxzrOfj6/vi2TXI8UJ0F62B
EQ2cFldVCl2tKP0uTE8+5OM5NqI0Dvp4IAlouPLbZs13rrZe6GxEx32BnsLa8euygIVpVuZHdYa+
fHnXUxT26t1CsRsVG1AJPWOLIy10jHxwO5B97baXu46pUXFdenUty65U2tTKke9stZ6d0S8VoQoq
F9rZ8yQkxl61zwFUf9yseolWSzTiH5POBOzwS4m25bl2muHXZFYXqoxU8gmweMMuK8BJqpy1o7mH
dmwVtQoiTI/IsXwMcOFiUU1Q7PyeZN5CGSQVTLWxfolCDLT91DMtBKJisNk5HpvxsDvpR4eOXXF0
M8pSgySJd4FZuaoAzEK3OPx66Ckcyw2U5W0POQHTvj8RbgGgkO0stqe+bdP3MUvw8hA3fSiuZhOs
4JdweGh2vtBcqafFd+KpbnE3eyPPJV9Q7IxlDERR0HQCOz7UxtO8oaVY98Zurq/n/kba3DQrLnpo
3ZhWbkTvoDSpC56iPlCDvk724OR0nfshv+8lPlwIrsm6yxFNOWaNUJHy2DmpPbsTi6M73cXKYBoP
RSFAvTaWOdFMsg4qjCFweVDkaT5UXzphqgnLQeOZA5uedSo4hYOlVGdHerNDxj1yABZVNwEWGaKa
+Jk/MmSSDw8FsByM/1TZZdrLE9AUw2Bg4Ffy+jVikJvE4DC9zSGTMahn2LHBHDyqNyTS3UlIDHTs
tMwI4tnj+uiJBQsby42y0kS7LlAbuY7wqbEoWvo0ixmU6GOum/VOsBdndAu4xRm7e+OEmtz27Q1I
Af3/CmK9OGnaZHLSR/4+LIevNGcfBMfzF3lGngkK4+dbaUB+pgqefi/jB979yrj2Q3Mz1wz2nSZ+
VKiqcNZny99JaaeENF74jVXjsdb9qFPIBidiK27VgJdFeG0v9KuMdOz94mClv4Cw3MCQ3NDlVjC+
VGvGWrOhL7PtLq9jWIYt69k/CAtx1HJ2H0o3VUxTacWxau75utMFI9VTbXHK9d4qCcVqmydsw51t
AXXOwLbz/Z2kOhWZMLZWRbKscbLnj6cS7jUammfh+YZhWIXQd0p4xMuWhML7rcBalEKjdrr4RAMu
st4GK0NtopSjWwTSI9xPs691owaSDnOR+SftkP5YsstDq63QGBz5xIHMjV24MR7Ylh1c7T73rcdb
rEu1DYIxqigaKkeKrpJEkZW4nGT5gBrdSYVa0+ZztpIkV1lvE49tcFvA1hWSqnGc2aBVBeeYvR6k
Rg7ox4d1ZwVdqm6zSBtAHlWXKpM/A43IFotmdsuqAbDsqsyZSKhhSKRshVGpx/ZQqWl85121+3yh
XwRNt1gFmAqajdnSKBp16EuTOG/9LMiIj0ZNjjRn957m0t8Pm90wDcdXTNvl/A+8BTRgBIAnAck5
rnQSXGuk/4UuYkDNUJN/DJm4kDOly+B2mFmU4d/XTCFJ4Y4vzgDRE4vC9XR2hMCs/L3k8ZLzbDKC
gpruUgHG3w4LaGG0aFaA0ao0zsdW3bj0TYJc+wAjLvXAtg4NmAOkMgbgzpXMPlIISmuvC1SVJa2M
4ftMgWwVKZRleCKa33T2/nURFmYwnjPNMd2Cgp4z91PGXzcmmCEo++NEhMKU0Doqrd35XyyNr2Hm
rbRRTf3FE4ci7AWCmDDQLsrN0adlt6IpToG31V56njWWNAHT/vMJuJjdFkX6BzqAOLk2aND/LQHU
C/GhEh+FFtzw2sztbd0/9kYWHXphmW65A8fxKkw66aPLWQLr86cHNgUVfnSWuholAWa2Ui5Zkwbf
6QEoK5WuP9zxRgb0S6s7nNw9cyVAEY9NbLk/iFpz76H0V0Oqq4vj5Re1eAT+o4xT+pG5SzJkbnDr
6TC4cffZXj6ReZ+28zOK1vbq6/zwkgnKMXe5Maf+75LSlM3BF3HN01FijxJlIHDqV1H6vnP8F0Nf
RiADPimX9FtEMU68kCx/FdMIL791HX4rqjRZ6Zc9mlDuYSX70zCPG+RaVoAkoMWeLZ1D80JVXWVO
Ok7W7K6VEqlDj44cU7nrsTsRP/b91+PGjfS5txkM4qLIfq0VnKlS5Vd0BpkMNzmHOutDUIW76zKP
k3bAXr+m8Mp8Q5zBdbxi4+Uozkp9XztpuqhjKwHrPF43IJyhpBadz7RWzygHBAwtnxzrZBd7Y40N
eh7J3t5lW0ovIrnvIWnGb/5lxbK3ZeBjMyTcPZEgMD+j2YTFiNoK61/FOWSIzERX3/RojIa1V5QM
frcFsAs+Z8O1Xm0h+0h9JP4nN6zyqWU4tbl+VKpHZy7DdWq0yjywXwoRqeIW2CvtXMD0vwn76zlp
tqVPyxnyHBduCLKKuXk8zepCUiKFtzzmvt75sQ7r5Yz0ZQ45GL53egbbMG2Nypi4mmo0bUuMaoAd
c6AVPr7oU44m1eId23Mb7RU0lzPeqrxW4HgNaLy7kI8WE7OXA9z5x+da+pqixdCNe5ugFL2UuG2i
Fts3HtKUX6hnU9UbYhqEq2lKB7kL4k0EnOoto/3LlCNe8YKkCYBtKb1uzpXntKsv2NuFs5pApGBP
sBWaxylxy8xq9ANOFPf670VOqcfEJyNGCBTe2DSAe+b8vhMbwnrxxPZEhLp9c4VW00daQh0vWTNP
9YhAiTBhLeRx8SPx9Apfx2aL37xd1ixduD9sD05R91/sOOSz4nttyIWi8pnWsR2coi97u2sXktvL
ezY+rlO6lFrDYUXujjwJ1IkNtUlgZ/TFb1E11LSVu3+b4TclfnwAc2GQ/5fIistkmDzZbjvrmFZj
976+X1B5X1uyReKOM68TzmHiWY25e8gFrAlw1T//1487qKgeHfc3cLU16Xo11VSzZctSR9/YIk6D
ROYDnbSx0XsNoQjQRvBy2thvBfQt8OLF30fYsXLsyj6fjyc2hZXhZcZKjN0DdTeWlyrr9j3p6FBM
4UQCm8j628wwxGsPzTQW5AHVU4fCCrbd7pOnPuJldORKCIxqsLPO5fENh2vJVwbdD0/WYvsTnnxD
ofhiE0KdwxjZp4UfkhuB3njRWpVWKrgR7Mk2vIpBnyowlaiaJ+Hzvx8CMc4qPJsNe74vn+3KkOha
miM2Bt4vUOBE/hl4Pby4CbiE4mm/Tqmp3ffXDuLOtVUuTKzEzMW2MAvuGOc6Qr7wQNF3zc/dK39P
2cpekY2d7Y0pwPMsumxQLoP9ca/AKXvazf8ia0sI+1NOdnysmveM3mTit4SzbLDMJGsApqRblUgo
VoU1n4UTT9HP7wgMayMt9PkVKU6TksqxJyCE2oelGHbKK1Z3RC9axA2PZ68n+c1RCFtXI6Q/KJb3
QuBa867B2xlaV7gII8IESWp4+bDrIHP4ndRmr3gfOuzgGcVFzKbQtFcaAe7FkcZYBon4BegUn/uE
Fsn4ZjPkIiZVovq6emF5XFy8nyW6CBq8FsV4A0Zc2PVBI3eQHtLgLJU2UEmJYOVeVeyit0lW/+LY
zJrp0oJymYgTnWuMAELz3ZoOdAxN8GIdQTFIto5hlN27bnL2FqRD/5dH1Nn/oF0DKG2/laFMZlvs
prksho/yWwtJZxR4tdVJwUUus3BGru7C0e7pXacOe7Bfq0CV82puqtyfknzcjMCpkKcfPSXw+rEx
XlvXxvm9tNoE2ZQWjT5eo+w51eVwZiKQt8zVWWbN6oq4PtQEflsXCRp7brIVSIEN7B4MkdAnchVH
KhIXXGQwjtSB+reQEIhW8zzi2y9kTyuvYM1hAqUw7LA7Wnkkmg/sj2lBB+6qAZ3d50P1PDMukaIb
D5Z67MQ3ujRG2UlzNe3ShOlkmh7+W+HhkTH1rR4mt9HzKZnYh0xXxaG9pqEAQdNFb4Ld3OS+YpZJ
4+npIZlB4dOz+JFZ67FUifvo9EdZ7alL0VlGztI5pfm3quIZUEncm3A4ri4Osk15NFJyAzq6+oOn
6c8w66dI6afJbh3qImRzPyghs2tgeSe/SitdWu7b3DPTS7o8oa89b+Z0S+A3tsEmoD+VX46A1Ysi
y+1dtXovAp4OwkfMTtd0kXPXrrzCtXVdn5n21Do3QlGb4DWvs05tUhj4dlRieSmRNsg7AZuld/dr
PinZbV1tPn2lG81/YbN+t/tUGwVQY/cCNU9qNIkqpdRAJQoZ/apiKC8DGt/BXCkZ3KMWcAJL0MY+
wl1lG9GHdcBY5WKRC/F+MrCnrE12flIKB5dRUWbZlFqBlX1v4gw//VKDyL414dkYOFhNwJNI45UK
lMLO2S7z7UhshWgX4mRBMksltwSo7CLhENsXd300BnrN8ds91CTg35VHDdPaRyMtbr0OP3rqKcJ1
CUtVBh8MSk+eTSvHBUQjfD1dsQeTYYx5tM9oivh7Ty/sVO4I4DLzll/LzUM/Q7dA42GSGap/6mow
GPLzqD3qQlA3CaqShKvFYlEoXvTRhOOGmdIQDkJbrx6axcCZRlT2kqKQ551b729Ixx9DZbxMrqF9
zN44bQ2ZIZhq/nhhEJzMUXLWKGYyUxTsaFiHMhnXWUPwwofTLF0nXqI/fnqBSOmEihTxa3arm5yC
Ph5dnz1pGozg8+fhW6tbDKZqI3vD34EbUCNadMF2qG3zIMoFUL1h/1maj/HtH4dbOPpaBqIlTS8S
zAT3YeQWCIU1g5JGZYse8GJoHxhc14MyNrPza4d5oVkJ6IcEz/TE1wrOYbW013p1eq1WkfUsnoi2
thnYPitnT9K1OjxJnPZ64ouCmJBZwxpKYUDiSqdGAHsTFslOqcCFC6R7ma618DugLbxYND3/6SRp
RlSImi5vi6/jJ7CmfIDxvVszqoJ59grJ/L6fz9IE/XvPamHePWdEuVHUuj31hFhFpl2da2dH+HQ2
voRB9axqnanhcWlJv8/nx+wjbbIeY8YyhKL/Q0uZgUBvhNzxC1pYFHaabRMcexlelPP4uISWfYhX
puJpmmOqQBEYdRZk1Fng17oHnMdPWzchQO1RojilmL2lx8XhsY/XW6GBJsqX6/a8tpVsen0E0gsy
WfHZYiDdP+v/rR5pD/xObWbJ1dqmDdhWDvkXoKG2iVQC0rAS4V/4HQ0okNAHExchuTH9inXm60K5
xToxqQ/uM5Ei9A4vCuIvW4R6kRqbOoqkOgGaVc7xu7p6v/i/cjCk8MIzU7C+OBv2K2AJZJvVY6Ld
122W5r1E6IgkCvY8G4Gye60Wt5aONqbGTjmgB0YiKgpJ19uc49Ha0NrvlxB9xfzmE558TqbJkkgy
/lb+ecruvv1TtzvVVDCn9APVxSJiZH5ea7i3VOc2iYazVUm/tIR23rZQx7ybx8XOQdyqa39QMbwR
3Xsm1cSobmOq3WEqho3uyadqufgsgHd7TwEbs4tEmpEI1aIEwJyZHXnERh/XVIuitgml6wBAeD18
lYfcdaWHkjlzxEkYika9sF+ixEcFtO/i0qA9qetbnbcGIKy+JcNCMugNPJjqYzvis9LtIH55pkBG
gZ0ajGjMUjaBh1pTQoMTEB0K+AOjiO9XNfs1rBr1x3LaaUc1/rCWBF85nXHhiOZ4Td6TESrYBV0g
YRXSOKCYEVNSnzqZ/vOshMoNXEh0ZKhBuKRWzizHEPogAxI01mYjgl+OHmHLgKIv3jZIAfFE+nsC
PGyPfvXdJ8Agg+HTXr0YyMua/VKih79p6AQAV7XfdyzmVTgF9XrhH8sty6foBlp1H8D7yXJMN+P1
uDZ/rum9hCLRtLCaPOxDR2VAyfkLK4qyHl56znDxRVPVVC1yKyMOwYLBC77G7jCgjuWtiPBEaAi4
bAbWbiqN6vVsvTMnU8ALpx+1FDpnSrHFhKW0mw6hmm+QW84Ggsh+yn78mapK+nCSW/Qz0K6ghnpo
00zctOW9OjOng9lZDYFsc+KR/tqipIGYC7mfHZaQdzaTCtfdW8DEQidFZjFh1xA19FNPkQyt0UHE
U5Fh0jUVI+TmZRZLVWOse/awjYLFJyijgJxJs5/3vU2UStNA0lZQglaRR9gyPkieAGSTkDUkvCPc
kh6jsa4qQ/C57TqUFXMd8jh8lxICD77Qx6aahrNYTVyiMAqb6B34S1Ya25UrZaMcqKYBKZK3VKe5
ZfzCYS+ty9tcvBxcO58Q7dToqf2/4l7SDoIjZML8BoIvA92kRJvYETw/3496rPrCnajJjaT26pXd
Qyk44FdGK9mMzmM+z9wB/cTMcljiqzMI5Lc19ufbNR5Lvy2663WNLSXJ2RQcs1ZNQVG9rvVmvyZP
YoWt7f1Ke/VbPgPmMvtz2B3yUBah8i1ZuWfa0mT2Ajq7CtoxSrq61bw4RyXR5GWXN3sIrNPeaJg9
Uh5wbNQr2uFSQBc8sl7XmS6KVFmn8A612/WeD07cDdovNuz3mQ+WEpWkd1MKfcRpLYUJDhV5ioFa
XKPmjP86sJfKHEFCu4fcuYVemB0RalFd00imar3in2wClhw218HuYDNJLs2Hw59IXkHgs+hA53FN
/zJ8kZNPiKyfviwlOn/ZB8zdbCUvvynChVm0KijE8Y+gddTYh4GGGLIbjprgRn8T16mdJLPOZXPb
d4kTICVnKJ6BmICEANSQxYeCkmvA6Ex+SWeMhEqIYWUrWH+SEKGiH9uigoutIR7BjBlneggD4yxY
Z7pW+5hkkD8L7YFlHtflfLL4LOEWxc4lJl8DALf+tGsMROUfyXSWum6YSTWULi4iwhPGtZ4b4jy+
dYmI5jK8WuAalsK4azBnoS4DpD9NgE5ZWSCKBMUo0WpEeLTgWqDBMWlci0yx/kfuMJAVz+3Ik/yX
1yYIJpg+AwK0jleY5XAaRnFNrX4dZ1NITwwgBo2fliuKNbtb+/MWXcaIZFV4dAdGo85sj8gaf1wH
ZwhO42k0QoQj6WDr+oSSm2Rs28EOy5tCyk25EI0LPAiwwrAaJrA22WszqEd9xJ0LN7pP+DbtWkEt
C8LjNf0eddl4/3ciPNVgcU4jyC2AO7qNPRJI9RP+YoS9NkCL97AImD+06i24kHwY4jTUW4TwebNI
gLIzfMPbxdOdi8Oz85CQcohGg5aAFQBJM5bV9Gaka0hYgDfpdpBaOrDoDzkzsop8038SZB+xoFb5
wtlyZdDs3XG5Lfi2MC2qNgkYp9x4Hkj02O/q3YwpDkvSLW4M9mbCCz6ifGSJusXsfKa/brNCmpJk
xF4m+lmbC0hXZuZCXPn6fWSr65K4qYQDJk/aqkkrx6LGMUBfa2J6CMpclevUimb0QFcqrLq5Qtx+
94GCK4fmk3f7ixuyEilMWlMAZWUxalJU64kEAAu/xlT0yo3rlH5GDp9MeZ8iv/Bz2hcGgPTzUcnQ
HUjVZVDeMUwMqQpUU/Wd8fjZgNSvD/y/qxByeoJPBXrCO2L+m2IOYu4GHWWGcCxynThojWAZGjD/
KbVU6FHCl28J67yWwLZ+cOs33uib/TvkK9rxF0KVpUvdXfMKROIJOpZ+SuLsQ9Njwaxi3vTF+im9
hHPZDatfrQ2mJzuDQDzWhiPbCWEDxviaCYltts3zf35f39Rz97/IBkzQQYY8X2pN0xVzWdlPp/Qz
vkfK7keMNOOnDL93GDxlhpW4TQpGOAxXtksKqaNGSCuxiQoLHmzC683c0h5UGFjWRM5mj+ohA3YK
NBzabrJuCsV01VwTE+HQ+OKNoNU2jUWewhtQN9tbnf+ppQay7f3NiP9CpXv36kfOLdFvAQyhIA7p
Z9jKpoDaBH+Mt995MHhafC6QeNKOFqGhPcSss7SZFBdjSdiMdUcXDYoMMKhZF7pr5oFKKaduqnzZ
Thl7LZGi9vT1UU2w4lPYY9rzyVLIGjFVSK1vRfMWiCbtlAQRiuTMQDNeeWYCI7d+xnsLPPxvpy9a
8Ca6A9qWfI5+CFp2K34edHA4gLhi4lmjSPw3iHl3E6V9K7/4PXpusCXXXN+1KhYTkQ8kA7SZ06mz
WM0F5iBpebTBQxsIUs/i5Gjs/ltpAQUY5t5GUTmapMUYGRgk6q+HCQW9kzh+DtTNp9LKA9L4iHuf
/OBRQNttDdMbh9cqtWY+glFQv77x+AjzfRW3R14W/xXat3a8FofM2LXr59rgVLXVneOYPMNPw2hG
c+KBmuB7yilIKyjPEdciwK6dstEWFq0jWC8s+xT2Kb8Tegb6BiSm43mMyV11MlsUEYR/Q5mvVHqZ
Qc4uxTWzaVgB3rU+9U64Sj2YoN0+ZuCI//7a3aNtY1elx4sjASKb8AR8jZ19UJuLZgnwAxDWLuWe
P16FKpK0EBhnh9yWhmlBjM+93ynX8KRPl5AxHinCBCaxSqUZqRJhqH3y4bplh0IHbSrLMaugQUMX
2GwDTAGpqVeMUHnhhAhmH94cBYoOHNSVy7ZSsL78kz+eOkJ6I454ZD6ivp3OLkw5s6E+O7GMVbZW
n+yhM3wRJZxlnmC9oXfAyrFAOFaYanjhSt5Otf83LS1nsQF8SVPp4n1eV95j3UhLeTphA77mA0Tg
Rj/JHiGnJBa7QjVT83r7hmQ5VTpZ3qu+bAa3/ZR9c3jdcJlzezrOSamXMGI+JjmLwq4xBHUT3Rai
WjVquA8G454JgozawvEDxfBoyh5CX2D0nkvS56/ZufEWW24Qmhssgc1Xb1Q2LXW1VQtK+Y9iedz9
1UJGoG9Edp8xAvZynLxDYn0JrAxHgbWgKlArndrxrFca/9qQ5Xpelik7j3vmkvF3HGIDLym7cL2E
ja0r8ZsBLy7oIPFdFvDX78XO88K4TxZ06Oo8eSU9H19PsUsnx+LNjVDdEe4To3Xp82HfW6a1Ndw3
LjCEgFaanbKIwWOKreHbzyk10N8VoSSbHlFjyVSKu+4bZNkBdJF14+/DqNVyOdYwWsnjFaR/P/l+
2HdYMx0RF8udnphsssO9VnYBE8UsNRAV+42KunZ/b313QsH2vTtgeQGcdzpDYRORFmAJvPc5qFU6
aBGtzlyCiYo/LfV5J2mMweY5OS0DlPqHKhGS43s25qCYDy84yEd3FNtLwHnXcX5zKyLv8aAlcebl
LIx0Gxw4xneTL1cs9ZmmLKE3DLmtZb/Al2MLo3AKbo/sxDf9xD5mgXUgvH7xsdNzrS+kdjJ9I50h
ptQIK/ORgoVXQ2hfST7XX3l7yG5X3mP/QmAXQpLKZh3AhkLn2FrcU1FPzcP4YTG9EAwOKTSk0V88
pCji1QnPYEHpLQlohhFfFJ/RSanlDnuhVRP6RTjjWTT8HCrXI9oq84xOYHYfgyYaxWDODiWaJqbE
9sIikoyxAl0dotHMDSBlIMJfLOQUvkPkn4R7FDKmUfWymL5mhTNcF6NbJmozXRelWEer6lfhk/Zn
I+bAjKLbRj9/2uQsmUuovOMxoq9xqklneXO3jynTjLVVb6R4s/0/+ViAuAF2n/MZXPLbbku87fnI
jnXtBLa0fnqoX/Phh6aHG+VoZeZLf29KI6bqCYeOTGv9jAMdiSBw1zo0PGw6Sfla20NQDIWBbLtI
JS3Yp33Q5KldLRT7R+lVMS6GAeF4dEIZ+jyWcT15dwXvf2KHDmQ2gWAvOQ6SfWIH9KoV7p2ksPVZ
xEkUq68ieboIOonE9s9nvj+KbZVUBlD2HRqAINu7MXzBnQEwZYhWUbnMWdGZBllbC0qk2f3Qm/eN
KXsWS04QQqaV+bz5tEeQ3XclYuZuXecWSrpN8Eg7OtabjKfrJbKmly/dNcoXtiDszPYTyi/O6ler
JyObzHGkj49ciqWoyo7AOckPytzRbazrtpF+NlLELBY/NlHN0YbzugPU31eOz3md6lwbDFHg4X+A
bzi3LbjF/b8En0vBcNQEjCnZ/xxSuQrKb7uu+meTF1HKvM+hF67wjYdKqKo9bv+3k5DM1sn7PEd3
K273rNuZuxuXSr/Y8xylarOqrNso3KKYxiL3+Q3AzOZV41TR6ev9O7G0sUhsI211L6FiICIS/wnK
kNtFUKxn8irKn5aV8L2VcIfuPGyzLMPcOh6i0O084AYZynYUczegB3JsZAvhT6wJUUU2cEnE+ZFx
aiJUOF3RfYPwmLzEpG9A8D3/qMfI3s3QpWNXO6W8ddn3CqVy6q2abd01ydhin/j1g1qFqYm8xVfa
hYpbBkj/rQGxgiVyIUbUxRUXwSiIbmMjDdnMAWyKbXbEJdP5S4pDa746TgMwVK474ZOayN0qTae5
0gywYpXedVIWPoYMu/ueKXTTlUGei9nAG/VNMjSbyyO5Qq0Z8GO3qJFCiJLK3tPrbIo7qcGY2N5D
V3N71NsUVLQQ8b2bRWpu9yuodKNMNejlkV/kIvToJmJryzqMVIf0rmMTI7LpFPr/9Bet3RmiCTKb
GKQO/YoW5oKvQJZdg8GjN+7weKz2bYL9kSt9FZGDvU/SJC7y09VBVHS7EEYm0eMOOiy9k9B6hdqX
x3qrSxR/3dksBLIb8XoJTQWc8sKWYvGbirREuFTbubi56i/ZK9tQ0u1g6aodajQF72OPB8UjgG3P
BkKgC18TEfn+NvXS9Kssdq9LnCQfkrZFmmmqThVU75C2msTs+oFRSERRYVOALBrjFBGWTVlFl8Vv
xR3Mi5oAKoQd7NQ6MIL6nFLaGnmXkl6LhiXOoUBVBCICBlTqh6nw33+4ITVTvEQfnMPCuX36ece9
HviWYfUe4ITWsUKSbQIn6LZPgGnU+s3WO+rEEZBJvcf6FS9DP11GFhSFzdAW7GFsJAMen1+B3oY2
jbUQ6XlszRlxGQw1EnzgUONn17lk5O0y1incb+LLj9erWDenzgVsUQ9p4GWjt0GP1FHuPlSgRVIi
MZDBh1fU7hWirmXhFZU0EnpV7zoLV47H4SDx0OEN6TufyXJhZMgvApM/g58u44rtW4PmpnfYbAPX
a7Lx8vDMAJ39V9lOkrZ0z7aTlxSJ6FXKR6DUe516y4c8Xr379PdSxfig3QZ2p1+bDba1w+CZl2Ve
Xz+6rds3A50ntWjLRwhwz6ZTF8pdUpYNcyJw9aZEFE8o/wSmD160yncZ/QNRX7zCQDUIVEKYjKz3
zm6nClFPvGZMycPbhYBO3CDnkk7nfEXt5hGBy8y1FDjDSYZgCbJstaXcJOdzvnBUPlJh7lVp/qa7
lcfVLXFHy+OEF4qqHiWPGJMghrCqvNYR9Nn2TQwx1yySBFfzXFu+pdCmcNKLicomIUA+rgw06OtS
Ukd/krB+gb1qq+2JF/DOu84W8rhoB2lnwleA7xaWp+YKFUKaZHNljV3YWxF7jfnuSsntTYaXZxgy
1GTz5AwuxnMz2yTFh8oJnw31E3cqlGt9lhfWkFQQqFoUie2lLDP4D44Lyv8XPddtuZUtSlOOGBeT
GCf8LMa2dSyntHhEIcL67W3TKk88CiIdrtqcw5ahzzmzvJMZlFmS1NNc7EFd6imIm0CFejgTdgBC
AFjPNlV1wRtJcGxqK2eBXWY6n1ngZ0ZqJT8NoUy4uR3QKnZl7K/hZ94DXlK9DP0xlgZuVDG/pLVe
Ser3L0s+xLWeLXYycQDcpsOp669mlYijuxFamtuR4dYbRJgWUFq2g/qO8axZwVRKiDCRMU+fudZr
lEIEGrr8+Tvb/kqrYdcJuEMIAbgj/iuM+2hwHkyNCXt7ujWqL9By3fj/v+Yra31AZ4Q7FZgWOon/
8WBmVYgokf1TEBt2CsBsW0flrmfKBIRwk0DLeoTqQVppUEOX/ISfMnYIss2CdyzfcK2nfwGJJFT8
P0EXXmFpnoqJl/cC6wpaOTtu1VctljfD7TDAfa8yBk9dlJV2f3zUflOi62F6HUMTgKcZKtdPNu12
F/jUKtrhUbLB81aHJ8/MdjXP4DTHiIhHWmK+RfkWU0WMGGdWBbA8+1+MarKZq5z3GoraAlGivvmh
ZtjHtWOckQ1C9oHl7kW3HLpD9ZDJn4MrfTaahai0M+D/C+AqQSqoDU56fAb8tY/1MZoiZsvX6zDI
G9ed/HQOXYTs2Q1ahyaCB68KrGMQg6ak4gdsbM8nlBDyWUjMYAqaYCNxjYKUSROPx6jeWL23P9uI
5xP7GV9Uk/Cr6QLqftAToYFdMlk3vQWqASkdBdlGjMCl3uR7s7QFeWXfmAI5T8maAWEoQgWJ7gw2
dpZLPNWO93E6s2VadFWxRbdDHKYMmv69lwdHLNtCKTKzIGoLUpEuunFMT1+LgMKAeVuzx2aG9AlI
BfHzE3xFHBy1rsGZAob/aveXAnE2Srxd2JvB5qNtJ01BoUUvK+0MQKXbCu2q2Jk1K+YvIo2uKUdr
HHosKy9Z6lgx2J0RmATUsZ2ZMsGpRGKNHi1yXNW4albgrFrAUbXAbrMY4co6ABWZf3qpTw3xqhyK
iymLtl8k3YXLB6YMdcUrQCBvvqYQpMkkvoM7DGp8IMoENn2CMaThaVTw1aGwVH0Ezm7ue0JUGRUW
LvVKM6LDhRMBXot4cFw0dPKRPBuhZ5Zou8MXuwlFhecbUZdDdy2QnmSFsqVJivnyw1d+sDL2cmpO
yTALYI+SNyQPZqMlGWjlMBMewdyrHFuXXIBdwFMCjfojaAZj+e8BSE5DQ4mph8APt8ELK+52jLkW
A/j1P+2eZBm0go5b5sgpqkJ/oZuFeTkjvZAjyJJSquyfQN2FXkzEQxHJdcjdkPiDTUSPK/VM+Zn2
LKYTpiH2Ct6C+oPtzuKHjrnZ1c/vokKJ0YDdRT1zeYSWB7UBX2ucH7U3JV4RTnMn/VG4nQCGTfKa
XXTeHUoSz4M0khTkL8DTtvJa8RBviPyUJjcne5bWc+MCaZ2/7iPqDOycWZgfy5/Oqq04zR8sMPIU
YXWnT1pRnlES/LHy/lsSgfQh2Gr3qZCVjcNUjbRPs/HtITSrqIZtkUUor+f/fbF9ea1Ke3s0qqAA
9o6+dWvEC9Jnw6sQifB0tEWnQBwIkDSshf9vimvbFWjs98jwDhae6rED12lyVP632QD3klv97rU0
U9Yv25Svydt5NRMXy8WqmlmUXpHnofEHNXDUfO0AuD9jJFuT0VPHV0Pbx8A3H+EIqgIgAtyjpFof
BEKZD9DUqp0UPPTCQQkY+5U4ZUDz37oJ1CbXjFnHI9+xCYWHKV+acoeXYcP2J6SjOY+bU/zplJmp
IWJtuuhtW6GCUl+eSkNkDLJMCU7b2OY+9y7XmpELO16j5X3yZig5fFWvZA1xTqeyGltetFY8u3mq
1r3FUM5pgBAHuQ8GgQin5bqWjECM3Jb0up/3lQBxaQVQXmCWkYCpSWW1+a6bpaEfeWfI3josj9cw
8+R0d1taLRW65RskNfxvL/Trw3aETdtQjkNFGO98liXote74Oky4U51XCnS908WSN2xywX3Tm7U8
SzHcFRQDVIkXnW1NABVBB6ByWmyoenh+WV3ndioNCRK30GnIGlcvcHPzNsFMXd6ICYV8n+Idsfjk
7BBDOx07bfey2Sc7kr1e/ZsHsZSldDVswM0T2766SqZMUPRTuTSHG+1zjeKZtf3RDn/JlYLlmbrC
MzBAT6D4zZFbwvhTATM8/r5wp5YRaYMrNgW0M9k/n6rfMWY+wukz3FwPmqTWxQwNyyPRfZSDyrV4
RMjMih3T4TPkOERmHBpZQalEWBi+Ma8MqojK+X9Rpl6ME6NHJCpMbzDdmzjpIZuB+fOoGs0eCUXj
cshMJdvfH7pwxY8olJa5qGER1cwcDfdHDimRJLi+8Gw5GV63qZyBMrbvHhAvSRL1oxlIwvyP0yrb
eRwM4eSGk8UepoUKjnBQN56Unw3N9kzA5KbmqLRo8aoMSlDRIKkmza6iI2Gow+esbxmEsSQ7z0Ho
vPXM1aJF/skhdHeGJ/t2RmSI4AHva8IHUc8J33dqjhdp1AD+ZCYAPMoH9sN0hGnGX7taUOkRCIQW
WV4V5wSpv+BQGl96iMbL8vwRBg/Av7Ai8U0YVKxkdqApy6P6E7xAGiBVNoiGkEbGabfTSfElR/9e
OIUoj8/X+ioLgAXYrmu5TpbkqF5AmXiD33jP82wkVzeoJQP52SUuSr1Fy68l5v0q/mNJ3iLbNW/k
53/s+66DQlrqiXa15omXpOs+91m+C66tlbWpZFY4dXmFEu7roumKVGMVdVzC8RaqS1bC6Pi8JVaQ
7TYe2NrIL0sBMHUoaREFxgLXFy2Mu95fZdllmSYpDMYIn2RZwgFVWe0kWBwLh9lKIbdtDqvYSh5M
hpSAQ0NK3ceOwRW2Z5Md8aHDQnXyXI/PFTnn2V+xxy/oHHQmws3Yx8aa8FKkMTA98UzLUyc0Sz8j
hoX3CGFlXGXSN529jaNIzPJEdhR1MbweuUp9rTrGz8vSN1xy4c4FLnMqZNgQ83bKGNMMTfDbJm9h
eD+ygAY5xPqlgWCvNP9K1v8bfeFlFXzlqrZtKHev6yL2k7S13M+v2BECxVywNv47UHOHs64VE8iK
IOkn64FyBQV5NTvQF0NR2vPQ4jRE2MgvxxBy3tMhrKyNG2gLDBPZn0eTjUxp/uLdTnZngXKKYiGB
OmRbkWwxbVROp1f+zCWIPX4/OoS17rA0Mm2H2HKl7Bdvvs2FX4pwj+mDGBJyj0u2n/X7716zZtEz
ANZzSlRRZ4LrVHEZw8SJcB6mQs/T449SjFqs3HGpS/AyUFdPVu0x2tND7Vmpuz7LRirYpL/AWvA1
ZhbURapQt07l0geMaMOz5ZzIXVYkZh0t/sVKujt9bF1CTOPnlMhu6EsfBG5hufmfNHFpHltrmcci
FgKn5wD7QfbqIHPg7zy1TcQ8d/3uVrD3wdS7z90kEuqhqlFakf9EEvV/LlIdZj44aZWMq9zlpO53
3/U9T2wlEKspZS7RlwiSs4UvkFiCLmg1XcOil937TWvPDhbe2yeEmNbc2GQRQ2QiAoNVcKZiLyto
2Tn2xU383dklYcQMBBhY/kcvmXwlhTPYidLrjDeZL9oCVoSPQqNkZKFFbHkPJwUfFi/ndO9MWf26
R8heHFDQYOGzlc/NxeBrLg0aUqfM4NBXwOWj7zWkZqQwG3oaCOAg1qP3qORTLz1sfZ5G7Xr1rHRx
/avurKDikp5eYzFmlgxDIGMzWiM5XrG0ANj56OQngLB7W1tSr24JV3DgG7tA3gh7kI5NIOWqDtUI
nN14A0k4gPgKeaahgU8jwMQBFws4D1q+wpeWext9906H9X8xOtdr5P8O1gc6R90XktFrxX97LLfW
lzXnJQpz72V+XPXqxrf6uO1gr4dvvpEW1RuFZNwcDG0SHq15EHBGgD6cIWB9OtmXpmDC6Z4/3Od3
AMVx/++PsOsBdofff0A57UEsgyZOQRsvoqGtnxlPHRZjzsegF+PZMMR13ZeOjTsrn5e09GVy8qKK
t4eFa1hUHSWQhpsag+wT0MBD6gBF9HQ/duHksSa9oTmvlSSqZIhiri9sgdA70kV3MUbrjjG9Gy+q
MP3Dv1E+ykNlO8wWNp1PeLvtivv5VKBzKkXuAXtcIcXmV714sUBoO+KZ23PGhN+CYHG2arLvnLcf
pMBgk2eZ4E96u56cIh9MJdd5C36zsWhU6Z4n5FK9xDzh78/fJh77sfAAFQUAGvH7T6QMmJvG0epf
cxghSo+EMPEq8FjbeYt3B5XKizggZMluHlOR9816lp+DOTQO5nyqp6mXLFgQAQzYevvwBSF0mrjw
QlmfpSiA0y33m+ahZh2mEnr30enXs7Ge9vmoZSaoDdsrLk60ew+jzHe3LQbIjGEflMFDRaXlQdc/
Lw1Sk0qb2lsC5wn4EvTLQKFdGwL9nz/46pGSevUvUqVjomDc++j49jqIoL6x7BgmTkEptV/vscub
LZ7/lyHrpHU4Jup3oRksUNcxURkAe8oasrSht9DzSR6VvLwmbbPTO/3rrij8qyV5GkSnMSgCzsgX
0lgsl9nP79HTI7B0o836jCqn88isBqwOkf/095sZrqqOfcof7sqYdth3JknvmlR3VXgjH67ob4uc
r3uO7UbZH9rEVWptfHronvmk1sai50SQqAAhdpyyjEhAbqHhjnXyA486AAsgva2bMPRBEqJhGqOM
RQiL6oeD2cK1No2Ix7QhUhncVtRx1NUw7PQfOEsEMR9hhLY+ZfBe2rcxgBoIR72bExehbeWLmWNW
axOz6/ck4Qs7R5cM+cJe0OdxSSJ+ezJRhq6Nosc5LHwR1gNWpfPKwcsUq5NTtxZvS+IGSWAuCHbW
PpeRa4y3wchU8jiy5pX95ZKgUswpKaQs80t26Yvb0LkvdrO+FrHYhkk6hEt1B9DUkrixIi9AgQ/a
XgWK1nawssDGgOZnPjfk5C9W5GjUxhvPRtE/RHgR5+bUsqlHTN7UgKTl76GpJvrfpgCPal+BwUAv
y2LQCqj+HUkJEwJqaA7hfq9GNOpejS0i7a17wf3JRL0AoqtscjjdPj/B+sC9ieQVkPvBuCdpn1KS
Gk5RfIqoPU6RhxqIPvQwUw3fUdPuel+wjhfAIO202DxEov/hqM8rNKKgCCUrai0FV7RLeu5P+nKr
1GUXEss+hESlEpyvjg3mkSMfF4A99nKQERxrsVXoNm0HR/OUEfAgzh70UP6G8fmlDQXuUenpKXu/
LVfBDYg1Ku1TNt6ZzRsnHOL8auh7fbuLf82ZBidPIDG6+ebPk8sBTSLn3HHcsz1boeVPREKf+bx4
0atZh+yk81t1ArHeao98txzKrmzAMQLq5H58GNoStRzpDe2HwlQj4mnHoj8vbNeTbBgoOgVaOMlh
A+2sUCUHzEi2Jpil8ClHTk1JGnv3vh+Wn21fpYL+V18502AnYLYjXozgAXS22esQc7PYjiNio9PB
w4oZ7sSQgF01pKw2WLYC4RCNqOgO7WuMysccpcxgpN/ZolKIcIfcJu/qdnkoayiLEETNXAFgS27t
JtmWoKVIZ1sSyxDXfHVDog+xk8EUX8ELRBBpIFl2lK5KAlMr324aAusLU4MdJGQwk18+DokI4U3D
ymGAV3cIFeLCAf7zbuS795VIV3VzOnMAcsTTttkiC2NSPFmm6roXSlbZUwkm6Bsj3/N2rY9yfnaH
IyHf9P43Jd4ctdt+amRY4N87C5/S9gQx0JRX1lll/6xkEBRPYIoIs4Y3Ct5uhYQVkcrh3/8wx6qA
yUh3sN/5N0Sbj2MbuR7hR+3C7NckudwvJJanKXVoZxoFsHVD+0Zm/Q1wMvWCRUxYzk9S/CWbqIb/
1ifCEioNGWxhKn6iTJn8x0HulGIMfb2rGDk3asleqMmZz9kmqMKBCKcb0Bcs3LUL9RX4yeoxsXjV
k78kLGN54yfE6SUGMRdrQkvr3xjAjA7CQ6LFuRBZxSuKtj4+nZK+bwlEAqaPEA5ZV0hghKd0gAGb
0yctJS6YlcyIB6sJgDBhhJOajIgXccNiVuGQy+OSmXJVT2/hDnrt6ZSyoyjiK2bJ+X+1xRhaB+dT
AwZK75Ol7HyJ8LtI7Gc1Aq7j263TLxIHgblwX/9h36grNXO1X3O5EgXLh/GpaS534gJszV7nMczH
Gxbi37lpzNLm8AH3+NwrWUsP2f+8m1NH41wsXjL6maZy/vDc/3Auy2mGOLddwSKvo2Ia5EhsCUgR
09X+1eiGuiMcu3zUYn2gfSt4qdD3Ze5zmA37fs1O9S/+UVdJcahjF0wdNwaCgMVEvrRwgan20XbD
qWIOV8m/K0D0stAGgvP5KzW8DFBrspuZOUNT6MxfQ2JTQkb/FqbiT7uHf0IA9DnZw0VqqN/YvQh8
HXDr4ktWlYiKQFBRnCKgETu+2XCxHWlSD3CYCMyPkde+Ex3iBXvZiFWtw9Fs6ePkEW+B0Sjcq4qC
JjG934M00l3yRXAknFXJd/gXRz5oFt3nvbcXnsqbyHgnvpz0LaANhshNqeGCYeF+dT0j+c3YjKJt
temL6Cav3JZJ9limvusTYHa/hqaIzijTg8a5ISby0K4TwmSPROTG40YMu6k8CrAxXxYtN1cq1Y7O
aVUGU07I8HONC9BCkZOxUXVE1LCV35Kg9Tx01GH0XQOfkRYJfYEfQmdZJFDw5PNp1AjxzGYAmcDP
RKfI2cImsL9aGLzAyjA7Xj/wxyZq+KhVxWwIsFGZqV09dcqoKep0w2QFWpcBvK6pyxlzMlFl4OmS
ph3NN28RaCD6OJ0wt3SlP5WksV//JhJ0jI9RHQ13uCm8k1OXoEsAesuI3Phq+bLwDxq8AZ8vItW2
9nQv/Ii6F2xyft7zFUvewk7dbl2of6VUELWGx8HRD1ffvSxO7EsAlBnsAzCXDuU4qeqzYF+lerSb
9KIR6P6l/Tg6YnrbGL+OE2HUraW8VgyKXJJtGy2nMv1rEX44oneLC8dZiYFDHTJ7YdunA19OiTk0
58bVk//GPKPrqRoT8gNVatiDaQtBHe6BH+nToVtnaMjKysWSeBOqTOMZ23L2A9VNn3cLapD++Bpw
w/qMvYDnLpjIvl1HiLTMvkJCHysZalh/Y61YvKHn9fm3q4ejtApniNmiQa+qf266B53dpJ3buk5b
9LfP1tJWFYjV5efI6ykyZn6FJ4DmqIksLwo2qqWXOFKMzvvpq0KrTfYj+arK5xffghailOlyWqV+
ifndecN5wx2MZH+z4293yBoWUt6BTi1BcWABN+V7SqukFOHFeIfOSbOzdpcYj+/B0s3zacXDaRXR
x4qac78BIu9IuYPZKj+5X8i15KbeouzXywzJQfb2GgMXpRg6pw/alK86cJT2WEAf6oY3I7XJ1HK7
Tlt0W6sMezQ2toCaL27RhAkHQjmn6BR12AKT9gczI+AFZpBwnDXbhs1VPTtZ15MKDUDMfID1lFar
1vUup3L3oX8AuTeA/mjHVh8zQVHokqdp8OxZRDa6YblxSDuYYYNjT9BEG87mqZ7U6+SQ13SR9f9/
xHD03BUfmDWjPQZrcqUUYW00b6hdeTzwXtKFws8G32kuTQG3T1RGioa0fO8fXiQB6RDScgsh6IMQ
COIo3lldBOWmOXkJ5zB3hwmhw8fCL8UuWwht+TGW06pqzOWVSTv04TdAgsRuJheCmWvwrPrJ8AS4
t+YNkIh9QLF+ol+SHMa9zfh5Nt3ga0A1NNLBxr7AoCZu6UfAyCKkQWv6D2qyRF9EzStki55MrtVv
eTMD5etG50FcHo0AG0znLl0+neYD7bkkkmWjAeC57pvuXiaigRFW1rPWWfDBIDQnn3OUAYOPVRXQ
Z5sXSx5BHuPVzquCd0MoDz8ikFTDEbqQd1yO2nXmygIytC27c+yoedEDObVEdU3XmPPrYA7n0H7p
yADtrTCu7og8M3aPC8xbbiFfjSFRlmqcnn4VyUMPUTLCo3Mo/cxMqOq2y+591JpYnKxTuHWtndGY
EObVQmkhcrf8hvBe+XjFuSVTzJYn7tH/IYyCtpdFchBNSi0S7K3Z9NSZmfbHA+aa2WEK50McnwL1
yV3yOChvHPusbX5xAiAR3DfNrHWa7yv0hXTT9UDSRUajkaS8hvL/0TUUPYlIT6Qlo2c+wmFPbx18
ZLGyhpzpvenaseIoyHbFqzg025fvWdzILY7h5CWbcNe3VA+3RKKXX6rI8d4Wd0cCfb3cae/9/DNZ
D5oRlaxG110WWsE/cjgrmBYrtYuhkcx4bc28usPbSdeNCLY1GPUwMvy26ebLiUU7zbVcm155ZTHk
rOtc4WoE8F11zLCbM7e35//fFix+Of81+aROvyid4fz5+gjxpZIAe78l8v38wblBi8p/g2lEMK1E
/37736+cbcwqxxypRjovc2U1vUAoKvcqtVL+DIFRONqy83wzk9ThQ/xHFPqx2wAUYnwZG0M3cLmb
R3ja3RU8U4PCz9dxzkzljsboD4hi1wJDEj+vrPfIxzGdMMj7/r4j9E98r1uB8VzJrWG5PpS8/RGb
801FTD7+9b8BQdL8JAupyM3YwmX5tzMsuPNFxiFk0Y9fkf6736pWPThv1NatZ4u/mjP1jGwLRLY0
iZmCEmkQ8ftz7asyryNv37Y/okYbJD8Y6m8O0XnXzrhqfqQKIrj+UshYxTQH+8SHB03H9LUupDdQ
VmXocjxWzBGy/sK9qi8Mklj+GptDbPW0JItWTBYJ23wMUJ+O3HF5URBHSYyWe0WlIfijaV1cJzee
f3U2A9GGeUJf9M+Dq0ADZ9lXzVEg488W2ZKM/2h29zjQ3+GFsu9lZx0+kiFlHYyT5sbAbN+bnDLJ
P9zvAg6Bx4oFc9W7td7CaiZa0CKH1eI7+CLdLvrn7p/0sWflPWhEMHDTNRlpDl1VovClb8kQFAx2
+RP77ixfK3EGSuAnKM+3KvH5HO7EL097kmhdyJC2NZyXxqrkZCLav3ynKfjyFdoLJMwWS8eoqL40
yfS57EE4qbF1yXAryu+7mF4gIoP5qR51AymB8tcwdqrDcpXDDEf9SErY7Mjn052ABlUW3HoH5BHi
tNicU8+feok2WLHr7F2o+TUCn/EMo18K7ZE7K/zs7dR9SO8qUsvkxBIarUiE9itHw2O+EQFZe692
RceitdGmupVfFHBbLoyrz0EXGo3ZDretUC80ojUHwhOOYFikp5FentA0I6TXGTQY7wCWBphD0zmZ
aMXCMGjutiRYmQAIRNRn+n1F8iHKwuddSDDw6oGn6Ctc2zH/Cx6dP5UcH+HF641pYn2tSYa/akYm
ZV8/bh/emF5aneBDOOtmLdEq0BMjvqcO8z7Sx56HEZX1+68q1w5k/He66XFyJCBY9cHsREc2NAHq
a/TzbmnjH70RLm7kqFbm101Q5uQOiIQ34wYPrmj6NPQhcy3btwicxiwuPpmkzjJ27rvGtJznUsOq
/Ees2PpFneEYxQenyDqn8in7Z44o/Mxkoq7VBY8CqF4+QhHlPh5JKkFv8YV+5IvzC0XQca0whLw4
61b9X5jTsVwIGvB8OdYi6w76M1wcoU4zNgzfqH8XxTffCtv6pwnUBANHbBhxn88TtGLeLGnsxtjb
81b419xaD1+mQG8s6spZWDuxIqub4vCKeuhJVZQC6qk7BMOgKe2NuNaOUkc9sAcXUsDm8aNQ/doR
uWz+O6fw+oqPVJwBSIEthxnkEsukl1r1rmS18ScjuyV/10sfjIabe8/tG2MJHXhpqd7wFj7gTRPH
nJ3Vg/jWhcib4uHdBw4Nu01rtNltfuGYk5phdhT9qhoWwG7um/pjIGgCuOW6auBlOE8gaMs7cY6p
SomCUzXDnX7BhJ605NCuE4IY/UVtGqU5V/W7N7Psz0T/CEtkoL3mv3ddh73QfG0NfgwyAwRQY2Q7
BczK2tQwJ/Q8k35wZ7oo6j3R5Dd+ng3nyUH/pt2yW5q9s10jSCzlcSKfv3gxXwqYwJCirLI3dsiy
FQrVjoQVjz/YRG8o5mffyJ+tfKOZn9UsY4QbGc6MQ15DU+Yv+VnEiJPZAaZXKtGs1p0nLef4kkZe
A3no1uLD1JJtqnzteuyGNIZt2KYQ65SMA3vIZCn0XqBez3Lx5/ynIbCX1ztRRxtjryVlTzeMH+VC
5Iqga3AmoaOzQEPT1ZgoLS90rEcyDn9S6oaAtSC0JA8GH/FVjMb7O2mmZ8IAOCvnN07umtNd96L5
NRIImLV3QOiqlsYJRZ9qkSNN+HA3t0JDP/M/kBV4XEC1Opa0ioPR1UoerJ3+fQEK0zFDuvgXgTdj
0wCZFXG7MErxpe+C7v4IWMZW9bHhIqv8KQcYlbEmrpMZn5W8DlIySIINLXSWhonAj3fFYHF8Uwkg
CGSY2llP3hyzPMqRSry9UNLTVQ+OqhghgkYYc+MfkG1mLI55x9sTAtvaghfgXeVZfOijBvXPPcNj
o3aozHvci0ikceZXFaFOR98a/p+18auekQ+N8+t0tZfk1tR+ygg8mS6Y3w6nvdJPqZgkLQ5OmoE0
djtAo9LheNf5CZSMFp8RWe+LdDt1KoxUG1Nl7iY8z5mj3LTf91AZV5REfGawJFUpy9MignJqJqd7
BVqewYyKiv+RqrWkN4Noz+o3Mov6tL+bkf2GJ86Fhm/nRk7/RtiO6IiEF+juY/JkFqLNbawmvNh3
K2gVeaU5iJmP9YVfkf4xFH6Kr2PsMQEKJVOAzMDub3yWWKrGiYFImavxOg/zep/c/0cgTprSaudp
38WUbxulo6DWdTYcF5tI69mIWv8aHVI83bKKY1m6F9S0hT1VrYtNY82sYJu0sZiqOddA3R8f9lsR
0Aqle/8NvMUNLl4Li09zrav6SVdJ5a2Hm6Ty1LbwngFFpUhjaTdOorkfeSX1sVHIRj0k1XR13+4V
WlIB2ZNR99hNU9axPSak5B7o+h5+CPenHKckAYNUou3d3AzLYIXc81YEaMgdvPYT3DpvkYFiUemM
k6KBmesHiHvuRpQV45mw5EBCxjmT0Ed/IsEIVVkP85uViK24zrZv5m3dmFIJoToExPGYBw4ZhG7g
XQ0k1hz12DejBdX8z9EtayRmKofljBopKFeLFisTYcBbQIkQxf12Sx7ejH+7HaOcmWEmobHNDtm/
OhtlTWORFdlEOk2vOtNk/T04o2CMJA+3shtVzkaJ59ccciUcMSrQZhQiPBq/o14Sh4iH6uhbCllS
kOW5I/4B4PmQCg7oIgi93aHl1UV7xL0vuDg6KuGzdqAu92YYgIBOGPLllYbdjB/hXloC+TYBpLqY
rWso9utkfZWWKuXRX5A/fdYLQGvXnsfCS7mV2buktAJXxDfdH32RmqYPdKARpfEh/ZhsEW/TUR1W
u/Q1QFviZUyBqOM2buX286UbWMwoaUUnoWGHQaQhxtyhrWdhi7GNE9xEMXajk9500U5Te44/wW6T
fJcrf4G3tb2VTdg+mRUGWu+smP7slFJ8TJqIsbgQoKb6iQDEM6/gotUBCKShCdJwmCdrbAxf/Vn2
Jl3UhZeEzwHXL0Baaf/8aOKYAUKFmofPHOSzYFjJEX7s2clECh4ubVMTqBt2ur0oxG9NSL2j0VlU
JmRDdX7EyfpQzbxdaMF4WU34RJBX7IwHGuZkIn9Acb7p7B8Ar8ET2dplKtBYXX7nDG1XZH1tUPj7
zyYErPXqDFgvafa8m+PBQvp1zWRTSLe0BX1p/CxngldHFjiSId+MIPN5g4AocOS9dk5IEeb+ACRd
6sDYkxaMBjRJDBXlKEqaNisRAawj7+tpZDcmk/MkPzQZkapLGQXSSbVXd8P1OV0WGhXj6AI7cFmG
xaW1IPv37dZWWEI0LXXVEL4LJzyqUV6UyryCPz/GI3DPl509ypZIF/Yxu3MWZSMS5P0VPj3JuyID
7qnHHkBtXYFMz4c6OB1nrkYfeH8S5q8QChII5bgBhwgSXTsyEBp9Q+uYwFnVY03h40E3JATvkOJj
QvCo6gNw4cc6BrdVUJKUHb/bB39SUafajIcXR1ysQqw0E5iUBQLd3PoeYWRHRiqvY+Cm8KLbnSFf
s3XB6dbp3z6aIYC2hDNvPfb6T9ncGdpiu4S71mJzamr1K7WkLNeuKUPQlBAgje28qIm8UTtEfHX1
UGZOPktyYjCEYUMJQxE6eEK3RuZYRaRhJN2rSwQrvPvpI+owWskoFd0bHQ7rQUukUoYWAWwf//1K
CePmjsmtow/xxUvE5BpWe+eR2RqJb7gleBODhx5swTarPQpDOol2vld4/P1dssCdRyICu5igPrUF
ZgntimmLBla/FsFm+MWJPwU5gqnv/TNrRtkj4LYolg/b+ZlhnVRe1RiYM4HalOFaWjdAkyMHmo6Z
9JMhd+/6Ljlxv2zsX2k1Dueo6gJmgSBIcQde7thqc9awXQ44VDHKFErwGepCTERbpgImSvuwqvcM
KRXT86HBOYqbkIjtApsPTPphLCaOgXjViYwFupnZjJmBqKyxvHHOJYNJUnJ6fiLWgCAK92DMi0x6
+hS+EGvADBDr0JuhCbcJGfzEk5pOEhZFeST3u2KNYfCBhlNUylywbQW9FsOORrbly1lUWLdSRGsg
byx2JvqGfD7Xv2XHci8RUOIb1pdSWvzDS1DPw8X/HgQ0wT4zXYDFiDR3pGrBYb8WwmYYEkuoLoYj
sodbG7RUH++NduiZqdeHYyPgZ2TPb1Y+Bn9PuH6IxOwgxcHMtPSS7+Lo6RZTtgAjjYGNQethWpGh
XV2Wukjk7qWtzkFVVKiB+8Kb6F249He/qcLmEh2+/zbnY9qrdtfgmqLiOF/wyLMWKeMVR/OTp1Sb
M8XrlZ22/VIAoAL3qUz+VfFPgBVyVnz9I7IsZLhqviWAQjZA/CalYtEs5kOUyWrchKi2HMGIWh/6
3AkoVzh+AttlaRPf94Vc/lArGyspL5xkNwGJV7QV8i9LQpoOrPVppujle3mjUUk651c01itPufZq
PzK6b+u3P0W8sw6ya0cwvLf+uSLrw8Oytm+xWMANgm6C7JPzc5f+jnvgjebmsQ2M5mO1IuGlBvoT
QphDfONQGBvYga1UwEH7eGH/xHDcCQmgSGYscLajG/wJrijiHYgsvCVHZF98qZZZgqbyTyG8MtLQ
iXG7lSfa1rqQXwWPObWVKcHBwoKM2l1X37ORif+ocoFAF8D+3I5DVbsq13zr/i2IpcNZFvHdR7NX
IrlNHH85Ai6aEQ2GaMBeFdZFakP7y07cLdNugzoMFPJ5xO6cKCf2tgDTVS6kGraCAPWf59jRPC72
POwQcyFiXKWytcyKCspLfwbWYCwnX3JMkExp7jgwjwoAY2dKvV4dSEZOErmLpx5TC7RqwEzwQZ4C
IhfrMkSBlfd01OWnt2cd0OuPgzzMUzGQtX0azfbpLs8cmI58EatZ3upCFulQA4Sj3XxufG3GwCtZ
KwG34lOOorQ1MdGk4pKjGafmH93fIbMZ5lUfmGq3F28+ITomycGNtiQnsByXnYsUYTwpZC8SKZIT
yvNDeXu5Epf/Gpt8inzqNmieiYspAolJ37Ivg20AojeuGPy/lm4rutAwcsLbPZz/QQD0CzGCrHCW
sAg0NE3DvSHe8e+d/yc90D7Qy8ILbgvNMZNrx+ty/0ESO1aZy0Y3nBWEKNCEosRAUc5d9UH8h1Ya
XT0pgTacbJ2s6JJnMaI3x3HDpIeo4qksfDvvmt1IH+yKb0nm+unVgNRtdRHWlIYyCsZUYSlwE+ys
6cIk5vHDIf9qfXhhC5vqVB+hYqr3hOhfY9zRgmDdzcnStG9xrRsnlxscPL9MWrq5mVyJEwgkKwC2
E1a4bEeJxDdRtzkCdcyf1CQYaX8R5fSyJbgbepu6fT7BLM2+MQ7hl4nRHRIWVlgCodr0Pb3BUGky
lzKqrCpoNWd8Xy5pHFJ2Npt+u8jXW6aLIrDrcjRrxcNJPgWmJkRRzczf+gWWs2U0v/fxcnFLAeSj
CXTFz1TQ4Dt2s69b6oNbROLPriIoC/CJ7ZjFdHPXSx0NFt89K7v2rX5K4vD4cINh9WJQcqr6h8gc
wRiaFJTfVXP3KOb+1tpcc8avUHwdTZJrlJ4z1RJ6GA/fchFOM76WEHp5YakPLMLpq3nO2hOyrd92
OZpJk4opyvA2Wu4SJMKaPdrbAz+I9xQoxpYZaJLS4d3woI6TaLpeFeGkFw5iNZROtz4+XCXOk9DK
Cy0s+Z3Y2XDHyei742ogki0uEiMHeZ6ljDMh92RlEnV2OiyeW8hW6b6e8qFEuQ4lU45hVWpDJOFW
KqTYjgIQBNlTfBM5VQLLe5pEQm6Sb+evfIIeTRgFFATJ63FX/TNaDsYGYCtbOfwcb1T6x3p0v5EQ
BNaUbB/aXv74vb4EP4t1et4gNsc9U0g2NySdoSz1lyfdcvh2wtkCoivnJdegkSRVPm8AS5Kz8bQM
GUNrqya5wWQfLt1gCdRxqpHkClwUf6jdap2LI2GWfAlhU3/egeAPj31LshCPlGTEeBevoTnbXpZf
1HTJFuYVQq1ED/n/OSZOHvyyCn05f69CRgMaqzbn8XEVa1pELnmpb1WJmWrUMjugJr/V6GCsUcT8
UHVLc843d/V+HS4WPnqGxQeLGNEa/eweyQ6sWATRFpFiLldbDNS2cXQC+sBdvRoH/IYbyjF+o22x
RscmYVW9u1bAacgtllfx4foDgR0YwTklfLmccpC6gX8rGGc/1n6GK4iy1HDj8uReaYU06J36wdMy
v0s92tNserKmBblkwQ94OrBfWEfJqYLRxNnFIyYU/scNxN+w2LWl2q3EStH1VtNhSr6UvQPlAFrF
vpyHDhKcgOoEcrbgLNs5vTgtDe8q69+TPDCX7A2mtoNKphNN6H6XIDdinRYQRsH8RujkHH6vg+gZ
yjv53VSERtDMZUZcz2MzCp75S00necpfT9sXRadjV1I0Dz7FJ8DnVzPUtkdEDREut+1XiceynsrX
f9mQpE07NG+gRjkXv4a7DwosyI4/KYiI9jW/q7BwzG3qZmMVMPeni1vAobHxGp8iAm32NdCnpPX4
QEOXXlAa2T/RNrh/BbVTLPbpEB8L/EuZIuNjzNNnpjphuExMDDwGMzTaNL3EHsk9lfmUA60rLqyT
tW78AbCWg6+AXyAUVyUWtpXHnWh7CGC4iZouxjKpIiKPY6TdG1LpAesW/mO2Qtmrc83sJb3PmB78
5FvWrYuXxaKQjho04ahtATMbfRiDxl6hPC6dYHhHLk3oUnzSel1vxIEC0RUohlR72q8q2emV5RGH
L2DU1vLZGJ3KIaHtPT+CJ3K1RsG0A5dtKZPI3wAmTpWIiqSHXmGaN1gLWGYsbwkQACKXejO5C6oW
342LzW89SHQQLbLYo97QK5t1MOHurHtRpgFoYU7D46dui419vZQHDy2BQozCbVpuZFKsdQpxsrEd
jm55HjwnUJJvlJfCHXdk43nk35Q0Vcn9oCa0tYaYVIeHagxbuYxIn+wxsiiNHjInbwlJ7+HYsOJF
FlLZtV3XnYzB1HZYtb1Fz8NAqPrbweCMoxnubK2Gjp/keioxIxlJG2k+ktEJOf8+SPy0KQ39z7Gq
PsNq2Qh6/Wh7JwbBWeecN9MEJhNawNDofU8Nhjhj+ueXPrSgIBeh/jCK2T5tXS+gd9/uuhd7beLZ
IpgZeVYKipfujIoB6dH5d2YFiDyGLDmNkOCVkj7YPDQkblhVMIbeeWNWaMDkDkGHQpK1p9qkZ6Mr
lBOymc0/y4JiSZ/afaRBk7vTnH8vm0DwUOM/WtxSDph+M/f+XMi1Tm7LH2JfK64sW3tXqPziZcot
2hVGwhJcGLRvR/PuHWP/nvXwuH+rvn5Bgn/wQtvZG/MmqUNWQsNB+NeV/jz25CPmj8Oz9ENZlF0T
G10zagIOiml1WYGucGljIS0Q/DelQtrsTu1N0S2WGG+T2884JGcOJWI4D1iFUe9p/dNNXJU2JzDS
iNgC/jNZ7fJhzb2P+aztB0nvWq5iliKA+ZNhbDfRPwJnmiseqxdktio1QAEIYAI8I7E6LJv5ZPGG
zdRb0CYi4zFx49kuDvaniLG+SnFc5HA1qb6YVLiXlGf9mkxP0aqhHhXcH3xvSY0wLPdzf/d0Ykhc
is4aKLLqpySY+7ovHqxAptqFay4Vs8+SJ5KRSHlM10D8dDB+9lZj6FOAPLPjxF+pqgCqZyAimM7R
3T4ffdIPn5pwIxKptPh0geOsnVmoEfUFqPRlZtrDTK3jd58syPuZ5ARoBXkKtLI0u9TePR9fRd64
r43zEdlryD1j/uDTzbb5hh05xjQLODWoUVIL6L/PR1treGa3uc4oVpgvu0utsm385uOg2b6yx9J0
F58GMLOvVeyEIf+OgABexUWy8rxbvO8cnRUKkX0EAi6mlCs5Gz1RqMAYrIPG8f5MS0qVn4Uy5s/8
mKE/tKSiRuQ6SzUHwySt5NcffkKJQjGQ9Q3UEfbGe5OcxsbGrOZk7nSuI13Uwat0Ho+m8NFprzOm
vjoYh1Y48IwJ3fNoxtN2SpPyoevgBjgGoCMmEmkYkqjqjddmDx7wRzyxq7Lco7sZktLzf5C/lIKW
uVxpR0mBOM9hBCDc4Ewt8NQl8ODXmjzg2vTouKVWTgrrD+PtmPFf5ZCgcmEtoRj3kfIKOeoSp3Jn
gIvpBcnihkR0BWOGhL9PUmKIJ6VaAzwo7XyUw9Yp9pGKpnhSMH+dtlef93ZMmpb9PZq1UBr/XGs1
Yywv48wQullcHQu8Jn7h3EvJIkN1iH2RMxngdHVZ1ZzXjwHEWIn1ilZ0G44k60HzT4cvDJA4RWk/
dSOBqsL/zr3VAHENg4HWf60fYRNUmL/FKbL5x/+bvqojzSQNg3l+NppwpSGjUvgbTRytjjBHmfbY
PzV151J+HL28ybGIh749+TeNW8u4u7pO6SUT8gdKq1lm3RqAVL3pXSO2SM8NJ/fDWJrxpGSIUwHY
ZH26hdWctFQqbKGoBvz1XeWmmTAApZ+aFoI32Urz+1YD7q8UOXDspyuEeCBn7uWA42c7qSXwPgu+
cWWMYu6PjUcvo84Ih5/46tQPDxECLQNmAKRAyOUrG1BGBgCk61hmCI1y9MGK2VB4oKBh9XksmCJW
KmNXhiaqNkQZrPbsjvXLNlYYNSOwTf0pW9IbIlofZV5IoDV27Y0JM2PdNiQebFWHLP5amm1r34tN
KpEkpGlwr39sGVUcukZy7c04xoWYUDNbudofbwGf+hDCak5kU3pCAGplQYp4NCm+oIXKY7PSwH+m
zUQW/5uQRGdOvENXRlCvmhwrX3KmsSz/jveLMTDDWd5eKPMN8Pqi9XXHGkNCNRuCMVWagGbp0G0+
PRnYmp5wdIYhvS+koohnwjC/jDA4h0QLwRQs+f5OJOjH9iFyZj0mJfKoSRy7k3Q4w/4Jq1t3HNHz
0JtBQeIsvC+Om7+wxQJQ+p7wvDHs54/DMGhCtq6J1Zk+Ojo03QQSv6IUIoc6mAaidoxKMUSAJ12w
TmIGWA1FyHDIVaXl0Xe9lTEWKmoyxfEe3hg1ARHhBaNIOKpRTNHKFfsZKkPjgY+/3FcZUOxd6QDO
UBqm8k/8qgHz+B7Uq+zjXnYEcMQMTE4QdnhjgGUpqnSZDlVmkgAlgY3qgtHIex/5loGUd9b8b7ba
ycRXhn3YXqBGq6x/9umJqJyfJchezOupeSgFko8qFboNvLXuOyu5dpppHoq5R1C8Zi4qJFGQy0I/
uK5UbtKXTbTxJa6BWGDNFVc98Txcon4BOC4pKs3uWx4EikL+VLiY1T/oFgn5Bfc88IKmo9U4g0Ri
SH6OgGtogo6EJexChCHc54G2baSJOfM+m7BMDtnbAvGBjRXXNt9y/mQDr6e2xYA+ywIqqONjkBuq
7x2eBFDzHVzf3Bm2imubtBBelk1k/UtTTWpjc7ybreJo6xMPaydoWKlIXVDGBSG+I/o5WiYiiJ7V
W5lTWNoHP4Dlqfbaq7vzeZn3G0imVSpi1qEMKbbvqXyQ9yZ/JzW40YvDfa0kW/g1YqaDnrcCQ/yK
EGCSK9Vn8ZbT69oElj6l1ShaiLB6GLUBTKroxm14amlcDQaVRS/ULtsGHURVfGYjuCGITaA/HQyd
UdawxuJdO6WNA8Y87dIztQcrsdIfguEkcAt0XWszKAz5USytmZGEb7YWUpEwdk0Ume8jpIL15MzH
2ZU/NtZpEj/SONyLGKYYqV5ix4OUT/4+N1K38wz1oziWb+qkiqfnDtTam2p2RsNNi1FIryEHUhVM
doGLkJOwd+ulFEPnBtIEdBYQXU5F8NI3oKNCcCpcmyDFe0wrqm7P2XhI6ERQQatqWD/cbRtVswIK
hLI4qEhe026gsStmt2+seVsTB2AecB8X7rct6k2P1cfbk7oJOGVRiPeTc13taPpebXFQBLsqsYnc
3ugPiPDg98VmEGVr8BbxbHLKTMLoqJWiSb0PfI8YWxsiFi3gJHGLqMdYguWqfPqE7nE/+qSQ6bJp
58pdW7FZxK8DSsqxYmLaLcwUuI9sB5vEFtWWkHfFI1FPlLaLZmD/Jk7IlHtlEkN70S0rkv3MEgsq
i1K8R0ttUuGaBCrSVo8B7nyNtBDtmvkTGSKdwYxMMdA8OdhHXD5CS8SIcEf2v+ywJ5C8ia56L5+w
D2mbEVmclBIVITuc+qe+3GVO/9hBS1X6P41JzWLxzNTFNTiij0NNdbxBXTUK98MeC6mMfwy60XNn
2bGfkezrdPFwkm6GDVSh1okksUF5h2+eQAE6T+STaoY7Iol4nGkRROW5qExQdguEqR/d9X5OyfC+
BHYMJy7GfjDeH0MwW+IgDDn0qcOW3AfzyurZGkGUkW5BkgzRfhXmWfjDgiZg0c3j7pm1jpAGr9m/
AgDnW1wzUraHznMOvoxzCtI3bhleh+OSr8H9fdPXDOkJoaQAXPnPgdIGWZ5OpmrqPCZCPxn/cxm3
ZTWMfyFoYPoVpmOjo+kxXffI07ftMlAuSbufxV7LaTEoKzyRZqXbY0pSZ1ROHQX0qk76AA9hLt4i
l3GlcYE6+IyzchDc1hsPj+ulfsG2qFOK3gXAz3w53A68SBXvsAHtvS8DVIzKFdnKQHS2QtK3CXcr
ZxtmvBX+8atuyqpZR1BLefa1fLg117lOir08ny1c7FTeImXO0Kr33UA6i9xibR7rPFmxzGP+Goi/
GANbmvEKLPIVa1Mdx4a2vJ4BUFlVLpnCC005920FtOcffU/pwe1U/ATDKCARAWkqHbnd/PzBcHdo
jSLxei32OTl3LDIwWKX5yl5/zyUb/QXfx3Hm9iuDZWjzuzrtj8CXUyhwPc1TM1UTGK5j/B2K0cCF
KeeTei6QfCHZ9yJou6LaBMBM9pTg+kqQI4m2KIh3vW6dbZ62+7L+z5xGSl4J2LQdJEEbrOSsJ6Q/
aNzmAHCGt0WuXLU/6doL8ckyVFY3QP2j93jrzS+qsq9S7Oyl2oj1I7U/NxuPStTuGjlNiHxxYNDL
tWhDt1yjc3E1DRdoULK7Q0xmVylT9Qhve2ePG88WmuGmbT3dEYWczBfqbz1jKDMycctFXqBvXlos
C1ArdqyQa+EtnQMtL5Oky/fdrvxx3Nhdkb5be0bc6cQiiaxU9h2W6kk4ENiKtBtiYsYTde6rO/LT
rbt+liZ0YAX+0p/xBDEPPIqbt72EEKqfD1UgTuJAG7LIZXV3/iVOO1Gv3gbjLE9Jcg5LuOdiGnM5
VotWlBnGoZuLNkoEX9EkoimLkS89a1MME+ANAV4leamnT92SzPoNwbVgmVdlP7gGj05sQn3r/vPw
L9ebzewKPqhdqcKcdiypnTFZCIYGOjiBW4zjEm05ri06AFrIh8cmxLSe3VckDG3J7MOPa13lqsSY
E6dVPmcX/x2U0+Qk4tzKlGEJ8UwrXGHgsGsidAeYGBMm/D4qyaQkz0f7sauz0CE3CGLsSvhm7Rhw
2RTX9P29KanZ5j39P8Ye/YvWX2FAULnyeUaDVkd7ZQYpTFuz7LBbwiI5liEuHN2g2rp/s3DgS3rm
QjdHGrTol/73plxQZGidq43hHJWwTdzVhVSTIS261Z9Q3f6XuFimun9ASXd3MBlu3o8r9WXV3Vrw
0Hi2kUpM8rUnbQn15A036TUNXa7TOKzcy45u13VyHj48FsSydMJvEipXf4+/Q1EZ0h0LqVwHkKQh
te96bUKZ26f9Q5wvxqBejZtWjrBjB3by0UKkRRfRdB079xepi970IF7Mus9k+B9qvTGm/WK3fKv5
jV+1UonEdNjGPgnmnD8CoJDOSggQYrwP7Vz9A+dtXlL1pPOwiBLRV/o1F+xe9OYXLVAD+9gfshkL
kmkeg0RFGx2lvQP+fpsOIpUyx4YQ6d3VglCTsceHuMU7kq+KKwc5si89jQdTwKjWL59ckIKIEEWM
SElfVhNLjkd3oMUBBNEVCu+Pcc8pyKWys8XefDiEyZIeFcWhGOhD/FZ0t5ipTohPNrtSoRmBTd/r
gQhco7OfXdT/tWa2ZXDrSSbfWw52U9VQ3VwZ05cIbIworptSfCNxb8xC3lC+MLNWBTVgwm8obQvX
YwNE6snBX2U+8+x/YbbMWDL03xNduvsVu0HHp2k+fxIC6ZnzkX+mukCPCi2ETZBlR8PBfRhlxF2V
tGJFP03IWpZMM76PfDoidqdDIzWe2wNiE7hY9tsRV+SlcXec34DBQ9gV7NtTAdO7kOquwmv50qx+
S1uA9Q+fHlkw00aYwuCzOnUKMYaujH1ELZW0TcA15BOgcf9zIEKePwx8iEkYMjlC9MF/PUNuhguE
2O4ArPXPJB3hEFnFpzwFEQz2hNjGD5n+nKwoutoGq/izo0iGbcFE5B4XgnrowLKeK/NCdewSAwyn
NSpUU+rMlf2ixB+WICUzci0rNsR1iR7Ffw5BWUAJi8alKV4zrEILG5iUqpL3EJzcHbHAYmNGMXq3
MNjf3Ev7Qn+DftMo19X2y3j5OrWKKVs1JF0vGjjVqGM3/Vz7QdsvL8h4J61tiXC4DVxayzT5V9q6
GMUHBW7Re9PRUh+N5zmXCMG22OGzOW8YFV59DylEKwE8YC5GisaZqwHFNgeDei84hgHDhbrmwe9v
uqPJFUTNlAsduQvQ9z81q8cAhnfnz4tQyGdsHS3zcRw0ELQ/XMA1tF/wt6Z4cHkSFq6zyH/3evJp
rgur1lrW6+DcuL/SYuS5WyRqPtd+JKSs4U91ao/J9uv8LJoiQ5H4+bXC4hZNXo+9hjXNDSakt5XS
Tv6mPz+tbrCzcRyI+Eop23YtG4y3/ZuZLVn7/377znfcaTS2r7moiDdt85Wqr67pf+eckRb2QDoa
RljP6glMp8tMwJoOvnceBJE9AezaOc2sgSpk+E2+jJ/5rVuiNE7lEZON4RNyEHB583YI+enONWLS
8ibxQQ1c+7HaHWLv9atDvIGdLjvJnbPHyPqhU/iuqXZlxeeaN0NOj0cjwG2d0xoQsO6yEnuKGnqd
oaiKU3kO8zM2R3UNjnAe7FYmZsEWHx8qY7FHguewfIiQc7j8UEjQuSBm517CrJUrlkr+Oq09iULs
mNEqEvBV5qzFnNEY+Q46b+/sDbfIYE3M1jFoiPy3UG+V1gSymppojX8JsRiQcBZH/d9zl1f9asH+
89AxrBN6d2wG2l/jqSdou3f0k1PfTurOwwCLulUCTpqywp/2z8dO7ALj01zWhJBbQNrAq1xBpz0t
vRFgWHk8XmgMsRVEa29tKW8TM9SJV/qbUgQIcsHI1ug0G0u0Pxz5t2S2UH5mHcxrAvNffeyWUxp7
Na+jMfIzVZlctxC7+hvrHawE77eC1KxdVWmBfD8SgCrHknWnf2aHEIKHp8m2vOwlXsVjnNhI1TXH
uibHxU2vOXwts872O9HpYW5tzrfNmEE9kRWtqPVW19QIBdc28OhXl2zdd0BIz0mj5Mg2FagonROu
HUS5skaA9ZQgCaGNo9OOYqBBPupwX2vbu0V/R1Bp/dHpaLrPRdgLt2/7BWz+ihYARIcf0HEmUkpx
2qjzKY/Qb1Os4RQrLZdJIg+ZpUzhd+gU69gVdsBVErMzhWJBMtlOQuthbf5XiATebyag7DOGlS72
s3wm5teS4PdnLamtYh32xZXDqrkREbGJhxA6a05YyaYwILSXiQeaW7ke1sOcqayHuDAsA3Qk7RCL
NBR4TulwvfbG9gMvZFLXZBAG5WUFrvwVk7BOhLLoSoKFjhn41aM40rK/qIMtao8sWyNVdyGVxLfs
l4GBEVc4uBBKYRUg1UdxtzhiZPqO2yyhPF2yXUdGW4JAtMfVQnu/iDEd/Or6DU92b9xvsYdmg0Mv
1Abce38/apwYQjJxLSNVxxRLDu/qsyE/JGD9fxLjLT48hpqq2svcnMdWwOzeSD7O8AN2xtslgpqH
+yA6clHckpKium4xsS6mmqvGrzJpxNnParogskn0WOwiv1sWfcrQ0UbYBlk2KMgJiCtVppirtSQ2
ZJLU75c800MfZMncZnRAdBF61kmYbpP5LrB35W5m0lpPJx4/3yxdbc8JqzH8D9CYdR5v8fx6aKW0
13WbpQwl37N5Mw0Mdv7Lcs4cbSRlHsf61828avVbNBouMF4kxTmOfE5ygqIp+RE6qUPIeuolL9hK
dbXP9pyHya+/clt37Edzv5KiD0KJMacJRhOrpA6r/o56GHFaCfyhCWEuS8zyd8A0tVY2Yw/m8uxR
zdAAwK/Rgq/951smwgK3JA98+csmXcQtGBLnT7neyXSmjunfsH1QwMXgnbRNJ737UEDLBtLp++My
lTH9hZ74Yr2Nx2ywXKdzRVVaRtv2nZvNiVDPO8JPp8Z727tnC71fRxEffkz/GpBYqXTq1mOYTHqu
GPrA0B6ShSVim7ZZg6Z5ltgWsGMlJ3Uofn3nuW03eUwVtbYziiLsIddu+07Teb4otEk+NX2CR3Lu
ngkXRhBsEYnbkPx1G0vOtjXA3y5yXDMSTpiK9rrFziQMMeRfb43DE6P1yHmTcn0gOcHJdrvP4Sop
e8w3fClT8faaogEMsMQuDXjADN4rNyUrJweCN5fgg7Omw4vbDFdH/S9ojyfYJz4J2zRm+Avg4GjV
CR6CraStXu2EesIKPDNAdSOB0OucKOo+eEP2eP65NRb9W4zWff+Im+2WpP81GwBUOLHgcgU6D1tI
QVWzuxL355RLI2jJfwcfQQ3Gb0fVD3u9Qn0Us3lznm5LxbUqe9ngDJ60AFDbWkgxEHvBM1QP8F9x
pFsE/fwGk4fs2uGM5Sw3I2r/MNLPmB2/hHchnML7wamNQz7QWbVhv13LMe53+mueTjDKcDY5AYxd
neMwoXM9vLbyPDzG9VcdfcrrnfkMqUjXm4xuvMtTTvVtRmpo2WqWEE5DXTOvdmp59B3V+vpbS9j9
E41zdWzvzEX0zpqIdPaCVC3EvN6XRxLP5H456xTmBxvcUnOsEUwNUhoFYGMc/ot2JlsudDqwxr+t
4Q7LqZOraIVa1CO8PF/RyB7r1UzGJYE2MQjaiL4ox5OtUyyo4oI+sxY/oUH4YFN8Ulh5he/V9PX0
Vc927SQw31Z29xAZA/Qpej9KyBlyY/ywNpt4N37YUQ5E0GNT1LZTca6Hzx3AiRfD4wAfb88FQk7V
sH6RipuydVd7hurMppwKXsdSDjX0Ts4A81hudqqaiAeYobhYlC5paYxyn/5yQM8impYImghYAoeA
U9ta+ZPwWDMSk6bxwETWXGlSTs1Y5r5cdHFIy/OYxFYag2LEqYY1YCT0mh99JKL3xK+4mG2ylohx
/XYg4bkR/W5dypZXo+mI1XkMCeaz0LKDXQww8lZmGcKsFfWxQfqbNCBWjAXOzHSOlKoKQbAkMX4E
/kr8xv8tZaCjwgIu+25bROT0u7wx9DKIbpGR6N/VvVYmroqNoNhsvh8KKo596nkjzcEKsYIe01Q2
8MKRz+ZUG5KbaYnzpolHx1HtOXXOwa2JeJswJ3LpP9e0pT7I90ysvxUoG3GJG2xqB/OhzRZKWzp0
NJHlpXReTgJylYCArKeBF5Wz6fbzPhPsRRAVQkLoka4qC6zqY1vToognlGNNkgHZ0m30SnJWi4kD
Jmf/GzQjQk6iWrWinaSW/PSSfQkEy+QIRvWqnNDoCzYCqwp+tYfuvvrlTyeqi2RZn04W2juajATj
ARKQkHap6WcBb+KQz7K4f3Q5NvsaoQce5KTm+xOL2KsLwN0Tf93dgl4WIbIA/OhMhZmHkEhHM+H0
Wur2Upf8Lc/JwSGGacbznUItsA+gw1UmeAXCHFekV5VnngAnqcfU84ENB/nYbqTaDo50i8kxisg1
0DlXSbpkSCh5/WwvNiOkqL5FQ15RFRoZF2stUJmaIQYgr8o5MmprM/kj/MLDQxv0hRHHkjXQeSV8
7u0ZitqaTSw3h1F/0d1gCFcC9woxC9sI3TcmgbuphBG5glNoWAGGe6hOgMCLlUwI3iYyHfDd/Keo
w6GIiNWFYFl+L6CNJLfMH+QYVr6mqHp/gH2X+ccw0RqRHg2PJApTG0nBg7/7cVc/IXxBwCPC4BlB
iWxgWVmWLGIc94irtRWAHBMZcKPDzYJl+5XHG+4mx05l7k5LwaUalAuApXUhtN5Uqe5IAfL9To9N
QgEcnbHJa9+9COXBRNrXNbiktYpKvOa8df0wyv+rSwZgGLNtfBIYEM+sY7PPjiPRMtECLsfoKcOd
RdP+SzS4qktKrAMvljwQmQtyDeer7qr3WDeVEhEmt3VJ5t/+PzljpHK4XSWE6MCblVdepjYV1rZf
yHMJDb2j6YDjmd2zVeQsBWfROqpSScQBvacfsyuzH8IzSk+5EryhDuS5Jkc1/W5EPEkKuR8JH2I2
x47aUxrOyoGNCFAu+Z7qsaPbSochTUBL9kpq/v9NkM0k+dbZrpT0ddKpT0neOQdh3uZjPNLQHOiW
nspeXhWwVwvoqrBQUgOCYDvjaoYAWQb62IIpMaj5h9gu22KCQhC9tzTCU+g3LrkFL/dLBDaNpD7T
xJDXOvNlisuqwVPnxJt6nhfuO+Opx84bhbuNqMMg86OP3hJORQaNowzOp87Pn1WCuObR6Ju7g/EP
In0ybmvFxanwu/tahd+rSnLhVlkRvu4Dhy+DnLCMlXG2tcDiKIN8SjcXFnrVPvacjeXapFKYhqmu
TrFKtKReAfIPOZk57kJDW8xn7EEMjUpsWCyWzr8mq/oqkC3SuP/ay5qpwwDQcyMvhLcjlgoT+wyE
pi8N8uLPJBZsfrc8z5WqkwfvVo6IzHtYN9DixGpoeHNaRjwwwyJLn1xSXffUtvUE7Iv8tUAcdRUH
1z3lODV+ozzPKp7Uu+qDcTD72ThTeMf84hoKBowdo/4oikY87BJ3NyPcJSHqP/C39b59emp1oduL
uM8amTV9aTE8ru4Ur9omUfoYqXDVx9xsvuwURzmdr1STlPkG+QeOLpwQ2n6nyPTC1JYnTFzK1dKj
xYZr+F7G0SQO1LMmubs0XV3tKyc/9m1SGpvocVLx/yhjJraVagwhMYfW1Ly5v5rk/ILaxmZduVo1
mGnVnVxBIgV+znLzh24bCVij6os1xOtnHgtWWXANCBsZOvoFtO/ab7NPWvOnKe5wo3O7iBrHZZf9
YjljqjuoFZdrXt67q3rFRJGB7K4/Vbui5uyPdMkP0vHIT2ZzOY0dFQXxqW21ARGDI86oaK6af52I
KLb+Cj5fTbW0sn0MLU5/U0Nj2aVZ5ShkqB7LtAEboi13BVSt819LNGJXJJPAHbQMEOk84OPbpnPg
gl8//IbN35J0ql8nD3/Zm0Z51IlXbZ0lTvWoa5gomAhr7ebjyRaaHM6rACBE6BrOlAuFaOlcaFbO
KYU9I+v52NRcL7GOqZrLxT29Doyn7GQsXm7zUH6MAIOjQmFCCPPvTwXvdNs508p6hMrbGcouMukp
YpdMUmx69hjH5gfsH99ISG7QZ31y+K/1HlsTF7KkOdDSQH3VzSlkY1ab++ZfeCeYlcdywCzI58O0
CrCRvSjrggFapq81LGqZz5NJmNe7zrrI7Ner5y+Wu6wKVXO3IAeIBZ0trMj0+7TEnaZdLG5kRfIy
TQ55eCs4qYO8tiETSq5JhyldmEYVOhhltqHupKaUqzeiH5DmYMVGXWr/BwZW6V0GyiPGL0auXO57
GZjL6KcwOIdwbXlZxk4Kz49s/qSRLs7kDGtSuzohwZItK5OqPpf57ntNtNDjxQkZW9cc6E9h6Bct
RbETCvsQiXq29C26qWa+ajowaQdntfUMCA4i6kAYkd/HlwA3Ph7rep7gsuyh2rujdf23D/4BTkrC
4kX8AkLYzduV25lphclSThD66V/o8gNfLMiTUh3w7z67xEsXZkY2Hopx2H4uvYn2F3TG3y74RgDZ
c/0MUloG/kHBVp1eTiZygcSWene/t+N2uvkEUrWRjyZ8DV1OunqvwLqHt2OcJ9nWI4sPUZMkxgf4
5OBz7iCtTEgPLQ1toab0ZWiDQlNjQelGELn4c5zn5soLTWi7ALTHkRe31waLwKumBNILNXUx7ZWQ
gArEk2WmXqKm1IXWqPtoKpDWpfDzSMMdTKFlVRYgSfXDygAfFTFLJavscJdSVQUktz7uCPeTMY9K
qKhKUxIjQ5ja0Lc1cduV9u7KhHHK8qAbVTN0jOMaPh7O7Y6nG6iw6fo+THRO03tuo7zUTYj+eSpX
YzofgeF3UDAnAUmI7mjnLzlPG0NZuW41rW6iRHwQO/HYFGnLuFhMGwBvawRbu4+6bxvARsCRzbeO
0RIXER6iQn6sTZrtl0CbgcwDdTpP0sbB+mVw5jDwzc8BfzkL/26ad5+ktdDCkeBOMKnv1MSF9rJI
A/0UclnYA9HrScLe6odmNqhcDR3lrlTVX3gwAI5N4+YL7KH9db1s2heNuuaEz65T4biGDHv7HfqR
Eiqol4WMSKRZf35yVQQlZb+bbglusTN0WLxpreWR8m7G2gaio1JltB9IJwM+o+LfArlVS6n3gPKd
gQTxbh2+LUdkWNPCtYY/MoP/I1SXyL3k/zqPAQuYgSPTOpcOAmNJv+RvwI8kKCSjo5UfD4E5jqol
uxDBxl3UD0CYp3Y/iqdkGRv6a5KSpFT14HlLTLluYsXG6OI2DOJDjCiY946pwbWAlV799du4GK3Y
vWiA4rYOnBXTqD6QOE++K17du5uenPIOkdXDPCZ08ZvUvI9yMt8ZbVI+i8S24QubpIb/3jAyaz30
frg0a4hFILrK+6vcDX8nOhYMrhiUQkXYEFTd9BYihnk/S2ucZVlPSBlMH7mPATDVGlAgNBGJrIg7
hRzvBTXFyLXlnpgvAxLupV1PWxRwAAwpwHazOUlQwZ+JCFr1wcnxHdVKgohEZ9gf/d5Y1QiHs60X
Jwa4elR7n9NsZvXera08d/Etx0VDVbFXsUpuCnNgVWXwtuCej/bRemFMp+oen2IwdbNpQ3y4WDmI
kxaVcrnlambFdkl7SIkLq32zbFkRPK8KSyHqiecvNVw5Apf5A25s3h9tStjiWM05gXV+Gd8tEJ6P
YSFCjBT4UJaimNZ0fMq+puamU2Apbn4WxLAwRMpeQ6aWem0rapCRKcuZ/mh6XdoDeh4WXw+HIjSR
M9IM5v+dKhCmHoCow6Zn/vx01l3vHHugIIC+fAvvQ5OckLX5WpjWx9OvH5oLBCIlbyrgrpYd+cTo
M81/Y4Wx4euHybefyhvMjXYYzCVd2iruLFgDf80O2IlLXFb5BjLg42WXD3ftwGPHkk8svK+WTapB
Ya1jOUCj1EorU7jjXWVDGUrhdZ10hiyn8jmRUzXU1DtEwCsm8WftONo+Qsxw92LzDdJfxMhPjkKE
mKHWTgv/B9+Ria54nVFlIc3u30Fhq0XPsAJPMZyiG/zLqmsmx478X/hT//geMObdmuErkGlgO8ce
76C25fNKPWyzCVFa8stVM3iSrArKM32i8b3f7a/hlCBVPFKTAXgouQXN+ga/u/TA01XEgFEdUqAJ
W3Cu02UMHZpomach3gYJ53qBsC0G6ioP2emYNWpFg6mUeoGLswl3OUOng+VQrylFg1kBNDaIcuao
HaTQ1tCfZbctp5fsDpbzGVHxnNZZHc13nc9jq/yFFabD1jpyTd0cXxF54Rs6O+FtZsrPAShLqlTC
ZVSfItpD0m3dWWokQuJjgcbC2hdR/C/K9WSKKfu83CVdEaNU+wyywSjxKvibMXLA3tbOBha/Qc/7
2p8qu42vurluRuQXbDtK2ObGawezomz5aV+0FqPVPQqOO/4WdKNEV9YpXAIHk0SVN4/mqvAoGXS8
EAmTvmqclwvOKTA1cYQWXZs9gj5XUSNGFycpRJh8vaSgzlgbA93ZwQpA0/O8IPnvJ/5kTfjUhA+w
YTUF5A3cPQUFVKmmu2JXnKE7ye0t/sJ4iNUcsYxwlUPcKf/927AvLmwpUCXMoCJUe0U1ixN1jECh
+7bnY9odubaI+tRZoEW1H3DFEF2rb/QH/aQI0/2x/k1drYZdf/vuvsv8mmIIjblu8XmrbiR4ZsEj
vZsM0S4SwRSouDwvHW/3vnLDtpBjWjh4j9qiYqkd6tE1sniakvCMDkBKTPR5Xz0Qitkmn3RYPMVj
aqdxALX8H1T1aAuS7YZGRSgWVDKmpBjtILCdm69l3kfzVGa4fv7KJZ3YclD2Qygw4B+MdNCHKTaj
Kne9Zw2oGDEScJpoieU4PYEjBRXQuDKOECJsNcl6isCdR/jS6mLQTl3L5WKw83igAfvJV8thKDaQ
79Lc9q/rZ7pMqGyr2dMkvZOdJr3eWMeEABR5WIVLDQXSh7UbOn/UOq5Fe1Kv1JZMxSTjfPpTfLCw
lmvJcbVNDYQXv6jtYF4XS5lSsL246OGg68cp2FtN7i9yuxZ8TXSgA6h1haGQfYgmo0SgmI6yc7k5
TooJwbyxn4qJrrP8qQzh/DxVBU5SsTLqu/wRw1Ife0xHSxdvmeTG2WK6URLI4z7sJv95tgiGFGTa
H/KpqoClW3RL3X7x/OjFercPyntCYy3UCrlVi6YOA5qZCZwLoiNBjKtNVlYEeQkxpn7ZqeBdRNRg
9oSXxqHZ8ENHaEcogEFYuARoicTnPS+PBCPb0cjJLBSrqb5sgp4iu0jurdtjmktvUrpHHhJ6NCqk
FL7Sbd4bw/0oD7SlCLSy2/rSiQOtmcSlCCP4yAQzwUsVMrjO25KqGV5bwOKrh2q1MiSYEl0Eui5q
0vdDeWQSyyelJeh9uufKYqDihOkA7InvFcFd2fOKKeo6ksLIN7V+FjzXGkm/XNXzFGLZRFqdv41q
ruC5QFoAFtr4ghAZJv4Qgaa3cm7jnCZN7KzrvPy9HGmsyZqqdy6KXN+OAucqTVT5Zd8jSUqWJRVr
V4Q5aUL/rga+Ne6K3se/J/vedbT3waxMPbxVVQwxJYZ7qp3iw/CaTBbrXhqy5PeEALS5Q+XR0eZ8
yHHJyGlp3pQ0SS+4nGTdYdlF/VYc94Sn3UEW/mfNX3ojAu5g7oTk3vKh4s0LXAfWYJQjY+wYYdfj
PYPR9h1Sf/SLu+gXhdLDkxGGyTuERw2OAT/t5WzTI7N50oDwq+FpvIhVNgJjbUUVXrWM3mZZFETf
AZFRdCmto7AOiXCX5n94JkjeyB7tZ/POkg6UQLhU/Uzh8MlbvYkAAsY8IuCkc5j25VuDpuTwf8RA
QNBhJZJPYPHUEoquIC8E43SgUyfiVi2GkOmJG/0NQvnVw6CRoaN4bjE07V07a5Pgkp4WKuZmir5p
NcuD7J3wKbA36+55PV37FQGu+4E6oIJIIOPZt/POwVLk3fmhjDaVsZ/3IeiRrPZJsBYXcnMb2il7
XcVV98IKIv0T3P/+1MHMsvbT0uXF0JS2t3zzRXUju9Uu3GBm9Ex1HA/YKNSz12cgwpm50btemkB+
ret4dqXboX3thQUK6QDEa/Lfmb47F6GlNHI79QL0Vo78EKzQYdNWbJUjfVRZ8nR2XMUq2UHTWsBb
jxA9o2i+Cd2Yqnc5jtpVfMUGhUEMzUx8zoDhEW9m1AzO80pz+8rFJp6LhWzpDHIfgNvnE3VKpli4
lWGGe3MAwZdHpZeBr93jOb05ER6FUUSy1dBMevWRBMpsi3X4hFfVL/kTAwne2qx6iSkf66j3g4oM
3B14KIbkkHip2P2XwcLYaZyBUeQPAqvrWdH0zy2xAJ6seYZlhlmrftXA4wcg3MR8fZbKxbRuHxKs
tcBOqlqh3FD5qU8BQwYL2yI/x9Ste64dCuaJ0iU2/F8QyQtY1kvpvZDIjEmNOjGrXvV+MUrCe9dm
4d/s05vY+fSacxnjkn3t1q3KuRRCmVvU2SaRSqz1ExRBKSBvTiwQw+8BKBMSdKw0210Uwlvhj/cB
ilJKznENJdF0h0YJemDMo8oMXJvnmqOmEEE8UdDxOLe4rp3ArLfVkzPC9D1q0Hb9Vk3yoVRFJHx5
Fxwh8twOhINjQ7w/okvxCbJU3pXF9seODqXsZ0MkJYhnFuZeUY+frHCyN7jWO+UV5DhAX3IutnN7
LIuqedbeHYNa1dyhmlevNzzIFbPQfFpIj2Ok+GeLXprIOPINWYQJ/c4oMXmROb5O0QQ7D62t8YRu
XMl5prBgv2RVC56AFqpcxgrIlb+zKgfcuAxXuFthMZcNrAjnqxMldu+5YYouJZLCEuGGu4C6eqmG
ePUspANYnxPJC9w39C8OkGXC2GB7H1fSyi+cInQRcdaGdCrBA0PLOBvRnu3Flqfh6OsV+Vj0faqH
44zh07iDVvaBFCgF2tz9mPjX5eo3dOJw0+EoXy/SAyuCBgLJ/WUs2OQyEDgWrJIWROhsG3AdXH4E
7h0n+l8/DbyuIqvVAcbZCPC9gCUtBaxqDWysKplAM2SuTdDJeXRNUQy1V7svE5Cx1jgTTQ8mUPh+
/NErXTzgGNDhBkmoVCQygp9Em70ViD0gBFQNmOiTXU2oaf/XQaPXUD6quRdnlZkZLeqLEKHsGrno
QzZkoJgp9B3P1mlpRIvgkt3iQkP2LrZvPS5G2eggBE67ccBKd07h4MSUjLxtx5JSePtWjs7Tcnm1
xjBgJ+rS2DgPxhMO4u/+nD3IlzLEBolgOPemfXYda9SoYFUeYQy2pohURrDeRCzsO1GTSnVXF0px
+hboTO37VnhZKzEPiu1OyFVuoxgh8Iuy0mF+taaDfCBaZDXKtq1d/d9ylZsCHlFkEJrfV1FcJo+n
Z2/plhREshiTRkiRydK+HHVJUj/PhMek0epZ+ytIbBTaTKx6ZOlm4Ii2ETFMh+HaVr2pJgxjbc34
2jbg9JNckO500RjaPfLZq3SKZMFyMAo3X9+I8xWWFQmdnnvOdtarRN8G86HEnMBUp4EpG3U7EX8z
f2jJv6R+hinGNtjXlVaHf8ESks18wcZGghisyN2+Ft99WwETskzUYyiU052AgBUkxMKog8CpSkTH
EqFgq8c7gOoiwXMvxU4w0Vwth/aKO4O5MxmvAyHVzTEH9Xkz5r62NQeoqxohpkIOlUTP4S03j/08
M8ASHP8xkt256rDtJki+xUnEdEv7VaXTVGNkyDLjZSFh+sQ8W8BY+Q9ybi2rgvbKEIv3u0VoqUHP
Ld8FVQ9ZVaC36yz/KUbZs1nUZmld/ouV8CM1t4/TdtIx/dVwpOsfikZxvZmXxas8sO6TEUiwU5hC
SSuCqTn3XLxgrZ7hSimZwyP8L6DTbBvS+qZu6GP4tSuPctMmWa/DFrPixjxtRZlDrl+Mse3n3DuB
yXpvkhPjIEptZ8X36l+oIHrbsKTOeGz7v/DjYbJ8vDqaZasGgr9B0/Ij67vFf+g2odMoX/pAgNG0
rTWDFMeSc3IRjLowmVcX+rV9U4/h7XHuZs30EfXbyyzG6VGHKMKnlITqihqDU4tSM4gKiNUnt7gt
SzIqHAfCQOKNce6EkA6kvIAdO5u9LjAOb4LFcQpEzGtYm3cUVdjuxPKgh4IoaGKXGURZA9tnL4Mq
pBdL9e9Gr1rm5L+6rG1uw5gMwV/5gWSYMZgUdAFx9yeM/l0h5dBuH7rmOX9j3AzHhVzrMff/knf4
D7p9o4vmFOSOn3+5XJujn+2/8zrd+6urFZWr3TfPIiCyDUZFcnk5CRIX6yWwocdAiKRQCGS45jwH
Dq3u+3xUzrefaHifbdAbHJ68av+enmh0OWu1v4oUfa21L431wZY11EdA9dVjn9vL8kgpSyH4r71y
rnUU7jsT9Vb2f/edNrhsx3xbKXpIkqr38lDLLlnU5++GBic8Av7EhepRMqbp8FakNRDoDgMilrW9
QZ8E215HUMwJQKDYzucSJHFt9mb+B2gTcBRIpyeAMuBFIxk9a8XHLOmU3QLX588OKO1pi/iauYU9
CIdU146+q20q4DBM97QnKHJgUrTbOG9chcGEtCfyhrYZHtj21rSbdg1+jD5ZhtXoAHxA2/1rPBLh
gtAfi4Nql1Vg2N57GavN2Mzp3wDo3rEoAHTndpAsOSBmXg4GYeFs9dpngoKmjqr0lz5f4xF6MxIF
FkcYLxJywTBNX2FhqO/cbzc6lmYkycht4VCMhMq3NaxuXjhsnulIK2I0CVdrgmEMryt9nviQPzfk
d/2WsYanN+UDYsP9932jjmWAuInyg9ln5cYcHrltEXf1dp4oNg18M2FZQpjlo45j5NWlYHd7oANT
YavDERl2G/JPsoVX2XjKGe8w9n28DvG4WApMTn+Ls1FLFKDtCDdemz5JYLmugAnQn41xn/SwZiFz
KCUhS7w2tmlNuYChT2qQVtrjykjdLuj/3xV/Lffn4uELosRe9JujrDHXFGgt8Awz3Or8QxcfMCfa
9c4tIvIDeudQgVfUeUEnBRNG1042iWr6e9S/yiwOlMV7ZbTlHiburg9aOHfYpuspg1rLI8cu2wRE
3cDs84uX9xOhEdqVxbfbgEdwbpjC5eJct6nEXhoL9/NYfRP3F9xWlRlnDbUjfDPBlwQY7GP89u4T
kGn0h6rb0PbAqGgbsnnMs6zm32UdYde0nba0xbItfRBCCeenZjMjiWvibAJepGY6/I3KJbhDaln3
d7A9NfiZTCZOBMvtCXKUBG86Rp/EMIK+CzbwEleDRgTuPaCM5drpT6nfGenLki/rHUUnIKfICkuH
HfuxP719dDdaCWDzuo4kPPo/Dp+BswR2KeNJ+FzPZ7CGCYvkXofxq43oVxVSV7urpD1rD30s5d1k
SYUndpa9bIXpzZuJlDbhvbM8WZaQzEIPUfMf8WXranb6O1g/GaUUOK6sRzQRBUUuyM6y/GwlAREz
In4CuYur0rWWoE2wg+/1TYk1P2KigAWfCD5Lt8MUQTg+MCpDNn75bdlnV83AAxRQirRen8ErUhIl
r+v4ushAlU1B0Y+EzguEgxTFcg2zIMNeUHiIIzbirtkH3nvHi4ViuVDUmlYTUFVxCMEwoiWa4uVn
UvuJ6WtTHmktDl5SfvCXSfpXbzQgSak17ZLxTzP282Brx0+rSxmu21TA4SD915b6AP8TOWuolZir
PS2X03OfwWBWgTIkUV0Obx0x6YMs12bAkbt0l89rbVjxdsESdiJ1mlSnHRypz05JyYt+Oq2ha7mz
rWbtaGnSearQClKmHWM8AsLkE1G0fkyKqqsJEqbSeknSAVEx3BK2Y3IFjMYss9QTUFlx0NXZ9Bo5
nIA0NrAsaTXi3/Q6396RzbUB+5OaqahwuX9hdl7V6hrQFjPq461q5/ykM8YnJRNWfAJ3KNXGao/f
5DYU2H/51/TNwkuNpS19p02iAzEVI68yQq544cSdhbcdRlreNKxakInHY2ovm4nBgXFeUYfaIl34
JSJtudrxQonMC/K5uV0SueQLHT2Pq9uV1ZkpBDpbz+ZqJCHPM3SEpsIVpiNYdUZZh1uPnUFhfwGJ
usnBLSNsWY35kxvP5drJU6udpVVBYFx5UrN7YAsJq/PiE6XNHTjFAQ0YszLTtTfqg32KFOIz6i7Y
ASWFf4ZCyI4YA4NHexuXQl4AtxqePrkOEuR6Zf8K08UnKfNtIFimXHdqA9wsWKgLKJmaj3y2IzDO
oH05k/Ngiq5i2h4E1u/qu5XpswfyYrWfjKdyBs7cjIEwzYPy2q6IPRFjejCQ65LULOBA2cd60Qut
FEbix9lqKsKdanU0LtBBDd/tTAlhx3zjm6yBcoWm6RvZSEwFb73QTX3AhHGBAmFrnzmE9Q/WpbEZ
HHuC1xzSXXBbCQ7qaJA1EDwsPVLuUa5qa2eaO04B4VK/JrvjIfma2GmNOUr6C/Xo/tUyZYctyN3W
TowlS9ZI5bIVWvp7ttzbKTr40vzzbNzgBLQrtxd4tyu1rj7NgHkoAZ4mbewaua9wdjjkmunyuOk3
oyA3er3h4IEImjSLqVl2LMKBRzfa4YwLRuZKGdkCk9EdjivxWgfrpD+fRvRipPMrotKGuKN4rrqc
W/YIdKkJKnv4aXcAiqlaxYuAW8lc3s+p/rOstwg+kNZZ5jzsecSTFsGgMXhnaBeiZuKVcn+zC+0A
uf1/4+R4V84rPimbMdYHq40sq3wI76QeVl7PHD3V3zzhpVhNNOXiXGMPW+FNihEL+3v2aSJ+93C7
aa4X22GTKXCWCDN1e2VtFmwl8J6E168nEHUgR8H0JQVtq+LmwLFILIKbPv5SvO8KxpuHlWX+Dw98
ncwj0jMzSM+tGL0c7bcbaFZ7/CX2OdmCAWcqR1xYnt1zDPdXMjqII2UCfUdJto5p2tmm7vc3HgLC
NZM5MHx9X6iNbF4tHoL7k49WCL/xkR/oHhTrfgFAL3uoLqOd6snst5RZBcMftffYPTR9O2iDF5q7
0XXKw7CRrot9oOOTP4/eIKvnaNf0tfVadYDxwOekgTNRmbWTDuodEyK2FqJOdvkcBZZ8i6oW8fcw
GmFF0yShXyZj3ZC9iUvs7iSb/CT0aiebCfIKQhN4LBsP55h9IkSzlnZmisdGlrV6IZzj70b1A1+m
BNR6GyWzT+6TEehCh0sFvddQePbMnsda0mZvqzhKF0aQDLnyJVPn8XckJkL2t1Vn+FAT490dtwzp
RwnDMTC+T73GTXXT4Sxdl1DmF35gLodNuiEAWopfgZOhqVF+72K7DbdiGO1rCqN1Oo+/mu+qz2Gl
yxVE4rTQzt7DFB7Yp5+hJIs93sRC1//Uy6aFouCJ6N87CVL1Y0CV+iHT28x9i2sjL8kiM1rOJ4X5
xvCW4rv/DWZOCLTN/sFb4zIZM5lCn+AgaN7NBgzo2BgWaJKhEX0EURGkojo+qBTSgtgMb03adxt9
ZAa18x13p2HUbdGSCyYpGhhiWbQoWd1M0wtCBVtsK8TkvVJqs4P8nD8oWRDOCdrR3l/6Z6yaq4oT
cUyW7A9od4izEzcgMegX5NcmvdkZsPv2GI3Mjlbj3EnAm5YzQ/GuoJaK/o3Su9mqOrFDJj5lQQv7
mFgdXWfcDMzHmDrWJ+lB26UbkxvDy+6CTZiyOqfBEW4Fmiz6wY9AvSO65szHWQie0i2mz1HRZ6Tw
xe2vYcnOFyxII4I20CjQPIlxrpCB5NHjCRJWItI+wGK3DeiKcz7lFXyeWRCP7iYF+70HHHD9YKWv
S4qMPZUif/KGV8DZEyDUjXgsu6Xtk0gCwljhUo/zRZB+ODPF71H8U5o+120tetgoPSqQF/Dvfi2H
kuclSdH30xCgVjZ/ST0UXbUazJ9N4/fVQm1Cop35SArYw9+n+pITIR0/q5ylot/5wCDKcQqNZgKs
mj5FXJppk2EJ5M2iwkdcfmtPaYCRh9c5KIbbT45SvsobfIabMmdk96ASvD+pnVDGyAza4U30v9Vp
0HXI2SlMmleItlN8eGJb+0pCIOZkZ1he/RPxfOyqT/KebI/W3QGFckxrHSPXaTuhr+GMrqNgYKCB
NhnR+2Ry/BvnCV8fQZQHqa15f7mupER/euU4ZdTL5BVYSOLpozXE7jtQkv3itCXxgZ2i0ydSFU4G
nN20WLTTiXlAk6xzmNrUXGEuIIeQy6GOQnuod+VbOhwITBu4uxZPxKOonVDkJVYLdhaTuqG7UXR5
yoPhQGiyfTM3aNAaFqgMS6IV3llD6LeC5H5Mw1H01eeuuOOvc1zec1pKwjTr1SWhfQyQqTXfyqgE
QqXa3nUb0At4hd5qDaT8wtzUGPGyrA7EtHvB6/hYN7H+nMjnlwDD+0O8h4ukb+xhAcw+wYBD/T02
1K4OB9Wnytcm7ypPj7VdHNX7aqfEc80Ebeg3FJNF1xNyfSXlJsSejWG91AqyD81HGQA7H87pwUnZ
8pLswdU4OCY+IaiMm52Vt9K2KrqL96gWidelQVski1sX4ziGgiqR45+XELvpUVULZJ7nTsCRQlU3
AA/FatJ961e7qDSDYPp7wV7U7lswqZR68VCfRGGl4rWb6OhAn5+8Rd/A2Uop6at0O3PKhWF/se1+
B9Z3y3Jtnf5STZN6u9cHL+888PdY0xNiUlFH7KKh7WCMU3YdzTy6T3yiJvci4XhmeFIFjW6KsdCL
XzSyjkg5WNSTRQPLO41M5Fh8HT6130j58oowDGfjk5vSa2gKLTkdDLkQy5tZl6G0a2vST2cwTUMv
WKonvSOsqbUGfgPXhk3ZkdzcY6MHLRT500De5OfN0I4HvLoEDDxrcienvYcbyjydpTszMknzHoPp
6uAkMPDtA5Ew/0lTtVZ9VDx9Ym6E5QEY35VRJxkkjsjVhstByFxA+903GzJ7YRlm7nORrQKPYAgi
3YHUjFui08Ip83HBYZRx+UXIZ0ik7TTVkXcJrn68sckzorZpFbNK86qkYyKT3An24uX67Z7WDDgL
0jAswPsA+B9j+W7lFp2fE6i2KYcAK9IVnSo5H1uqhvPj68k4VE/UHMntiHraeJBlZ1PetTU/tAIe
rrpL+LYJF8ikExZP1FqqMARLAffWKQJXSSQUQMDRAEnrOUcLi5shmahWNv3/lBI3gRDe5HE30Biq
OVpmd7Swm5uyoo/uNhg74VWThbnjFmthrgYx5rXmneHR9Mip8upsE9UFOWWiI10Yg3HVa8wKElEk
PwZm2GLgmYM5WbNGBpxo5F6apTGDuShuRVOIIjDQyorcBwkZKtc1VqsGAUNJhe8wZyzYj7mcIC9+
hTfMjFc15PBg4dlRJZMxhPKDM8yPvWxGygTcvRGz9Lwu3/kA/3v0q/BcfQZr7rTLWaJmwcvCNr9d
NtUHFcceDucDRlSmnHKDhQvDu8/stuv6e+mmZyxf+NgriSSyj6p/Tea0oBBMKq/ixP9xiv1uHZQ5
RCOtPDlGoPyGNbsLU4KbPBtDc5Mc3rzdB8u0FEopZjQ+gvBLcjnAIJjrFYez5sHBzLQ24QPiUOZd
vRRn4O3XtD1HjLYHYJMubIkwXS1jpnOXG4ZeJvSUORKueD+McVEIeIDlkKyBxRkvEptHuCOTPJYN
fF8k0DBlpd1jCWz8kXsvk0IpHA2UfKwvUvYS+YOCizYnaUtQ2gAtwXlAjU1YHindgxOGZEIH71My
u1jpLLdr5TZG8c9WXOtHcolYXpqkIgDcfTJtpuh6JBsYeRKwLOCQA2nPENyfkp+/nv4pAOh04bN9
AkcFy6DvaYCK7vEO0yk8oDkeGsj38KA+n8Y6yWmW7hVGSfqOePEZhBNyyqU2zOnNuXqKLDpN5k7L
tw2lwGxE/dQoiaIx0ptWd2trvI5n7Hj9Uq/ASNgY8IPFCkSlVMQrssx5avDXGKXqmoIVIB7ytTn2
silPWxj64QwkZ698/m+3RzCyYQNNLrr2v2w4/keZ9jqcafH8A4rr+W2JA5GYtyy4t9D38/E+ilXW
BJivV75A7SwOPy4lTi1ZEqQ3V+iWqTUA4FHLRBsnahKVNCOl42VT9uBqyiF5UPuihCX4zE/1UBPS
NgC5JVJTcyrTBSM6N4u20LYcaPAXh+Liv6bMe2nRBTctRPcmJ8ZtNC0WIEhhZMO5OoTN89OEo6Gl
jKjwgsH9gnE3o+A4jVPX7u1apPLaZoqLSSdJfUFK9cHw1YZTDjAzxatNb1m7Nqf0w0qWpUt1gORJ
ZpwWS7FEg9fY+GKUl4n6iefCiDZ3Q8m7h3IQIpgZOmwxLnke8o5Cvoc9ttMxSpXk6V0fEl5Izm0j
i3GnHwFn4/n3gjqi/UTajw/RscLHhIn27P6pnzvvaQmEuDlUbFXh0k6TB0jaFqY7s3xS0hXM2T52
P2HVvIDSEJV5Q705rZ0atLsTOZ3gkxoovDVjfepvKj2DR2+NzeljsmGOFBGj1XILt219XsBlSeHU
s1VM/eZG84Lpf91tZhgxFt9wp/0kcaIrBRCUrTCT2zg/1pAoSUHxpAYPKF++L3TLkX5Yb4vXgOPi
k5J3+6E2cbJ3vZBiMDFGjzBn0jbQOu903nTvWTZWvFrPILKMNKCdVlhAbwgL5h+omCiTPhAZAOL+
qPmDJOBH9/zGdkYxASAak+C6TN6xrhkc6BYN40Y0MW2SjHnr0MEeth6ZRsV5SP8WGRS5scybZxBj
22YSnj3uJX4q/nSLPJgUPxFOSxm/9DfjAfqPzyGA0Q2AN08jK50qmXCIp7603hsCpF43iyHu7+Ka
sOohtmSiENZJ5B2iL6iK3iPtx8tzfWJh7npK6Zz1e21As6G88MV+MgTyMJxNgbq2ipE5LMJkPzB2
ns7ntMK72Y+Or/hwo4d9XChLsX/RUuOEosu/lBTIkW1eCGLJT3NSrQr9DWNMLH0teAawP0xXnWnw
wiozo8nIaugPpm0qPF71/azZ8y/iXgmYerw2vmnYbciwn4MvjeQNVubTBp1r1Zn24kWywRpG+m/R
dzNa4YOZa4BJ7gxuyUfWhc6ae1Xac48TR4GYD/8n6YfNAzjUPFCCNM1V5GzzqL3iW5/D2y0PeTae
oVk2zfdG9c33cyxcZwzhL9AvPQeTRJfwuFgaz18/tlkh9l1ha/lxYwPvgXO7SNbHHvZOzH5mIYsd
AuD6TnlO5oVOYcrFYq2LE3cttkVoHDs8LCTJUutlzPpqzdT6ckplS6jsW62N6lC3HpYwUqPu8vHf
K+WbV/zWCKTPtZYH5vuFGL3ScPEBOVFLH5wy13wh08pF2Wq54/kGK59ydcT2SQax4o3Zjd7pFrfZ
o7mHJN6sfa+Thda67qzOQLlLDNcpxLsJb1v9OOWgJFa85IMgLO+Yx0x9AfDppNc9kcVuSVCJ+jse
3LrFwG8U7lmAUzqHZH7JrD9LuoPnfVgwQFlxT9TTgBFrAPFpqh0U/qCUwUMtfe2bnQsAiG5Hobut
cOd2CoFdY79TUPWTIqURAGHAOFZpshXpnv11nuNqWDwnKRCv5gUVq+e9qbtkf3ix6/ADgFHb0ZJ6
32sXeT2Ouf31zgXQI0mOjNuuja+Mb0J8bjv6YehMMpM9CICKlbLHMhBruTrem+OcJBtLhONx8qZa
PE17AwHObNTZFQNc7kjpsJvVM/jP/IpZsJCI3bp4c2s8UpAYgXh+Gd6Qep5Rn0LBfLapKAy1VwWB
NwMyWSWPZWzt34nYoSgG+PbVJIkUpMyZe30vdfaGGg/3oPywGeN4IRWColsR13DIYuoAUxb/kynp
mFVBoM4eUD5YG5esZJ0SFuhHTEeEIAefKKhNa+LqPXS5nGenp5Qis2VY3qtQDJDEFHQawFgrM0fZ
KvysycjxWMBpxX9/yNM77uwQ/jCEiBenOd1VycuE5RBT71z6+pYorABfhhZ4+IiklQnJ9xpMyTLI
KWT02uqWgcixZyCHwYLgagTRW6jQbxrYyRfMfc7NPhkXpyaUQgeODsNs4CQqRaokhI6IFBpbAkDJ
w3Cl8Y2FBr2AjyvrKv5/3SxIP4Q40VuCjgWKzUvTcXpoaytobfvA2hWc2GmUXVfoe1K6AzHQ1Mx7
7QoveL2xR03JXYUiIIl7JtIhoLxYbZJy6dC3kvofMk6tGd6iONuj9WMAeelhX+h64qx5EjbnaVfI
yXdLnx+HWS8IEW8AZwWJsco/LTEpjLTbLw/Xbarxl01Lms94VUDpxqXUqEjbGmGYQWIWdz+I9hCS
y3LVDePWd91z8cInt+HMGmCkNo+82NTFgU/3QoSTBNrvzPYMM/mP5edhCDkMvPJhlxWKEwxv6cvE
N46EvA9oUcWFmWnBOK0NTxtcspl5RFphkOun/PmiLqPSh1QELvmlVO5AmlCfIX7GGpobhsc0W7BL
GVRQRYyXRHXX+1yJ8utnDKxA6lh76e1AhNDQSaOvp6ciaUOueCsCSAtJmJ7pyKCbvtycgtU+9r3p
uj38raDIxvfn2D53dwQRZUqX9JNI6ycIKE7cpi13RTqi7n2bIK9F8dnwRcIvYeR+8goANrAOJfYD
vKdCnaBhTljU/seHraWtGYG2b6FbQbxnmvq0D/oBd0kREZ2H8wahs11CKTgO3TdbesUg21VbjAE5
QZv45UM8QQkFXBpDpzr6oHJ9ksKzIy5DywDH/Y7puxpnEyCdrxVSmn2FYeKEeDCXdx9o6Mk50Trd
KZkDDP524dx3N4qLa9CXTVsndN240ZpAOy77VoKdFQrFQlh1qGLUvPH8cUugTJbhB1xKm4jLGUYw
Xf1+sFg20aNUHDItmh7x0woLP9lQ7wkXJ23nDIMyjFVHz91v4QYnhfwyl4x8/JKybUi2bPk52+j1
JMWlLtDXhttR2O8rdnh9s7CJk8yDp6NnzoIBUqoAdJHmMomq5h0skHvlfaatKae20im4/TIVip3R
uV/egz+Gac3KMch2SylHvaiCzq0S/thanO9txcBa40a/LwuYMjxQeKtxI4oNXTg4P310Pi6DRCzP
Xz8eRX9LvvL4BnKeJ0Gwr2LAucOHy97X/Y5PFdVhNetMjYrMOWXmkq8hNNOw8B1txx+nja2Ei9ZN
HebagiDAsruelFW23+g4lFhSMX7gHDOtJTMsy/cgBb7l4G7+i5QgLdOxzXwPYqIuF18VWL3zloR5
QI9dMXIFOJnTRxSdJHal0QhTwNz2yM/pPxb/itBQuLEKub+ti8Gs0YhX8hAPdKIk6WvdfmgZbnDD
NIXjNpGFaW9qWy85USZJfVz+JyPveE+lDpaipFrThceRIqdyK0tU8xRFsRjcc6k8/6noYZcW1Ofq
DsWuxdiQSKAowND3gMGsobbKebiS6s9uWwGbPtiA0uaFiFFctUxqez5e8Bt9Gm6SixFXuCuCW5UW
2+EPdtYspVl7VLvqESZGA0TUxU4WSGegClk7vUEUfH4k3zQ5U3uG0y5Zs3xUb70XK9Ff2PE2QBr6
ow8OlRA+dZB3Nlhuy6k8QRdAA/MOS2VaBYgEJYqHg9rm6OCOF2sZYRFL4hlPRIrw1EsdCGof/Bc1
2MrDBGC/Be3LDC5fzmUn92gPwMGOLerQ2BykiGh+1DEHsOHDotvSD9sGeHv4NVaQL6cyubpKvQfA
ZE6CncBD2yeGDEn97Ao4GksX857BlXDzssceWREJj76O/z+7i/CxyDYWm+vAGWa+bY707KDLADBR
Fw7WE7ieWo+SsN7TpXIq3lL32VHahXNdI3HjirjxGW8zEutMwD1BSuAfrfg3X2QVLi29Uz88D/DA
QoQtaAu8Isc6crcOjRKwVqeZtiJ4Y86n9d0mBiWzxSJzLKFyhZx6/ni2DPazkRkAHrNmSit+0+2C
1Un41J8Kw+mxkyQI/SxUp1U71/+zUghGx3xuAkqUL+yX4anBQx1IqqkxExe6gaLw+3cZE8OYDSST
dKKm2FEbzMes3AqvcVsQYyHNYcJ7eUhRtYE0zh1x3OsrzvH5iY+scFMEhl7CO+sKei73ymaUhnwI
hoabFsPIV+UOhA2o6E0eyor8qCBv5PuG/ScPuXmTeWpe6QKfl9EQDv7SQXE4ykBCg01QEQVcCeyC
7fK8USBPrszcO3R4L2JQW5Wuum8TkONd2Sljq01Sskxp0uYZVUEVlI5KyJaWRznMP+mCnfmDM/po
0zHvQMtp8+mABI0PVxhz517BIFLVBowTCK3EricCDOqBDrq/b38kEgkDWohnXEghF8RSq9hbdRMH
/WhJOroJdq3bUb+tuLfKpOl6+sAchuWrE7lxLfO/anGfk1xwWCV2auKheYDW/tIx5jwJN+1LZK5Y
14y6wl9jAUVEluY28Ol7h/D9CHe4zpZ4h4VYRMCaBUgmUxvnR1/+2fpmYl+nTdZDGot44mX2ERvS
Rc8Ui++Pz5HoUzjGysxQz1sCqvRKI2hBq0wfxf1bl3udJNFvtPDia2HrzrBtWCFMYz0l3Rbk0ZmH
xYT2pnhbVNWY6dEF9Nmyma5o+R71Gz3szWsCAxAdvISEisTLD7LyMRZplG8CqU/GKM86XCRUsImd
Wf3rz1eYydq9Hf6loEQcnps+HJXn84DKDE/ixUzXu5f3N/q1Asritx+Tvy8q+8GP7OiloRA3fUjo
HihdBmccnY18C9164p/RLl+cIQ88NW8nAwRO81CU09YlChNyvfjSvtJv+89JvDbgyU/7MAk2s362
gKYCBcCRQZWgFbaAe0p9IAij891frbYB7wVC3D42nrGTUqJZdwxaqpWFIsWikqzcYnrvWB85SddL
bItMQctFiWBPwUOVDdmabkLs8faVKHObodt9lb73/vc6QVy8O0R5ohXnb56kXt6NuagIl9IONRLf
WAm8Ul0pU+uIp6jNQv5fn2zaFKdAr5s3DeuOeVl6dc8/RbqKlYJPpvboJ82vDrzjn1UfweUiK/di
pDG192JDYVSjNx+GfvdyCwkUTKQVeEI3iaUSzwLwzdAXT5B55QU+h6BuWBrWihdeBKlv8gLc6ejf
D2DzE00WaMHqH5WrfFDjITT/W4GcR+VbUphK01+CBqqtWqcYdnxJh8pcl9sBsXv7IPhoxlNIAPUG
+Sjqp99HQeqjuqymVtIEpkU3V0+fWrxWXUqzCRV0kcPzeXsl6h71zvyBAdN+hecCE16wSMQ4mS3/
kw1Ky9vl4crnTYtfAbgwtIMvHr7VYTOWDOC4M+RpTgeawcf4dSwR4mX18zad5F9OcbYx3GXqVF+0
NgwIRCG4r04c/HavOWCinYKO8M126JmuGQRgd0Llb0BemquEBWAdK9bmmM2u3s3Tm5F9rIEUYNah
OGV6NU5dfGcLknk5vhOiZVXQ5e7SVccKvzkWV4/tGI7pEtt62Q534BANpdxY50rGTvb32U2m4qzJ
BdJcbUWGXQPFEYYGyFZTSt4Sn5XrcplwZtm2qOJTl5Pc0EAdNOw9fGweOvEmKxLJRwX33DtJkUOI
Ip5wu5jSBOw+jKKTnMIp5RL2ilQXrL10PZm6KKW8g7n9PdVM7qt6DWhb3Hvgm0w2zF6UH7bpFtRP
TmGGBAZygR3/F9aYVvm7lENW31vF85kjA8zSvNgHqx5Uc15kALyi3DSnIQyLWKIENqZ/lrbLJJ7o
CP3wIBCaFkEJOf1sZEhB5hbSQpW+rXo5snTg10XCBG4bLXUVsWy7DwkM2ewgd8VulWCgF8PErb4o
q0CSGy+5kb3COyQI4i2PoiphFzvd2DUXNb0yqLZaXryL+hu7xxpV0RO1vEs7fmOPmx0fr2da40ut
cvdVnxE3u1xyhuWQQrcQQofg/0yJANRc+gLv7e/UnM8Zgs4xFlOp4IzIpHpM1s0L3wQiNpW6LXZs
0RUPJjv/xy/JOx8477iDPfLQiQxAoN70t9iF5K24KtRsQ/T3J0Nezr7LnWIk4owsewKGUfw9rMQ3
RaKg67bLskuTRDJ1Bv4tJt8i9OTpZYI1OEMnOwnH2O3DZKWNhFdSyEX3SMSJvU641JFJastyRLt8
WWzkfu88UlRt/A7imAM8wxfLTQuQoQ59o88RJk55iL1S6gcsC5DHg8Z4yjpycQ0HhlA9J9sixlBB
sowzJ8uEaYa7R5xLNiulYeAKtHv4edD7QJp7vPD79T0/dameK71S0x2+socFO2DF8qtF6kXBrUf/
VAd9DXjUhs1k9WfbDXWW69Ee5X7vfxzwVdx72jLIJw0+6agzn62xAZf/W+8lrMC1rvlPrlJocLMH
SNirrr68pVNhSyUthCqHVWA14poE8x07XjQEpXFnZRdPm7jJo06W6wIdi8ZRX3GcDRqprBnUysj4
0F0YGbkk44NKao3G6sbyhifHH9+vODNbjbrMXaEzXiHKdcngOqxv04RZBhuePnuFyAApinZhtib+
vcPGWj8k+UaVJ7QOdGMayldaNM3adBXt/lMFiKuSYkoPXNbQPUo/q0mjnuRqGO+JFfaEw6Y/JPcR
KEiGHGi9o/U2neGeAsSswWAG4+S5FcFT9X5jD53h0Ea734/kRyMBOznigJWvQC6UZ9K0Gplz/vq9
Hd5bsPtRxvnYWbMvYhANsEfSS+6snfFClYLD6qdFh0BYVjAWJfVAZ71ejonUed8hHuJRasyRUjid
bgrXv9yQA7wDQroMgpABIE5qGSKqn4fWY/+41ji/p+LbFD1MVeFiOhW7h6WgUAk0YV4zQ4TZwg7m
zUTua+Jqd5xoqxpNV4Gi746BRxwRw7tvfbqeNWHXIkaPH+g/0pyCqXhK3N0dSs0XlZySecarwTfK
qenAJnQKQg/LEAS6QYqeo2oF4W9IrgFJjiak+V/m23joJYyTw9Zs0FyVk61LnT3U/yPMmMLPR+8w
43jctU04NP+CIB6bRMJRuvoPpjC9JYuyBl7XUSElyu1wJGgOOXPbWMJvemgzF8qcC/oKj+1WPP0a
dhwaZj30IRiIcg/xbwCLs1Quh284qtTpGTe/3FKFHa/75vbZB7sQdgaGiVJenTkfbVZfIJzHBRsJ
tFJDjNqeHnjj6eIopt5WCaEkjZ1f0Lkydf498I18+IUvBHNkN4TUIkdaQKaNUnXpGm4Fw/xfktNj
HwNRL9ChDep2nrNqNSIyGC+oy72Zvt+7Uj9EQdEY9+g2lOj/JfMI2ClhnAUAZBrxRyxJRC4CSSSh
fA5eSbF8VO6wFvyh9yX7pgyYPlrMupw29JpRiiBCh3vEJ3zFVgDbBQWwX6gotei3ipeNsNmmGGYr
ZxAYAzv8aOZtXo3ZZKIxP6d6vJmpEHz+XqtFNFm/iNliHrg9Bo60K4lOp0dcKmp5QFTyvLQc98Lj
/jTRzUnGptf8yuvT4zabu7KquRdpJUK2WkpptkOeK0y/OSp/Fc/hbq0JjKNvHvBreBNoUN7PBgrv
Z+LkQ6FNnF06c66fZEJBmaJ/M09IfmGTHLqroWbsICRnUzET3jTiVc+jZSOZpqJoeixmNmgBpEZY
0oGpajN9IW7NgNa39MCOj20XonLhmT8k/P70ya8LWxaC3I/nTML/7nrje75PYJsnxyqLfK3QH2Z2
VmzWAzG03Yauv/hNtmb2SC6ytEDha0JnPSgeiQ0FXMwDN9zl5rqdQp3Fsa1KEouJ5knkP2o1zxLo
1D5wNL6QD/3DESQdAw8rSgYoH1Y9YxC4bOEPnXtBwKbCwjKHLdXZuDvI+wOCFJBoIW5sfG6N4zTc
9t9HM9U1awwPkBpX5nuHkD1JVJ++bv8c17CwCgbfHJYO3oh+zzJuRTNJHhIf4FhtsCcG5lLs6h3J
djvkMl03Or0fho9de0Ik5OJ3gxctxVOkHEdL6HsYmPvVaGgaBXyYLoxH3niRF/pGLNKVNZ55d92W
sBfdfPq8IBkTE+uIOHEUlxSURYFN/GeVknZmXY0XOscauBmkdBP5KoxRsGXdIfr4xo+VgGj7STP7
mrzQh9jRhhK2W6t4fitP5myR+xPWoSTZVnlVDJOLg+T6JZQalQYDkxEWALXmaWJ8z+ZkyBwVLZG/
cwKBfJQzjjQN0iglLA4nfavOt9XpLO7a1uY6eBWZsuHzWX7HRgh6V4LFwHjkcF5sFTZeyBZm/rtO
JCIA2KnA7GXFQB/np2Zou0kRXq5STtsdrMjhNqMljM7ffw7xnM58qN1Fue9nXuuEKkyVDPi9tnnI
xrSDosh5pva80fSB3fEMsDZ0G6/7skKMZSfY/8tks/FjKuOKWxswavh39cVeUjOiK/wEGl7bCyB5
TQ5/P7yFZfcDV3rIzrFN7U+gNTRlauQOvmR3xxuFuRi0TSerkAUZyUMdO9b60axq8f4F/dXBuhjO
pgWx9sM2D+qqMS/a6kNROwWMfIElU1JajJuVK/vnZwkMe0+r/9/0y1+jKR8jK+VK4Q05HIkOXe9R
TXL29gKULk02eBAt0sk/5CUTy+W14vbZqvscCyKz98Fp0+WxkOutpqvCJaBDn/vGt/vSCgH8qJnk
IspxogHTP5eN4GYAeVFM2wrf40uHJsSPa6ZvbeItkbCHEJj9kvj8r55SWFLX8Z1FVEW5+WSJUWWj
pvqF4spfs7hrVE/ANh6m07kqaQMn+RNsu3ISR7lgCynYTjRUAzIQv5E1v6ecd+Z8OpuI74XjKmCs
aizjMqcLCGr7n/pvtYncZzqQpMYqCcu7zM6HvyOdNwNm5DRhGcTfTL7Yi/XZGYZo52ZDo9dU1MHv
uwzwUpFmSPuXu6FGXkU6bW1SEfhb9xtnFJm++bJj2xLiaEk5pnALKmL6aXlfuXoccELgI8s0V9Yx
u9I2qE2gDvb0YlyMffC2ApwWmsbSEZorq/azDgMfIdKq7SLeVsemkgXZ/k6GLjH1p4kqWPJ2ryqD
LD1UBWr2wPjzRaxeGkvkDDSYY8nWg/YPk2WVBFFOLryT3rbpiSBZKA49zxaBKmxTEvB7M3XwD9hs
oc87RUukBI0vm1HuTtIWBPlNAGNKEp3Xm70HftK8QkNqIeYK2aJtComqAGRj7wojPOqD8Op3J4fi
+1uhHnvSc1Tsqk1yw0fium1PYDGxnSaj0vSum/1rI02gaaWQeIM58xuiOVK3EtLa/wrU3gQf8zh5
2QyeUX+yajaV0LGmx1kkg/r8H179DAO49aPOau9wo+PfBidF5bZgNaqwDHYzwVdE/GyiBZJdX3p4
/nDvXpXXEoaHzcYVN1ZOJduz39wZOA+M4DdyxbUZOyTSwil3Doa7Bhtdrq128pZnebAR9rqM7FU7
c5aI4LvWp3hQeGy3ap56O56KJ/ev5uvSxh8oBkeAD5nEuwMNxr2Mguhy59oByYnHT/VAlc5U2oGQ
osUF4WNHAzLwH+0mbeUbzySyBpL8fO5QU8EPtiSZOKm+0WihqhV+RI4KjMQl7OJ+GGJhiHwDZeB/
p+1L569kB7Z4AICIoWZvPCgCFUpQ5Cua49Z6gGzBTNOYBWbB+UcBu+3LtZGImqWM+VahW3T23jrH
dN9bHx94RYJ+f8RS0WZ79WayslZ58rbUz6vgozT+BE9xhZ/LwDoaYQpyl+9dIDqmjyk636uTgJxm
r9wzI8Mffyr+BlUfQqY3N5wSpRXC9VdJuWo9ui7D+s7UjmiUgdaKYoZMCalRq98fU0NESm21rOBP
d2sdpAOJoqVzr8IoMYlLX/LvcOxR61Qj1nikAXa+5RGRnvBi5X3lBG+/O/tHj+Uq8uYbFetv7GrI
KueazfObih2L6htdIm1Vchxk+lu1ET+m9o2/FZcjDkhCnxupvUSUZISrjsbOhxWCF9n2DMK4ZtQ/
pJfr2gWGDeouFNhEcsyJvQRRu6U5jvKWLUMp02vPSoI28yE1nWQbhxWvEYkf2O0Rawdkqzca0ND+
jXTta41c6tfogfeIb3/RaHgtUUrZmDw0edJaCNPvvxgMkUiu09xdw3LQWHI/iqln61/PQonPi1RE
rJJOeIMBe4IHVUgOZzF7LhbPZAiTm6ssIq8VEjpOeoApga0IJ7JH+JxUMwBmcCwxStW4Q5xIcuVd
meGTbDkGTU+DSnDLMW3DxQNWGJYi/CNbmBXJz2E0NNDaQ+0yEzZSmpKm1CITpqA6x5VyXCi26FaN
JmA0F3lnMHxXsRoS7DqL2gmSXOir7Ywks4rZFg+U023HAz8H1Iik8/GErg5kJuyZ+d6ANd4fy3iy
tNihu+f5B5mVk/E2eajNPAupyytiiYzEyKT/XNIfW6XTuAumajM5hR9Cot4N90VBpjI5HX5VaAFH
S28armDTxcdN3G+F1+BAxLg1OrBhenzUTwa0iDOi/H6BkWnmpH7FxOjWBO0b8srw7dPJY/4Tl/Vw
n4tzDqjJPOOdNI0VyrVWx1eDote2IJx1lHPf3ues9sWSPJUyB29hBCzZFx39L8qSVHaI0lGODpKR
76E8nGIPzYFOEwpVGsOIsGFd2qGTBPi0MWauxW+38znMpMioSyMk//OkGGR7/hNdFW4iygTBctNH
qC8+YNeSQez/3/qncPWR9ElijklaDUQ1C8HrP2x5a/TuaL8nORXa72FpXWrvyOnX3Bjz7DCBsFp9
8mVRByePuYZHJ9CFEA==
`pragma protect end_protected

// 
