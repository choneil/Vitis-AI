/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2021_07", key_method = "rsa", key_block
NtAd9OZUX95s/dSCRNODTF9HgTWl+h4DTOkNb9Y3Ju8T8NsGbsgq1H0S/UY/ncbohmCQIVToM89N
haVItze+LvwnwYWnQsvE2QE3wSn2vHQBgtpF75htH3YYukKxaf+OWkteqlivrrYC67CenOg2L+F2
eDqr7yjC6pMxu4Ko0VI7zbm7JD6T/YF2iCb7EOvSaTDEVWZY68mzTG9bIUY0qZtjz6l6XTv3Quxt
aEodQdzA5VK7AI0QwWxXrcBvzCCG0Z+LBrGFhpzsF4KSwOHU+jRAu6uIF9Mtk7xllqFcpU95pCXa
f9sqX/ti/taMnyqGQUTUL6eUBij3vlT7VnLfBQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="QVR4QZEDqi0w5f9eyB33tNffNvNEl48tInsLa5sl0gI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 6032)
`pragma protect data_block
Mffvdu9pcmgNJk6bmxz8vU18PDZ83HTKZ2SnH3ElTrQQg90g/wweUWow2CetYE+JSkwOoLksx5Gp
dB93hH7iUQRgW4jnZ+YP6kK/r0qmDmsEBirQDTYAW+p3YsJIVvgzoWcFcszK7ZeLOgskXD3BwsuN
GYApBhvBqvaEy09+TmdbcgdMaxUbU06SKSPKeryw6vs9dk4DZKfe/tpfVcz4Kb0NrzGmlt19B2bl
ROL5CxRwuHl8VqRxKJw0FRyxBLk0sKVAGV8BaVn1ecGFouYwBcYLbIeNpyBjXvYbOtHcqMqeZju8
OBDY+7m2ZVZ2qzPI3aTKQuj4fzxh9NilkAR8JG+vFSxJEZT7sHvk5J8jPusRYRpDR0sklb734Wza
KbBv7QWHdEAf1dHYhNzuQ/6nePLwMzEKn3jfnMaC4LdHMcQ57mb4tl/PGaW5DqmJpMeY3+c5mM6N
Vmw/KQFhn0juxvFZ7ZkSdIxFQa4ACo2vPsmG/336UaU7ucuELxswio3tFtF35CTBobcpEUfGfgL8
kJCb1hXPkwOlje1vykREaswVlPTknvsWWpwVLjRVK0VL2VkXWnO8cPYRDulGeQaHQRAjP2YPu4Vx
/ncxWdrx02NkMJLP7wgj36QrrhE3IJhpEsyBx8GBvf6irDjHRcUJd5qhfNtN2IhJ4DK+GEHmRxkz
lTrTGvV82e4v/MHSgmt92NVngrGpsLQzK3JuweNgVbaCWluRdtD+aXly8FPNSAcWAcB+9j4JBJi1
NlDBMoIwVyPquUbtdJ1nkWVg/mB09OEZ+z/0uz0qg/t4KtUzh3L/fksU9q7kycsL9QzGudba3ldj
ZMFvJhp1slizQvI/WAmFAj/8SDrc7iLKMjeYeGnKGu+S5zg0S92B+lQZRjm0wP2tlKE+iWVNiGX0
TMT1/t3c06G0J8K/Zw+G+Ui1+UtZMarohXAN4RgRGrxljc+NS3+43Ogun0wSdEC8ebUHHzeL9Zq2
/AF0+6vg0HZuroolGY/+dVPwAnpOSrL58+jMUJSPwTydrQki8HNUS0mlWiKPyk6u2mq6HUH+Dt3O
sYR1sqoz+yCydD0y3JX8486QD70xag45DLHKvRn1ZeGgS3AjgT8xCAqIoskeNDGkCJOYQZC+Rtb/
dX+ZIqPUxNghMHUyGJJkI02iHwUuZsTBzwR1MtQ07VjpozRfhmuYWGBXZLrpOYb5+LICHHj63/zH
lU8XLrF7Y2jPEAF+B50qrSd+6oAFTlulLgY4uygCrSz2Hb0kXAVzFPyXVMMHMwCkbasn0ucdac81
f3b8ESVmvM0ZQl6y8+jZnEASz7oVJTYpy3/GndTXuDoqu+mTrQOwnCKQrydjSqli5zZDwLw+00Ws
9r7G6Gn1pO4Buuub4DKC1jE6tJF8Bu1Vovptp4wP4ByjYqQ446y1YdU1KabUBP5CX7g/DYYB8XRE
h7vXBc53Ax5QkeGbb9pIaaqdLO9+DSp0aibE+JvG6YpUw21UPkCn4kNiVrBlWPsm17QXFehpkHw7
xlo3QxybatYsqxiDv37iGEI9/OPLS3oqVOWZKFVO3duMEraR+tKZgHKOuxbE1cGxdpbYRJa1jc8E
XoPlxwewjiEqfGekNV4W2vCdHRJMywZfqDUVnv9M7NSmzpRPQJPORKf4C5lbz3cJoeIJnn9cMTFs
9I1T1jc/vhHdLE1oJ2o4ALR6HvgaEDa4yQytXQtIfoammx7pQ31XiAAFI5oS14m5+bp6N31i9dsB
KpdLEXodaF/aCVyRGfyHbP7bSNHHCV8gXnzGU4niOX8XKkt5dXIAmc6jGfsNhCsqnp0Uqt77oynD
pmxeQwAzx3WK8kBCS2Lj/6D+ngjG1AocOIOPEjcQ+dV78CW/4NCjRrqf+qSrLG72UtgC3qXX6KSU
9iHrKUIETWCF2NiQMiY6XSO1jTWMXn7dQY0FbxDQl9lMU2jyuPHirZIiEchK1bv/c9ebiH4bZNHi
Zk/7jGIbqQ3zY0O1WxV99yJiZGMwRRov5fIhvm1vKlmeUaRvV//7KFZpsysSSbiesrh1h9bNXELY
SpqFQOD3FtV2Oy0ZN+5EiGo0dahfy23WoLM7PppBhMLT8WIdtX+iW2vNw7rODhBO9y5br8tyQfUP
d5x6JXI+N7yYzGqOmQ2Cg7Vfam0e/o11YH8bupbk93YbLcGlxliwTmg+pMOU6D83kZThs7qcpJAw
sNea5oU6edFqwZcoNNHKl/54g59ktPCzl3bHF9z++dgeDeZgl+OKsLsNCe+jINHPcXEViZrLHlpF
H5D9j7RvrKFQ8iYk/b9ngnycWYFXCPHzgacpv24ufI7+Th5xLDlNOyRztnYKKO7Gt5gfKvJyQsc1
H32518MS9Qr4+r4wFt8iZQcmolIvpcTAT8OjhsaHvvXLNuoGP5FdBajCma0TL7iUtQ29pzv6ndQ2
CMfBdp2h0M5exyvZ+qdAZ5pB6JjOm5AJb8FtrgIW5mTImKUWH71aOH1x8lnKJBqvVp49/WZRJe7c
ybmYF6zligncooFC27imxRE0SGsbUQCW1Sls+YIBPIXhUtzapa3cPTSk40em8fGkTaNE3OdQv3p1
gMrBmBetzYwHmhC/jGM5AcBLzi/gFFszJYfbnP2TJRvZTV/zAC6tAgNGfJY2+ecQ1eNuMcdtCvR1
0ficbA2QRnQqIyv9sfTriTLAi7pqjaGWfcTPzFKcaDb5eu81otQyZOQ1mO9PMQMhagjtGe/zEnbr
cDHAu/Yz+Fy2SRcxae1S4E/UHyBe/rGN4bYz0X9L7Vb/pRq7yicGoisY4NG12z13EJOliLPvCPmd
HtvTQvpyj3Wkb42gMReJm3Kj8V/r/3qYUr1YHW5io9hWsy2zbwLIPAz1blnt6otpwuI/SNfubIjy
5GVxjeRvP4QqUXvoYdiwA+5C8gMyOgDf7l6OFJXHskQdZT5COLwt3HIrGauJ+3q3x4Uh888J+SjG
h7nHz3bAYJbOPAHED8UOte8kjyJFlfL9hyGLYMRBrVuebNS/9y6th2t5cOz0qVl1NR1rcj1yWXVi
DY7eGcKZxTX9El6TZ6kS42leEm0O+2peUif2SIC94PoPJI781627pKWDIauuZz5LoQN+yZv+sUQd
ArN7tNr2rFiLLBHP0y5vKG0iIWQlmKymuQA98hMbWgpM2KLygibdnX20LeJZitPbxWVRH63Mb0aC
cvjd4CpO8MBBurW6G/QMQt0MEhnE7sCfH6Ni+8Wwy6zpfKFoprQeAyeoMHVkyMOrYCvK6A/BuVcV
/At0GaJ609TAyolQQX5kSpuKBkINk11KFRrGWya4Oq5BaYKa9++aXMYfiIhWzd6AgCVpuB9wIXwL
2qeogjhWCUJfR9xyZNLX7kdMdnCFBNoDaYw+x7shlaJCM8m2aMvE0Y6kFaWN1WEsjfFE2YMz1CUF
ntgiwK9MCPs0vny7OiU3Y9ul2cjkM/eiDZTD7hxnYa4+6dhC1O2z+7xSF9sTZo/RrBfINTuNlrV8
T/5oa5tUzqcv/x8YWlco3pAhZIBlzAov6eBpqJkaWUMx0ifP4thwjmg2Iph6FHopB6YqNgy7gJbC
3Rb8RQsuU4LYysZWckaxGT04TGwWvjACvJrRcb7nfyTaxy5r8PQQ+9A1xwhLkkN/wF+rPzjEbq7g
YwWwIdSDezBWfWSv4DOjZvZc6LK2Ajwng9R/ZzCgdYN8JD8/diHpn2aBO+/aogZEVwdSJiH65ws5
ytO+2bUirEhhk5ob4mueF9eMeZgs9RMvhugEaTtes54E6dQ1OpkUAzjdNERGXU59mXNbW6vaGAn6
Qo+uJhPDUSOunjqttFVPS1f3rgQSJs91tBVICl3UlwL95zhEh8KGKXyfOkGlDxlbDA0gSFFyArPU
7LFZtwbW3NAAwz7tQbzZujqPm3uIlrrusdembkUa2UfvE5ZOFyjkJeDP080nYSzU5eRWv+k2uuhC
guNc9qQdj2zKYqW+pJ8NOd7fK+0YT+whtkcYbkj7Wjekcz1J6sF+oxSZX4gFBFT+C1H9SRmrlVzA
qhnvh+vTl1pyKDeFUFJMiUCZLWpXe0WiIsYyF+V5t7mdOYT2E/JJUp0s2pF5auRGRxC3cuIS6lHv
1wx25K6PqB5QznMXZlxO7OVbPLVGL4fNAdj5gr/WyujpwYrPEQRflXLOKmpl0QrWM0H9VbkTRviq
sVCyzoaPmmmZpLFGjY7QX8Lk2+7pcI9SJhkzfvETQGzbBjyH3umMc0bivUmN9KvSJZgJgXJ4Dv+s
u4CWS4syuydQuazeqWnx/H3sQAbhIkUFj/5Pl/JX62ZrWPnIXvYMPnqvym8hP9AyBJF7o+paZmkd
5YIRmSa7Txg4kY0G/LSPwH29iQ7/YrkTjKO/OeTUZ6wKLVaNntcjQD6fHW5rLYKVpXKGyv/KAD7I
H/zsJ6NF9cLkAYH71roBt2LHiHniW63DJpFRgZ20fQpaCTKS+068PtkMfFAvjuqrcomv9rtIUkJO
pc6fAaTI5FOj0C08jy0HixxDC1f7bBCaTIT4jDGRrbTvz/gCCrmnQThVHqTMdtmK81Nsa+Ehw4N2
9h0E/MdxSA4jpWPvwgFSozWcF3UjNuB1rQTGYKojczRcb0omJnvuxeI89VhbhXfNW+CAk2INzAeE
RYAalIjYadHdroJZwp6zxTKZkZ9/rEhqIYmJ21KUTubWMc+jL5AM59lhrCA6uZ/NZj13DJ794/Yc
M+7BiBvXAgtLWv2gIhHHg9F+OTVrbd5PQrkuqJ7HK2lwXqZTZK6u/5eSxnp15o9oSdL/ceCHAgGd
CPw3IoelWCZbZXBwrM2CwFiausgzECOXNdU/jVHBcn0eBfGlVwvOiRU9PQuyhvn+4tyNZaowtj3a
ItS7oYA3e2FnuDHy2PRD5k8W01YdDp+u584a0QioxS+Kjfp+WU8VZv5mC69HO6eB6kYVatG95HOO
RN18GUxyjf0U2Yrigr42Yz8vZX458dlPhdp8n3CxrdwrK1PYESD/2Rx3gfhRB1P3yK+yee3vwE7G
BzzuhJiK8QgjRKCpv4xF8km2jbHpBeEq4emE6yNricmL+Ojn3ZclKu9DEGzqlC+1+1eYj+lAgisl
0NfJVPyvUzKArmEVC13/9riik8ysTxaIUm3mRd1K3903BmnTdHFwdkv9hVEz/GFmbFfUueHb446h
Svpv/xm+TYNiZ4q0P73vFQBOQj4HEoskrzzT0trNQWs9a4ncZ5/LxJIae3s3N9WwsFUmIi5CJKl+
428o/6j/ueLDaWbtDvx0m6jWELbD47P9mesntBVbYpRkKsag1v1PihMHZoEMrH7Kq9CqRBbH1raa
xyL2qmd/f4cY6CDEm8P/h0RMj5oaiU0WjvJdRwnhE6M5YzlTKDqQeZorZ4OyDLB5lurGZWkYPe9y
pjSaWaBCss2vystIE+nR+xK7srMIWnCOo0plmcImi5YYd1RsQ0UeQKnDz2fVnyENjfeekizG6F8A
p9HT2besY8ffN8HE4bceDOaqss6B1/nQAWiISfexgNithLcmfUrqKs0ZHlieTN5UBHAyCsrHKEAb
roytj1vG9fdiZFx7ft3cG2qS/sg2hWHr3B75QrzWrEAZEuSnkJM3bsjYvgymwKXbRLtj9o7yOAv0
u9XyG0nOeTMhzDxQ77e0EtihYCVJcj5liKCQhhEBsx0Ab4d67tkuo8Pw6lrLOXHedOdO2dS3yaEC
MafCyV0n8XwOUmC5kg3pj83vQ54F4KCIJnrwuoJtqFrZ92FZkYUs66C91oYuNvDD2qlfVzow91Og
I74UEHW/rTh2O3l6RgDX/qCkKe5t6cfq04xd3UcLqNNHWUm9IWI0lUtq4ObNwTBCzzgXrEdsq9Zr
yV4AguY0rJaQM+tTKtG9G97m+tu4tQVQPlCZufCfEYrUpNbmJyylb8VoRg+RrX4xR+jryo974oXq
P83JCr2JV1h5ejy+h6TYb6ipw82L4UMdNYJRE7Rwh2Z/IgOHAQK+I3vOMw19PRlJBPWRftRt9mw9
HdZ8V4BjNKnvy2ANinT0xgHV4g4bAWN76N/77ngY5C98qLV10ItrQVE4WPyert1/24irDt6hpll5
64tVSTq9jpirzjqNk1/WXCRtzwmvth4VjxBmJejpZei/KkEwNrXJV1YjRicn9WCYHONlHUShec3+
ZVEvHhojArEzAgD/WkwM1OqK9w3swzZb3bOjOCb2h3NcpSdPmxsH8dXyksYXBjWM/masQ3k/06/T
8o5ukL8um4i9jLQf2OpWVU5YjpxE+aP0i7HluAxjRY77mDm36OIQI1izFodvvr1usiHofsPYM6DK
nRjNifcZx59sSPQuXcoS/CeE0QdyMVmS5OUv4PQUrpxP4tR8ILVs7W2moClsn940e5poGLlLs+TJ
/ZZ6Ty4F++U+wGp7spB6fYC3wTf8fU5iBRympSZUc6o0WAz+Rt5tfJyviNpvGhoqsDRWdG+BFKFA
SSen+eaPCDe7JsK9aE6e3tboia3eFXAPS+630jDqy+ELxHaMLhRnoWXyXYReScuzkqLoHJRFeVGg
F80kT08wxw/3JdbVuSWXsvczKZSIAOf2immzVfJHo/qKHWFszYiQkvLKNMLslkAgS9nUb2KmvBg4
dwTtrLALWLpHarnx1ki+0sfsDpyIUjvfwceFM3xb0tCvc2R7pqI7OfwSAEPbyDEyJYNLmR9O3QuR
lJazEaSULJQU385HcyuXvCMvhNYeIdlamA8tK0Elc/lHTOH3y9RrtWngMHrcgIp4Bk1aBcywSFO/
f4HIRijXXG8B37G095nuJPIvJFAYeewotW7DzpmQsyOCImgh083TgOb0BXZjB6zMFSXmJpKucsOU
fK2DmJkM2Ksky6fuX5foWUZsJoS86tSDKiI0udEUclxAxFC5PuL8sOaA6rfnATwNPi5KFivnLv1M
MN9UP40zgE84shLlXwqSbKSongC1W4ouEt3Fwao2R7B11Rrt1slW1mZnaW1QZHqDic51YSwUTUtN
ys0YhbS7lV7VWMIM+B0tuHkNqSSr5yYYzKWFYXz9NCJFnyQpVV24z1TY7MAYpqmSnKCw1q0+7sMV
1Yu/Y7d+sEjqgtYQqOW/a8UkZ76mkpBPrIas5354U7pNzru0E4H40/KlU7zzgIwZOTMzMWde0ueB
200D0LL4IvWV/I2met1Ocg4dhMIiuOCv80BzpmhZXkVvxABcEVICffwlZk9Yn6cjEHWAo17zwPPD
GKpo+Gc2gUQzej7+HXEP/ehS4IpYrre8eIUtFR9ILqSMlBYdM4CXijYEeqRs1LwLT8ofel0LBT0Q
pkaOm4l67uThWueiy02nbXr3z1oOSqstBkO5hvf14mLUsonPDFHfmmtyWaM1cJPbn6nKHfRRe6da
fULA0XUlQpqeDOkKf/tDfQdAhNv/jlRwtWZ3jY42m8XNTEx7Ax6UB/EMoDmMNqfEI36rxHck2BOo
uJCglrg/ye3hlK9vkizqB1vRO6LmXUA88udXjtpb6rCDXyu7rMAMbm8812iyzOAKvD3PA1uEramo
qzkqyT+pFyH4t/0dbkI2ET7pef95kTxy0B/sphz4mn6/RAfdW8C9coJYyOKjYQzSyqUdtfW0/HuG
cEUZlQNzLYDh+yhpk6Ntio+bomXZqu4CvoL7qcWBVPbMk9VcFW757QlBCSq+jYcOjzFDCGkWxAUE
Dj/k5KMTIcGndiJoxXiKMM8iAUx4uuyTb/RtJC0YdfVraNuVvRkZgDUGlPqVhIc5EhEQZKiG6Yl8
bPtQV7ueM3TCQuJCdKPJa+wJ+nBYSBuauvuy/6w5Y2HMwBmdQMMPv8n+vdoh1OWwlq3I+upI5/Zs
kDnG0N5MV6NssaWKrYxIwFMNXZyQyarHxM08PLsTeTFZ9vUmNS+tr8eyCLFYqn6SBy+DwXcy8ZcF
VNrOAO6wSU1b+B8tpfDMHNXbCqgTik0WqTEzZr/Avl22iLJtunQrJoDRjLGg/NTxvYh4PXlcXuQe
MF/X/sfltl7wWSSDUTBx+kX5FhYyQ67Jgy2fD4AaZdehmw7d9a3LQoxvUwTq1a4=
`pragma protect end_protected

// 
