/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2021_07", key_method = "rsa", key_block
NtAd9OZUX95s/dSCRNODTF9HgTWl+h4DTOkNb9Y3Ju8T8NsGbsgq1H0S/UY/ncbohmCQIVToM89N
haVItze+LvwnwYWnQsvE2QE3wSn2vHQBgtpF75htH3YYukKxaf+OWkteqlivrrYC67CenOg2L+F2
eDqr7yjC6pMxu4Ko0VI7zbm7JD6T/YF2iCb7EOvSaTDEVWZY68mzTG9bIUY0qZtjz6l6XTv3Quxt
aEodQdzA5VK7AI0QwWxXrcBvzCCG0Z+LBrGFhpzsF4KSwOHU+jRAu6uIF9Mtk7xllqFcpU95pCXa
f9sqX/ti/taMnyqGQUTUL6eUBij3vlT7VnLfBQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="QVR4QZEDqi0w5f9eyB33tNffNvNEl48tInsLa5sl0gI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1506848)
`pragma protect data_block
Mffvdu9pcmgNJk6bmxz8vSc1y4qDcwFKMAu2A1Tl7SURUV5S4qUXqUs9LCah99yxGlHLtVI0wBag
/C3pm5JLFDhxJ7YFA96o8Awe+Q0BEbUaPx86Zf9CIB6HcL+mqbqh3ap5lfRtqor6FIEM/UJ5gjj6
pnLeGbZTpHWz9Afv3EWeCe6OabIrAK8glf/+HICoxgDVA3wiV0/CKkLObJkcx7+4+ghskaDUCxJi
QFX7yIOXiEYgKLEHi1S+b8EGna60RCBaCtwLXvfdpCcsKAch2PEGXiL2fIDD2/VD2Tz+5vuRTowA
CByHet9QL93LbbsKlYPjYTJJiKGlCxSKdmGh1pCb23iPBaYBCIgf3+OgZeIdULHeyXvLsaH1dsUm
iAxEGOo6pQchlwCmll+RjybDLNgFFamWZBDhSsY3339AAUSCjFqDkOzatZhkq729Ty0i4vWxBykU
u3NiZS4u4UvvL5ARzZvh82BgXo0qXaVVL+ZgEF3TCueZquL/wwbg2BkmK+i603v8wtZQqovXzK5F
J5/5R5L6PsrA9Txv9JKqH/7XeQF/9umCx729i01o2WNe2ULUmHXK3pIti7miPg2FLyhOAs1Q3fiK
2G/0hWrzlTuXAHjA7Vzw5UQUULIWv+vbCpjtndG9I5PH6C+Fz4XmT66q1NF5eS6xB95lFo8pZF30
jtEh2v37y6YnZWfsCy5YnB/3CikDtLbegxEjkeK1FKZFrAaF+j9udRDAzQVmGCvp2vIbFIvxoX/T
auTPUhTljZtDtsO0OyyxsRRnQA01HxDZTug9+CTMWN79kmSaQjAkJPB1hu0bd+PplfKkqlewfioC
D7c9j3opC4G44aLTquSZfJwvXH0q836P5NMcgHHGQL1h9Ksi3MYCAXzmxja+JatVtItmbr8D1iC5
xHyCfTZeN6owwCJPwcGmGUw7UpLbrU8OftjHyzCou1ak5j9qq2Pn4MAjG7ju5QkLcvKXAXo9d2gQ
MNkzDVMNUdg45UxmPSG79LY1kRGwDNOo9pN4doKx61EVK5k8q3Deq9TA45LrWJ5Pr2lROFrQ+9Jj
rUGlKcTexJQNmyzRCG+5hUdTCWJH7aNxcn/YHeuiX4FqjXA62Xdt2t2b4iBLYppBeL972VTt6tiN
EjcydOLRNW0uEhR6WyTUeVFFw5+31YaxElf8R/F0oib48mDpj1SsrHhcLaOz0FibN1PVc6OPq4qN
PCS4EOuZWYVlXwTBWhguLQVdONyMSHmRJh6CF6tNcrHc6cxR0e4QPzNnyvb3Cm3/BYyg+OwbTTgg
5gg0odEY3MS/Txb8/2q9OAHXnNQjObuB6jPf4Dun7wegIqZ20zEGol6F3F3oTTTpMy74Pr5tIE8E
k1sI/j5gNcPIMahJ/pBV55FfAUmMywv7Eyoj1AtkcQxH6VMI45OLnG/i++ViXTTXMT5Lga7HBSVj
4gcdhJ8Nt+ofkoTV6Sqgyqwac3JV6ntCyMAw5GmMZ4W6DRRI51LEYEyGNzQ65E5ocqsjz2D/tCqn
f0Lzbv5QcTFF/6f38iqstOd60beDPcMdkO0wQgxY9jv1EGCemtwCVvLgRi2RiTUjpgiuKQ7b3q2a
qWqXlYkppRDCvDfmpdWfJ1X6QFg80OHvbTFY9u/nQQljvvCgLhWilxHhSgjeJFZS93g3e9OXPP2M
2U0j9UqpXF7B2IDvPF/uEAUzq1TruejcVzohmP6EKt+B+bYZjILfv1f6xY/ls3fs2GevodWRLBtW
jr59dG2Xj8kWWSeFhfuCYP/bQYqcQg3zAfLWKzdWHbczQDLoTvcnRGoGwTWNykymvtEgiRlVrffd
kB+7x32ICE97pCfLNNf+qbdikh9mseR3F0gZsVQb/BBKx31RXhTPGMu4yGloMUfugEQ7+qOuannh
DraQM8Atr4/qnFlixHOxnahJ1VpvfquKTHpWTRGQw+kxUOoWg0c7wL2/UOTvebnmrouA1NL6Z8Sn
pGFBDnNGcMasalVMA7UZXdImPuPc74ZdSvhQMUUoN42OF9GGGC3KJJJ1USFZUJv+IQOYUNJ6cYx4
9KdZcEVTjUU1blBEtxC3Nnj9WvwPCt7CWq2OhQ9On50MHHgfPfjaZqIhzYd0qmjgd1QSwIBAXNKH
iTlyetxT8Q9Py9qi8gDsOqLIPbaYWRPjb8bKELC2DxJJToPif0mH3xNpYVXlDOx6+127mXCS7vUl
KscjIFmod4xrx0oaiuOh4YiIyxyvTdv/VSnglTw3mg0CD6atIW7LWRDkzRVra70xFWkYPhy2pLf1
NxLSYXpx322B/er+ycz2g489YIKeQfhxnvHkfgRRbv88W46VVAHZ85p0fHElEOnJcimYMVRCEvKU
MhNhOXt6IoVGmkEOlcFXmDrgBvpKFucOHCS1Yt6Q9/iIUmPVz57SasnU/9q86IIpSvtHJ3JjmKnf
0NpEt6w6zPx2WEaGqSxuv+DvYsSRi5+HDF6HJUXR+f+CZ4Q7IpuxDa19T5r/vp0/7FM+7klxKBdf
FeYt00bI8N65XYCHvU4avziyHGSU1tzLQAczondLcJA2Izn0+P3QVLpjInuwPjeHKSvmzPmYBpmD
UXvUDT6Q2vdZw7cTE3B57tbgQJYgbuIdpVox+8BMUfFawjxb/A2EqTmeG+nCfMHeDJLDNfvG7nGb
VMNbsH76nfL8XS0FBJvgE5zCU4bV+ZWymI2GVl9S2r511zBtbr2tIDwCVHt3izR9yDAKKDJbWH/4
2AckcahidZNQKfzYkQytP0e2BeF8xGz7VGRAw+gutG65rrrYJFe/Wi/46ma2UU52CMqUG0nO+sCL
Q4Kg2S99VxyTqie3aKETJ0/QPGhvmh9mVTrUwNqPkUf9PQ9eF8iKlezBKVcYIWuQJk76ZmZvIf9w
56ez8ElKe0+Iuhkcc7xz2E/U8nimQqqggEijhG7/nKs8PwQZIye1XbmjnJGO+ajUEdo/afL4kbIE
S/e/gJYYT/nl0Vtm0WFlGvqPhtE+9oduc2NzAFDdyKsbESLl6CZuojnT8zzMm6QCNXSTPqZKoril
7kNu6BrMxvZyjdThZFWA4y5Mo2r6Uj/Ta5LeCjI95623CfHY01MpTbjzGk0BeExfN9zg0FdDlYvr
ZFQRe4nA3Gs+sMWBULsVwbSWN7DQxS2kKuFq52wTRsYHAhKgH1KfDW1aZ+twaXO/r+0M90cOk6kP
it5KSloJAo9qccLw/K7Nj3oj5O9L//MtO132n1IM45hCFfKa//E/aBXNF0ZTTtmBeECsqpbo00Xn
ae1Pkv5INfdH+lPsTzkZI5DqFnhKfMiJ3jDXBox+yKU36tnRdDmuvJxW8UoOthRGYAKCJy4Qy/cd
fuJxWdKY6JL+b0d+hKACrCp2/D+2mtTveY65D9IWVWvVJESzVkyHFbUE2/FsscwKx1ITnqhMLlao
CbjENTMLs0yfH2WgA8hj54XeGHkTcb5TE2yP/yjOjvMUNm6BtmkiGlGEHGT/UJWS5o5bK3D45lnJ
LukzhbBnIdMmRJ8edRvXd//KFzgXcQtbQGSgT3jV91BiaDDM83Ao6A3p+zB46KGv+BMb7xf/2MT9
7N6ObbMSU2LmvfVUDqzSIQtHlXiJ5zud0x6K86oG1yaCDLpAhr/hAuBWxEMAtSpgyMf42Be++JHE
UmlU8kJ4yX2lioGJcIcgapHrSQk44uYJFRsm/Hhd0DzkIX4jJ2dbGo64Fnd3viUgHqrWLh34pS7j
Z9LbJRq7EWbrn92/hIR7RotrtIZfFKKpKMTh06/BDbaS5tn+O0hne4EikS+gZbavq2JwocQC9lDS
oI7OBLfcaD2sBxaiXJjRx2MHrPv50LFrUAlg3S6lVvphLrsyLIIc1mu+FvqOoq4cyNjTzhbuHlFL
kq6SB1TNZ7zQLrQaEiWMZsKz6M4xIqUmiZtjLGLdae98rUOYLkh/5zXHsjwkjlKy5wgn0KAh5Yq4
wKEPlKtrSdkvHYQzPm1VQsyBwazn8C4iJo75sUAAap76jJQTWuUM+oDhTUTLdC8DuZADa5sjgkgV
z5DKUFMK9mzw81Q5uirDs3jwP7I78iVPi8IA61nOASFqP3ubJXaGFpbI5POLHPkPL+hqEccn572S
tOjqqJrq4BPSvL46kVgubcnR37gIqMV7etpD2/J+Li9JZrY8aE2wUpe1N5+hC2mGTNqkr9gjidxg
ENKxjLRNbslvV4wwlZ638w0u4vzU0/mdp6J6BjlRi7W2IuvgxBwuIgd+0aHJ/bmO9j/odHeK8iA3
/C4QxuIaq6BuO0KN6Nt/lGeNki5YpYmDbI6PtTTDluUIUR9GoKEnrwzlrRKdELd42MeD6DlBT4ca
zPLvIDdDo5XapoAxwde/pQQSERMBbTWsGLtBTga9jWGQOovRrvLjYuGn9PJzSWiidL5PN47cHHAA
OuznaMkcOLxjaCwzonZu/BiivWC5LMP7CahaGlYYvBhN45g7fFzaZeK9eTBI8MoIqrEwDUzLGTeF
2l5pklP9gQS/Rg+/ewc9S+7jgmfuCmyC22CPjzEutn/E145fUdc1BoJoK1H55Fd105kVqAvlZ+qR
AApIWQ5q8AZJz497bEmfextuegz1JK6dYB2/JxNNemhbM5ghSUx1/SgnwEgkHuD2Raigt6iBkyg9
+Sm97Z9jzddjgWeRHL4LgPTQEJUrWlabaCaJohLp0hblZxNei0QeVJewVw5hXdk367i7ABZkx5LP
koYb3eTaKJuYLCsxcEpr4XX/LTrHT8mjCF8tXpTfbdMXej8ckpbI84cMxFqKdaqs3g6GbGUAa4FS
Zyy1VYlUaJW7HwvCXHMJkC+5F5xDcGSPLV/+4vxeHy7Mmu+KyYPNA+b90eYRa5q/uuCxVD9S0qlk
6klcHRLZAuwMF9N/Med1SmwVPEG7A9UXWwKt6QHPU5ARRq/eVt8nnQrTxCJw/2xhGF5smGOBp9hl
mBT4/i2sguvfG4qFpzr8ABVLHBtr3rY1tu+WinRu5o32s4M6qzbyuJ8S12TgrvAsAGMF8TxLyCdg
1iNZJob8MkJGx9uZZfRg+ZyxF+HUIIz8XGPro6MMVb+ns/SgU7cfIDyY1Hygly28jzPPdJqpCgKI
vpHUNehhuQB7ibr4dXEzjISBna1ST4SXkS17s54opmFmbvZyqEwglrpCj1DXmEUzqHwxS6+E2ZoL
t+3BYZDy6cW4LeAMl+cU91YZDEXeivEKbfB+Qxwm+06JOCl0LPMcwdhgpBCH9V8paf+DAbsKReoX
4i/e5tLoVOWHO73mfQtt4GDPdVRBd0632/BfMQm4a71o1UJluApf7LnR/JqqTbQON3LMbiQ5gP1h
qyOFlCRkRnpri7oxLOXtKzJb0CSsQNV3wBnrtXW1xKNxwGjkBMDMYOPTbejXPC0IOj6IUk7/2ICg
6Pz/CymDq/ImWQekw9tyL3sh7nDrTz1sV2ic67KERV27b/QZ5ixYLSf6qwdcMcYt9VfS8+ECIUDA
gHVV/0DawAp0BHWOP9LNN58ejANt4jBl/i3lGrZySawSldzkcarJiB3UBOzMLg+qawKF1y75KfAM
YSbm70BLqSbVEFneQ8T4IlIws/6j3uUpeMzOqi0rlkwqQ7giLTBvIvLcgHjmV/AXtmcHSULFeCg2
/uAs9l+H2u7NdJuHIEzWZ+VKwqqxnkuvwB4H54T4ZRpDKDJJBU1W6IdfapDQYlAWh0b9Stf7HD2W
SE4fa36XdM9Zu4WaGoXROl2aMXgPiSNUQsesRco42ylkmr9Wms8AwwAByKQX88PoLC5tulQAUs6p
nQANkn0b4L86cVhWGFEv4algan4x/K6GtAgJV73VNlFTYk/gvxZlri2DnCt/s3YRkjEYRAEeHhxy
zw9rRLLTMoocksBo3L1QrI71bsTvjI7y/25NNK/ZVkamey0+7mj5Pw8a0GziBpbFDs779LlQ6nac
BMIG7Vv0G1MemKMBT/EM78NARtHfHDAxZisN0wyDeF9TO49V0iNOut7zi9uYLGPhJDmJv6zCbNtW
x3Y8KkANe0YsodLjgCjB6vcXGmSGdI+BwuAjw+ZBIQqCVG593p7gVii96xqhc0qJPz6ZhYArXpMc
B6uqdj5SP+jRrJN3h/eMF/KOaJc/kOi9gMkHpqptEwBWIMD/JZ5isA5y0kCRWE+bKIdl++JJRUXJ
eflBa/5NH37B0OcUv49MMNIm03FL4xK3ueli1wStMQYp1qtNz5R3xeu8hIMt082VaX6xYuq3+QMI
bPBle9rpZsDlvRs8YM70hE339UXMafacUoF0tXOwOLUNlOW901reAVOrNrHIcrCkHc1TngL0dyca
ypX0DfCGIS9JFLbXssIjAGGDmOeEcD/Am6oWn7cOVsR30gBD2a810Xt90GsHBoTSpOdxEdcFxLbh
4HwdvDQseThVHrVEO/vsfSm2sJ8AToSAGgSBBY+tWfOuxKAZzYFa8vJl0XbzaUfjABELzBxrtFA/
nfbnPXIlGWxn6GeOAOoJ9H2AlfUI1nLo6K8KKk3m7A16Ba5WB7J6OemeGz9PBkQg85NsNzWO7kM/
z2duHrA/pgdJp+AYMUNG9cET560NlJrbyKh6I3RjkvvBL6FclvAAVMmMTjSHZgmwwXIWS19P18PA
qk4XkyCWtQDG9hBH7N0tBwL62Om/27KUck4q4duVXW4eExn6PJDUJ7RWX7xM4R9dVGmoyqXZAHTa
TGS49Pk/6eUOx2xN/zam7NVxmG950udCVMvc6OhwNCUhv1HX36KTVj+mbnzBrlHMdjBJLCDVjOPj
J6sylPCg59WXxejfF0I/jCNKLW/LQxPv2tuRHgk4cbgeGJAnUsOVKBVACj1N4TfIEtw2jlCn6hBw
uztJHbc38+17ffiiJwfQaRyC1qmd1j0ZikoKYSLI5SbshM+cCALaX8EvwFZ24zlwTkIp05cdonZP
5bgU4BQt2UZNhlXqqSgIavictT1TOag96dxcAZM2E/A9zzwa5OnixAR98Za2fgo/N5WTQE3M8ocb
HFQKgJWhl8VbV7wdqRyZkgbqSRaXblgb1WyFllQ2i38Ep3y+F/ARslHVlaj0ZaYlmmAeMgCxXkKX
uUwF0McOfNqHHJyfKUapceR22I7pYpqi1/rRLVBFfGqOVICsAC4ZlDidayDZA6UGjQx+fT/cD9kE
BtuGwKMUECsimBjr1GWQQLMNbcs5OGDZOTRBaGYdLcjSW9Z00YukkjEkxRoxFJ+YOCh1KdeGuQyA
T3WijiWG04Qi1yB7mS4mgd+BNPeFE8jChyeIJ5TdMfMdM8dj9PDtI0ugE5vDIxnU8R+mGAPIDv5s
XOacHehZWJVzh3l0THTJ1VxMr1uoPIq73m+ETaAST9EuY4ASc6xBf2+pen8buDTetuURzqdmnAgv
f91n9Lx0cZ7FD2BAx7iQn5ATRACDWrKlIt65Lkq+ABpT2sBOSGxZARyIjyurYo1Zo8iqICqrF184
t0IDdJA2dGahzCrHdR/ydEEvQE/fyhbgbw15QBhviOdr+KntVnGJ4hFw4jN3rxlJ55y/raivzEdd
BUWvyFI0Bl0h0A2KK5g/qpyacjR4MbPPfcjMbvGkvbFDUAdK6JAW9yPuw0dquhRWh5htXrorDCxV
1zA22VWQbfZjFDq4gKIRzB7hX49jXOPnYvJuuvfVlo1Ysc+41jf3uwi6JRLnaE4joUK0KX/0fkit
xfcCSNg8l2QRnxU8v87IrMjTUO2ouW/Ln1/yw9YNr0+aG5iUh6ETURhXepKSZ3K4lbDJkY8b0/d7
yac1pCV2pCVsSR/ly1990idBsemiMetFoixy00Wp8DKyYRcBodfe/dc66blkXwn5h/SrvOssfP+Y
y2tWjXgFSYqNCwmnwIlv6F+eQV1wybX2HkrxlMZn5MQ1USwWGFKcwJLQ9jcX4gOnz7q+ecFTr3gM
ShRTFNznZuStOHfULM8gud1HTzjq2x/uVtk7tWSGcJcOaJcUCGE0QVgEgmHuSOK5KzmbemPDcbJB
dl5nEL5jbx3wEdwaEmDisSeqvir0dq4rpxx+cOn0cs/fk2IvgDvwlpjeYLqEGPcSx8yoKSs6yz+x
AfMl9CO+VcloORJnKd1uWBdypdKld/YT9mtO2GhHuH/Z+2alshWTqBCvf3o6/ccs7qB5cW2rvSbp
o4+vmYj8f0shKswlNx9NY+dk1B/yF41fHsed879lwMLXX9ON3DTf/JIQ7U6V3Kv58Bnsm1JUmF8u
oOprFg30tGhEbGtjogXpRf1ei+ELog2nQWNMARbbc/uTbGYPBM0G8me1tSmL5msvkwF/0AfjQTFg
PIUXS2o6dQV6Tw0pTE53L/CP3Kzt4OyK5yDXUD2aJcj3ZX4nVTqAtM4UJDxYdc3aLnXimqopm71x
IKn5caqkPpu19GcpE5xIYq9H37qPFrDypESQwI6ubnQLTbq98nwK+xTLT55JBWPEOn/8d094Kz7A
Pe3LzXUhQwazncxus/mfF70WIOVAbitFs4sfFvFRfpcnzqjFw+5frgSvBS42CpHFiJxYAA+ZL5ff
FrZfqRWwNcKIe0BsSLg9TYZ8/s69kk91UYCKnW6f5Yp7NOnxV/fdlRc1d6BrEoeie0+E80SJIVJb
mc8syNvJ+WjgGUBOLve/LyfHwGcZ5vAurmdwyFzvSVyc8tbPn6ymIqyvryytfL0OOMRPSNrMviOS
DHi1094H8lpH0tTg6mq5n/qO6Jlts3FJdCoZGhqz/A9fcnFJcNcsoCnqP8sO/3XDt4SC+YkxIRBJ
gd9Ekkn7j+AQ4IJWTufvQseJn2YGthgKaOAKXxi/NE8izhpyUeUnnDU0surq+mIfuwbX9ooGnt8g
bKj78drUULdQyze9Vf4oruLt3HhWDnOZ5qWGhPnNWA20aHVZgeALpZfTsgYQE9GNuxoL4Xu2Cgm8
3OTif1NZk2u/huDdfo4rZbjwG8fB8nPPhatBBXCjISJEGIZ9CECtq3W86vY5ciMLYgy9rHawQhQl
wTky6QFqCJB3V0HDVhl3UyZGx5cl7vWUxdODbyqYyAZKp50UizzHbaJWFs2WKKvEFUXNSUJdqYnj
JZ0LObAoicnphZxFWQ0gZdJWQaWmT5rhCret9P4eJ6kbWBDryWKgr5f6Uma3wIEVF3zNAPtd6005
ULlPXw++b4waVu1sBa/N+reseNg52L86EAEqARPIzLTcmyLZWHtR2w1J6X2Vwxeqs/HogjVP1Hxj
2anrijIdaQ4FLJPxKPkAKEFxbdexemHbnXe66Ujx5mx7rDW1A5zp1A/RWLHg5BmaAQgMm+FJnYfI
P/WEvbqe6NBkbwDtydbLKzgRpvhM68wyb+2H+iP1kF6/b7g/6McmUKaTYOzje4utg+nLPKOVVtHQ
IyX0+O4eUnRnqvjf48NPFOpUXohKagxX1Pqxva0iInG8dMh1F5+RDkz6hN7dFuIRJhGP5Mo94jp7
BBwn1VIJBzU7j2ult9MLwPGti6h3Hp4a/ez6aVvtGTDpkRSqrvCeasGPlsBBqRKFJYWE+d3br7bf
qPxAbC9Cp+FoTcvw1aAws3+zoUP9r1WGkMdnnYdP0weeS1B6YVqfKzQJHmLnBgIeKjMrHO00e6jN
7paSCnAVzdXaB/rBr7FDVKJUYTcXNsf2V5O0cVnuftBep1pF2re0qm1fqNGdHeq0wt97s3RuGBLR
Z8OigfNXAoeVEtOZ9YPfAodhdBkMV2jqqkp76vgwaL+0Jmkgq0nhtb6p9K4HTFBoU3mYuCuFADv7
SKgKBNYHf+fzbnwoynHHpKkb1cgd3WMBC1YB31ybz0qn94P94VPjmO3rVH2xnxHy+bbCBYXmzQFb
ZTshwxnRZnjXkIXRPut38QQZ4RnYbDDJyWRzk0qQo6r8fK9NV4IQKvP1B2VVU5dG2zg84zUHhV75
jKPYIufO1MSYApthXm4Po68VhkJotzqJWzdvz/Jik+w/vEFbAgjNaH/t6AkH2Xt6jRJQq8cR0Emb
cgFJjfI4yNJ09ys/HoihKv+pkNvx7ekvJCRH5kH1Qx61tFIyzCj482mtvSWD5yMckmQ2alQN+Khu
YUmeswBWnuMGujkaD2jhLsEcP8zYTCXLghYlEBczOlVHWfbHgjRAwmEkUQOP+yvb/izoEiwiMpiL
DcANuWzq3FIl9S58FzUQfaL4iJybrlbpk+ohSZNyo0s1z9tWcOE3i2i3ocFI/l6JpTOkfFVrr/Os
kIaIWexV0hJSA4z0Aon3mygobW9DynU5f5oAcDYFiRhwOEngNqMPYvghDBENoLfxKYiH2Mvhn1jL
gmQapOuMp4xxuJzW1uKgAJ4q9dGamXIisGSkamdsY4DRZiHWmgsgXUbh9I4W0IAeqWHLhrrvIPpW
RwMB18BRVG/SLXlg8xPwaoSL8XE/DGwTje0USVILNfBoTJ3r2c26ANcimeeCqNMOTYH6K4y2Az6q
M7smurYjXCGYi3rJvbZjudwYHEJSlCGvcfw+A9NeLkshDGd2SjACxPllQEFmJivex37CcqnqSdHz
CksY4J5CMIhkbAbCATXAJe2HFIaUUW/8EHtxaCMBwfXYk0/7C/aDJ9Im/CCaz8L1KupVturfXrkR
q2zwCJkPAa1CemiYi9KbV/0efyBzDegzYRfO6O/0HfUmiimoJR76TDLsj90blyMSSABdRvsFUv7B
+jmu1pPtzjMfSGnm7WeJm9SU4J/S/QVtnsy+TznTQ8b0Uvyv8lI0tmCj//GyQlIHL8ycPY+0sQqR
pI1tjzRm0Vj4Fk+j4Lw0mQYrikEfVluQXXiaSzlafLUgJXlYk0Uvutv4aMmvp8w8ozYjk96e15wa
MqRlFaPCioBVzY7b9IBb6I4/GCGbrOFNniOxN5DOeHuP8PIu7E9OF8RQl4xVsix6WeCoO+nIcYMY
7rDJrgh9nS+wosbPWNuRH3XzG3SWq7Fgb+FINwX1ygPJfgZBqGyDR5lDIeE0sNKow4/3CsjsBZTZ
STpgHzmzu8n+jKrjvK4f09U5AoCZ8TIXiLiU49/hRjWKqLGJQ3wqUSsoMQK5ZeeGhhpgRLXRDcat
IjQoY/61Ph/PRaeuUSxGAfZeY6ysRTzOGwO2JH4DPiSHXpfPlCaXUwiraWBfRf5kuII7f1h4atQM
4jesJc1p4L/LBrKTFKRmwBVhijssLBJBprCpFvVsBckzfGyt4iGGy4D4qr0IcNx1Z9BzuQFJNNgC
4E/MGbd5kIuvZpGGGPgAwQtuHSQLvQkdujdg/N6U48OkVMpIJWxaAowQJ+eX2PP4mvK3YS+DL38e
ldchl9A0Dd82ZPY+FXmt1pu148ZLQrUmt4Zjdofi+hdyrbvrzmVJhYAG5nu+RmSU+nHBhmYuXoeI
wVjzMyIBOdEZGI5KTinE7G8bxxRHyTADSbmi/ZhI/g+hXVBa7m93Fzt8U9mzeULGHNYD++G56KKp
3bdaAf12C6H1xVPH0AAf+kwubbKe7AWkkgSbpeRFbfDnP3k8t/NyyyExUdSRkgPaoD0EyMwgUxuA
riM37qz7Ht/m+9he7Lb4JRQcj1Gzcn9Pnz+3BaMbCpU5TIki3ScH7OWrCOhMFbe88sPPNpZeAipF
M7D4aCIY0KPOIvkg7lJRTTJfDe2zW3U45v6pTz/VElXu5Xhvc/WCOOrqZrYYPMqzxcDYyxQYWPAO
Qc0SpDYYweCQtLK9PFqm3YoN49nfUmZF6TpD/tsboOBVo7GowF9q+83P0cix77VVq6DxvSJjIqnE
AVLlAZ0UFJDbQ4HCwckD5cqeq/ETnW7Pj3o7W+KQ/ZwzDLmSuQejbVwSUSqpGaTAbIjK856ZHv00
+81LJqaidGf3EV0XV/KFqeDtRjpJqSer2vjoaen5t2LjFiD2kSwlRp2k4qD44+wmIA96BPeeYKV7
p9S/VvSkc3kQcIV4hygPpHLoLr/DBUZorLsShEg41YSKok2PuuAtabk8G7fp+tjTmMSG9/oCuPqu
Znb7Y1yAc6AYlPuVDwt2DWEgbwiCLh+Br9vnVRzx7xwuG1KqGhk2fmvKPdgr8YSJiaAWriiJsrw4
yhurzbMZ9jJz6Swvk/NA6nGBycGQFqAHF9Ct6SJfgCFFUQtOMuW7aNgOtszW2zL6YTVm73IxvZ2M
pSeGtXm9I69InTkrJnummJ8uYb9Wfx5M9T3n5Xbd+/uUL8NRB3+4ioegVQoD15H7JM3EpT6Qxou6
w65BMACu4TrSVLe3WDkKg1xP8hzLd9MRiR/UFuk3MNVH+NpXiUQ1bmpRnwhviE/4CHTQ2SXlrwNa
X8Lz0ZggmCZSEGne5PIYLuKPrHHzT5mmzsaYNkbA5zmd7Klv12Tv5JmvoMCmOsB+4ebaEpJk+J1w
sjgeqGNpNpIqJALlEJh+bC4b0nhFiWtuljCEgAcB/b39DwCJFvB5CyCjVLKsxsPh4k/6LWR7JDiD
v5S0cJfxhDrpse0WBOZLg9xJKhk07PzvE5zsagmY/GnWXX8jI/s2gtXT+aMpT1mL7Y7379QIuK3H
JrUEt+qACnLGg+/r/7UophTXkTlH8Tp7BfWtyY7zBbpoKStknRyxy0IKtdsgiff8/WEHfuTbO9es
Qe6fKd+0I+0eGjxeGN7Z8ruO7RMfjbDWjHrRZnbCQj6SjqW081BWyIobnFkPDmPmq3m8kLa4ENMd
8lwLgE1gUh9Cq4G/rXMrAYy64VTwp8eeWhVC4MUZ4KL5q/UgUl2Wu56UKU33OFbBg1lNv8KDoGaO
dAEaLRDkVv7qwxInzVDw/I9BheML4L+IvAfQcvwOEJfEogQ8g/rwd4k9qa8PC+4e4xwARIpYTfoE
BkrFE55TTyfa4BkkWn5AtTOwNocbaKRrD2t6zfJGqoWX/ahYmQn8VW6hsJAzTyrsyTaoJV1Qc9yy
S54Gpp16NsHrz5DTFRIoAfhiOoe9pGfrazCgBe/5Nap2nGAuK4SdxrIxEmiJUoYniQeBwgOqqhcn
llOcNynPQeYY3b8q4ZE25amH1GUom2ot2d6sCowf3m4hE8dbkKKz9V+AlB4SPRMaAuRPxlQ7lOrX
OTI97c+vLj98XnGH9Vam3JpVhzFPWbdJKqqO8TiYZ0z+q/2Ruv2hnpWRXEBxDJ62KfkKGQtt0GrO
CJ1BgvNorIkTOWBHgfRToc6aqIJp2NllWiSwF9hdhQ9hL3w844VSKAqtc4/qcO3BwUwmCOG4v7zq
p4A/6GL1CuN5MFwLtyAiUtiGB8UN5gFyq9MJ1moi2G4mJg4m/bSgPoAmJ0BsJQlM9eA1xsVxNsRa
AG+0En6iIn9s3wrRXPZZ2Xn1fpyXkkvobb4vgMX16H58tzUdOI24COQcgIfUCn6ttWNSoQ+Ga+cv
8k6Dzvcc8iKumplyJLz7E2jNAvNVd/9BifYkLjjaDlJRI54UaTmtJ+jtLm2xxrmG2incekRzxdjQ
ABliRQoUPxhg84usyHNgw5i5bdkwMbSBdokJ6P1ZfXSmGdBfkvGrUsRsSGRSlyihn1pPl2H7BLdG
VODgiWv8T5nUs2EEpxlyJOdgc7Vl/t6vFgn9CP/7ix56G4Cnx53NB3mDE8QSrzWKlMCOpC6UJDjd
ItfOtVgY7wUZ7TyDxQWJ/X89W9hkcIgo7uQdZ2aQu38bdoTlthW0GIaTLfqw7TANQCiY4QcOIj0b
8akFEVKn/YBwuuHvrgvXM1SL33ERcirSXiSZaZPsbMORIzcdOShmhR/8i7dL8kWojCYpF29MSuGT
NKaWltIfnW5rxhWSntQSHQR/H0Be0k9E4ODH0RySQ/0s7uBIPGcjYKD/TtFM8SWbsd/kWENPOgjn
RXf3YNn+jx5rsW0uL8BLb0oSN+keN6dy/2KA5nS/FLSP9CSIYmWeK2wpmHkN/nqmHVQWaFQmY0/t
BwJUCirtICk/+dyjs2v1nwUCjK07RpCnblgCsyXGwXH1/PHP8l1uXxwdt0V56zYp0E1aM4D0mSRK
rgrkogwMxS62eMw9xWAQVlC96nbi63ujqBYkdUTTFXigxWgWW04V+mlAdpjRUk7PiOASPkSUartE
s9MxOm2/z5TEpWIllnN/cmAryXT3pGhhfPtIPh+Ut5kPPVigU+Gl2+7KsXjEAvVSwhJl6/pN4do5
xN4vY4qHjT+dJXoLl64w4qJOaHiFfvCEDOPShxNdpPkmmHFlPruPSaLZcGugr89Qqx8lA3ZF7S0q
B9FElDm2T3zeFoJLSTHbJG/5k8uThBFxbT482nirVd9wI0MUvidzAR1lVNwjtEmMf5xq8ht7fLse
ZrssdMXWVeJvQUUuUkaspHCWZmT1mrTR/p6VJrs8cmw7MGV4fBIgMsjj6gLtGRPNPk82ilNsfCRH
iFhfrmeSQJx8wTd7wBouDxVi8MVT1NJSeb8o1+SlVrZmCYEumSe7L+BK+jd6geJOmg8FL5liw7iB
+yo0gbkvUA+NApBQ62FJxMpo+yUFZvYQ/sIbcGezcH09tkzIgFhBIxdrnpN2CpFvC3fRZ0uizowM
0sLPAP12qhq9+rfU/dT+YbEvVbWwKk3DEOW3RwQ4TpATOHMv1zLsKPmBld1KByzZ7iqziqhnG4Hm
Czj7mD9hwkRrzAMnCGllWeuZajZH/bKVR5hNnmmnlm6J9VgfCoI6Gw/l7qzT++QOZLf5LpCK/hfu
vK7g9KNd0AKLoTo6vGTmz8SJ+eW/B8+rpZ//uZinF0FbggHjI6LVON+9PK6oxes1R2Uv8JYWlTL0
eN4b6+E9T7TPFbyGMmFj1CsMInVXb1DZSq/607gftrHtJ2txPILq9wSpyfjz4L+xqDQsTvtRoWLk
92C+4vjFXw7ajFwut85wCkFt9QE0JViY75epl3qsvGaanfih3btBJAdV9aDzrC+nr+ii9amKnVAy
D9PESNtIcPdVXqGPDHZhXmZQnVMPa+zIr5HWL+HhaUPdmhvhtdwd2wD4+cnZrXX6xb7dOXeGeHVU
9tcZvjTw87ZMEKytbeX2ht0KwjjoiHbjU54pyYNiGUQbWjpwiAo/bCmtr5iMatcd7N9cwx1c/B6c
Z9KntS/RUPkSgCppsNIQjr4GVCz+31ffZKDvIrOnhoWJrYcEloGVUsCgU5oaiLKnTwcYIpyyh8so
8jUlxOLoTRpw0zVqdcuEaciedxBpbX//tK3eVgDLVs4NkLOICb9Ch54vzdie6X6mAZ1cXXcFAzB3
So6ffUFs4vhWzdzBVC7jYxHhk+Ld5wIwODmRSVFGPVAKIyvO9KVWg6cELDpd+8CA/6dpWArkuvHY
L4WDBKIp0xwWYphCctFs2ZqT8G+20F0r1kuZ2dYsc9wahnXa1GzPP1S1/DKQ9X7DZQkWt6KqL9zl
d60MneDUaKBB7T06BnTx5Opzxn9GkOSAvdcnA80EdSYqhsFnkYQIboA+IVyHvvpolF7MbRnUI0S+
VrE7C4rPnbuEVF0pqmlIcig9DcBS3SqXVLMKNGx3oNE3tTyzFAmol0RBZMTOFse/VmRnRLH5+Crg
8wlC7Jsgaitw+Xr0qjGN8HBtQZIcs+rptkYhLhVmBcOmngUmMZ8iH7sGhwW04c1XuiNB8n/w28aF
fwe7NvTCZwbzVMV2l7JVPsPeZ+ufmfDhladfYztVFuhSeaK1PteReZyTqD7YNYkPGCWb8Vg76dZ+
asJpl/rHpPeN0dso1tHDwm3QNeX6zoqJEmBwTxFVaPBaek7lWeT3/3oytDvriE37gjiuwWNFmdT/
2gWAgcSLIILxRKYe9XPoSAMLlSsWTRhmWVBqNTs7YNQFLQ5CDDSoI9/VimF1gePJazwLuCn0NeeZ
eWasyMt1rw4i/IzIndBThzbHXA52jiCjpNJqGuizbt3wO5UW/O+QmVBBBcN+hAuqFAzs3UGRue88
7b7pBhD9x1Xkk5LRtvIG+/Gpbild1fhQP5cp2xxTXmbslem+VFcE5pDvexoHlvcbTkDuKNoIUBMa
3SsV/cYheAqVfno3vn2rn32tGsfMmXKW/Zn+Ci9xy7Lf3vqL+MxkXPm4w3FRjY9gKwUWjnp60fyz
FcPbf1G4aULb5XmMZleKINMQSoSusOEIrlXGVI9ytyl3ROAib6cXcFXSRRbH/KxYBqYCiDArcr1J
9Wo2HcgaWVFulon/jjLBNyOCzqpYETS7MehU67NOfNQviO+ve82242ADHEwjXhJDAXmMzG40j1ai
vO/fj/EEZD6LSpkATrfn9sariw+NEnIVKuRL3crhKIgbAl6o2jxJpl8oAi1U5j9DhiaQJPZuQesD
jJPAt2luLVfsZirAfTuFuty7ecWViN1EDLmFsYRG296n3fJUayxYmWksDDKIP5gm6pFxyguQStAQ
89HGAJrKwNEv2c1KqDKtForwdQ+AhWE4WbwRJ7UwFkyhMwpMQu962qi5Y+mdNHC49k4DFCEOCPt5
uKt4C6f/rh4Djif7ucnxAdI3IRFtPQGPYC1QKLb9KFMSYcv2bpg0ikmQBYB7EcAxU/PVxs06pget
hiixP2coIu/wlIlJecFw0+FVGOYRDiIUecQM4sDI2J/eh/wzFXrkQZNpSE4h7dfMFL3/CskwL11v
Xy3VxDKun5miGeH97AY4JuUdtg4SB9I76pX+taXmF4A8gfi0tLdalwVm9q3RXRF8TvUD1BMvZRSi
6o3mbldrHTFpmIffXMvIRA6zk+RET2uuY6VVXSu2TOnEWO24grhTjHtUtNBplB1vpCbzP3Hg/mXv
LCsUlCpWzVGEiDslcO8mCR9yZiUb6I/uVSy/uvcUs0XlRKs5zLAqEBfBBsGyEX5sJabCvgqf4f6m
trl+uxlnPr1rn2IDvYt6QA4nNTeOeAt+TjwcZMmOK41zoFz0+F/zxgJJCkiWWU/2doEPZloUgisv
kTTG66EnhYZ2cnPTiEfxjgt69vMbcrWefDpM0RxZSABVXi4sJsFLGoAcGD0kFu41nBFQgug0yG6u
5dTAbCiCdHe5asqQ1KsbrEVRwAFl0mx+ZoP12ZkZmuSzWCjdGRg48SQU4AfTm8yOtEG+zT/bXuRE
qGI8tS5MwABWEgMex1U9Qv1AcfqcBTMK8Ro1eyQoj/vm28A9GfE7FVnihvVoakvSJ/llzm9ZyPUj
/ucvoV5TRN1PrPudNKjlxoXU58iNSRKilMKRpaSEi5fYxR1JFvjYDlgS2uftILBMNobCt2HZuMy2
R/+pFvcduQmZh9vh+jVUu6U8HjUmmnLSaTsNgq8NksnDRyRjVAlcbARfoWJ3J+8e8nbqbIETvzUP
gtq+2H202EwZ/Rukd+37kfrXfEWlLynWDEaoJY6TpXJOeGMUnJu8vsKzm/CNh8RvGbl/UAi6FDjP
CcYy3TtHpKf90Gvz4yYuSIaDNQDCIR2vKc9l/rgK8pTr6Mqaazj+KliC+w7aWJl7DrQEFvj5aoBd
urLk15XV/Li+7zelU4V23AyB8SljWcW33QrJCwAYoe2BjFG6iU7NY2wxi5g+vZJ0aYsuiF/aCfIx
Y4FTRcN4OQJoXCUeb62NVyftBpz5dFvsK/Dc9VZYeBACOVz5yemaroucie07+NRlTGwRTm1OY/SX
Sm7qHFKQIUGy6GKUfRkwn6w6iWOvDD36I8wV7AT+Wb+DiJwk/jg6srPSjTZz/pQT+RhqUf2RvPEu
SvJApW02yq4+TSehLISwypQ53PUII0/xVJkEysGUV1h3hkn6JytWv5yZoAMOrBoxSfER61Y8jci9
1wFn1ebUp6oqL83yMpvKajpMt/x6QEaU+HdSHCai0m1xoNS1xqj3X8R7pRBCsoM5G5B0EgzmQlE0
Wn2/CxpF1Pe4pvc5Zfu0Qwvy4vz21LO2okVE4mKxJYd4cVBegrvwjVpdxXDFC1qzyB64cwg+woAd
eiof8NpZRNBpkpDbLE6rSJqdqaoPsi2eq4dN2MXrTV0EJh4X5oinETaoGzLbdmNCvHp8x7rUUJR9
YIjFgE8tni+gTpweTyOMdPj8bgQ+f/uVzANj6M3KHNKL94uxZ2pQjgVS81m72QoSL34XvENDkBBD
swAJCAaSC16jFPflcn4f+EmBoJiW4y+/dtftK4Ol4rXW7m+kc8/qspeV9kzg/r0CYGE78kAEON/S
VdyiBQHgDpmTRKXkHHxoMGYGSUi24/CrP+MH4ZTttv8RtL9E1YHzktHag86NnmKid9D7iBg1GPmU
xXG1NySujHv2qlZWj02daxIu2G0M9QF5CGIy42SaJlk5y79idqh/jWoBlbojiT/n+d1347AP/NaU
GmvIJ7/5w061yAqG1b8GrekYsY4VTlRF7iPieWTYl+fcmAYsng+baBaLMgp30zvy7GP6eobjZlGO
ysYsFNoktEf/rD+cydBx7Xa8aAUdolbZDRuc1N0/xrILSSFv+VznxFcLhFEE30iOo/T20YnH62B9
Ha26SxiaSEzgAMNstrL4D5c75CPhd88QQVtcQxKdY/lsMKxbD1HMZzuqn3aodpPvLoUziHKg7TZ/
gqASSLzV6j35I1gfmM9QoCc65szyAbgAxiVz2fA1b0q/yfYl3U/l4a5Mr9OfXfFcIJuueIv6NIxJ
6VzuJtKh6vo1BqJUxk3nzkhTh6cgwdRyLJGeXL1oZLMpL5XBVYr3bHCadH5UABniwPHR5GFHxJjw
3wqXaCY44ulv91sa1IJTw4WlgC1qRWxrO9E1iT7RDPL/erVaw65+ZxYaQy4ZDAgqECOntcTwsb4G
BUUQw59X/+0sAYFdUs4OE6CDrZuugSYxRmjKsWuaxmHZjyvlFD37Y9ltwblV7HQ7aJSbXepZWSQa
CyF5AwQxpMk9qLbnnxtBhI4nnEt4/Td9TAXGCNezpv46Xa5xnup0j8xPLBCaCiaDypt2O34siNKc
KiPzlEdPS6l8m1DzoXOZfhoRsZmLpNjdV0WZDoZC4Rmz2to8WV13YrsSAq47SX4L8e1KEJg355oU
ygRzS0AbQMcJ1CeepWDx2mzVG7BFcvmgrGA+719D8ix9UonKgP6237Ayto3PgomiCOQenzoC1Bry
sxnQE+mxU2RDXeXGzoJuX02BOXUx2+7aF0CuEWWOMT+Y6r92jRsQqfPLsKRr7IHld31gPkpNPYem
p9BtoxfcaItL79ygHBFUfcTlXxLjXOM6EnWJoxQLXMKFLcITbLw9IUJR29BliqVbXY2KzfcqVg+m
Yha3JzjYzGopnJXQIC/ubRCp2BGgZLx4RNrVLtQU67CEevi4SZn2hKWOhblIFoiCF/3BCkRBqq+I
KR/VZbt0xW3vMiSvKtv2O1ZTMMjmz8WLbsnor7U69+sE4SmGzJZ1BjXqfNdUtUZI1/qg2f/3YQeR
TeP0iakTVpsbeXpXS3g3/NybivAbJ5qo9piE2XN8vyTSkpKDyLm/tbIGRvaxWkT54RWukl6Uc/Z4
sL1ZrS6AtinIWJneddeIkzJ0lzFnFRGtNrp5HBCHLuivLc9T77LS2VE7Kl2sAzaC8C10KS1d3PV6
FHt1IrgMzEVXqIO1UX/8XMUp4wEMDJNDg01BwFEBMHZBrR3OmIoqA/w/JCFKUSJMFJYbtbCq/IOW
hRV1frQuf54VT7C/Yl3H3LaNKo4za47kW8IBWbC2W4Ckki6/3TjqO7UNa+tiYfvTNCpTU/Qn25wq
g1x3PUmgSUTy60hQckt5AencURhlR/pVEXPfJu0dp2UzWt/F3tZS7IaEfjVOjRW5M3leEt/qIqoa
n6tNNLVRK4CTx9/v3hUwQPB3LRJ08uLDPo38u9iiKHBVBkCvmsHKOBIPBNwPFC5zY1HEt+bnKEND
hoffBtaqVlAQ5ngAEyTsIEJARBgxO197WrKRKlPiW/axbUxYJQHlvZjpyCiIwBc3ULZrCc4gYmcJ
lxOeUw3AkG250IM4DMsy9HFgjThiWQCpOcPGd8yrX14V5mrmvPzNdhL4pzXCbFh/k0OnbvzAx2e6
24eAah6STQ0e9TjKxFqbBhfucUzxLVFsY51aM8+LfWI9dNrEkwMioWOZNW+eZ6MysXLmrK8+HGg0
zP+/YMJtOdEwv2wOlHrDcrU/H9eZzOj4WDsDbRj/cqDF+QtGT+BNsshi+OGBtGlMElSRFb0fV2lt
KLz5dYizcKn2a3PnQaP986V1SZmAbauZJlzGqzORs8vxWudeItkhq1zQ1F7dwuHJ/RoZ1S6t7htv
5vq01UQtYsSgx1HT3zJn0sAC1A58edCn4Od3GZ1GRAaN3O6TRzWIZJyN5bQYIzJf5XaZ9k+ukZt6
csyGOxLRWDK9019KwaEruZBY9aoIxOJm2zeF7GQHLIPNlAvJzwA/Ixj0tyTR+RvzOmXJrpTzJvFd
YnqdX3h/Nvj4DqNUHLuDXydfXdmWOxswtN7ZPoDliLdQSQIr2J+CP913dbTrmEGmSoj67cC58/20
Xph0HyQfC/7zRSiZRTXqoyoMLdMD+vVEfo9SNrhlxEEFZ9QVX/IPpKo8A0ZnH4zSxM5zT01s95Dj
gdy5sgfjXWx97Kvc9PfVz/UAd1N0+KvAMskOxM2mwHl+ra9g5HVE5Fa+vHP39GrcSWFWnztipzp5
f/NAWs3TnPVPQsBXOmaNanBGRr8Rl4lT2pD/NUe8tOpYvDGF03/9Vive7kS+4CEIsxOgxXlt79Qz
Ogq9CwbkCuXwNipJ25SwISJm+0AEMQ1AuK4J+MtPL0P1uwGqHdMTWzEP8wYRbUwLiOcyneD560WN
RJGXWO+6A3iPZFrNddQGlg089Xer447uvEAsB54mbYkEfH8kuzW3BtXsQwyzVB5t4MVlLVhAInNh
1Nab+b1JlR7Gq/RB/s0y5ltWMtmzyd+UoWjbXvw6u4PY/yxHBXluHxv3zoThWAkw0q9Ro4TcrSqR
Ef3pWE7Oyv/2DsI9KSBUoi48xB6/BVTicWppzF4oshoOZsubz2xjqmE8h0XEXlD4umWX3ru+2IIH
h7nEbcHL4QxrcHR10gpR+i/1CLd1nRGtR5VA7nkp5meYpkSBMBfSgyEkTcn3+uBP7x2kcWUazFq4
COIKM/5Pq3PDY/jCq83M0t2gKjPX61Fz0D6cR0LVfqufMomRNBJnXl4wi/vUsz0TTOHb7nN/SLE/
VxkzIB1StFNxGZxngZvX4d+wciezKMyKXheLmrp3fhdqnp77CL02tGOGNh939ooLINSSM10/tImN
SYTSNW+vyV75aidXlypNNIM/px462BvUBJWDw0lFtiy8TC3f1ijg5lCZQ6qCm1tf7kbwTd9ryfw1
6H2iAnEct5zDfmemV9gMZW9HK/bFDsOQ2gDSiNXnximEKmwCI2bQz4pD6R/X1ZRjOZ7IIteJGM7M
IvYUP/KareHTEd5ScCnzTuG2gUZSjHiGl16aO7o1V1Xaz+j04xuhr6Hk+qRH5UTpr9E2nE/cko8P
gCs7U3rGkf13YypLu+2o5KCh+pjz2dPFeAVPUTqo/dTXKY09+qe+NGmr/B5opFxxkuJQNefQ7hMW
fj6vKcVk/sFs6Mwet9DvjSISeRpkMQEev1EiJdgcWW9Cnl3+K+NnQq/eVx+Yq/eM99kQcoTA7b9Q
+7tJr10rY8y+7OingpgXru99Pufk9u2xKr3elqJXdpOpRxTttbbZGgPCdiSJ/+onxjjtGPW28lnW
68Dekzt7pBZG+EZJcaV5AFjg+myBytYlXavcMHO0Ij0/ACAZEXnJW8w6UIPtxZciWwYR8CtGPNYG
/XZC8oObosbdyRSCn2RF2RMkXVvkkllSJnWWW9Gm5KQ4aFeyxdtG6J1mzo2wqjKrORQ/dTrknBW5
x2QFPhIT0oDUxWsVDYu/8sK4p8sP1DS9b86AH3Jjq0d/3UXdUZfrF9HHfSQtXjn3ooasV1qQeg08
EeD3lGPZLgLQ5h4BQ97c8wJ6IKhj0NUtAmaIBdveDu2q6dtvYNaXDP8tK2UjoLjf8gfKBvwcYwNs
RZOy/8UnxwCtA7tDUCyy8nNav8X6jVuBnHK3v48AdN30av+7SifbHlKeSrkkR4KQQQiWEvxasuTq
dFV0xGoQfsNAWeVic49XnFgDPTUSFixvPhwV6QmFXOjvCRYous7dCMZEtWFA+Po4uQE+LgBCoc0A
9LEtXY/KwAO83JgN7MNEQGZhTqBiK5AS0xjya2jCKwoki31d6BI/Szl0nivE9l+5KuS0WmUZwYMW
x/W7BbcEmuhEWB+XuZpLv53vWIwy9DDs/YPhdMKknoFPUiACYt3Qk8PQuCvBecVXKwV8P0r5PvPT
55VAfMtjPqdsjGrPMjYEZyZjJS3VLEoPlWN4+ysqe9xgxZNzmAry6HSeaYbTzAvsv8XRr5PlGeW8
cumlyYOf47ERolKYlzTWmhSWYQkRrGBCDIksFTd+HFE3HtNiVCKBlGa9d4qOANmgdCathq+fJv7o
r09lEalVx8DYghmolQOO4AEn2YJnB+2s2i3mmCRmitHlPGb7V22cKfjXrzutpfP/HdRA6FMm8HaT
BXezZFaEwzUXCNFjg6xpBDCqp+RAYHrVlKOBVJDIRi15KT2JbhvLOj3kC/PzVssgSgMLJgXkZrfz
xQUEAskLFm6G04UNPlBoI+yH9mkXjfMi7oButJBbQhDI937yalJxVwgZ45YmB0RieSdqrJOYG5Gk
v+sfk5GHA7MWOuRMg62M4bTci6Yd2DO+dPJjm6ZEDThEbAJF+nC0yM3IeXKWESjuKzsyzF8bVq7P
Kv/+kaj4yii07g5eIVRdUVXWOgwFXm30p/2m+DguZbQIlM7kdmtj+0/GJ9OKovsS4+Lks1/cEbbl
OcYweyeq9ppdZMPFWPCuS538+/80UWHt3uhxc2PzgEaqkpIDBgrtQwPUFPG4g263f4y+sjidUbpm
HkvSzsMXsAaLYtDUtL4FdoT7Sj/ZZYtPK5etP9hlDg8qs5CzUSo3mPepqUzO9e1kUOrLt04KKKd0
3HBbiBikF1c9qW6w2xdTyYo51sl85H2Z5yy4/izggBVFFaDOI6Oyh5hjt7CT4ZpbfH2ulBFSIEvI
1vk56N8I6Ie7qvkfwnddVL3ZpL5Cfybagz/0JGNqT5hWmPa7zGCql56NvzH6D6kLFEombt3UhDzz
oGdoB6L3zkNtqk0qVNt75DY30EbZnjqqDNdbkUgbG/NmlDzpKZWawzCSsa3ujN4BJXRqzZBlaLRp
tcT4AwaORk5l8a7zBQLeDRzO0C0vpuBKnNWN+3X9nwxtfW+j+RmPqDH4dqfRFMbTqsKbqkfPocVv
7YDOuTFGBKzfIQag4URpxu3yN8X+CtjCXLKKCT14d0Kj42uThIuryOY+7lWdpc1RonDjcBleWUE1
mjgCmPtL5sUy76SnS1f+ds/S6Z96PejoszEhUZv6ujAu4YQ7dlW1d+BXpV86uTGJbMSCQzYxkMkh
DSN6C11iqfK80RrMMS3vRyCxwXl+rhpeyiAXWFiG/uv1y0a/rpiSqNYwimhKdmwlsOI74h8kwgPq
VJWj3xC/Y3tybNx/r1r85mcAH0vFdYidLRfTwI4FK4fvHRE3Y6wI+EsXmt3xSUvP0RVBaFAHgfSF
los+G/voekR63APXLBni5Cj/S/6QzwKLJrT3FHN2PfEyvzLIw/leImKpsUU/418EMOKp+YAXlTnc
4UuUDBKRBNfBdgzPBh8+hibTqW1wUPEehuYsl7YtwQwCUPvNK09KKhK2u+rL+hxwM0qhh6C46CzR
BV3BA5OG/2ToHQSG+nmycLBFrVr9WNTcDHpfhp3wIUN/VyZNIG15MsiXMR7f/ONlBRXbXimaOrNJ
ZIXotOdm02Dp40xZUqRTJu3Pg8BkZIJnqAA4C3jEeb1Ue7HAC4Dq6vpyPFBbV5ZlVbJSJBWom1tl
je/hEO0F3Wo8fPKGiFG22y86V8gcdlCmv4kgpC+9vp2PI3aT4NkBROMIR0L8cd9YCmqQLfR6jOpv
rLD1jqPrq3tgNSuS3esR5PeNKgjTP6cUF+AUR9+Z2zHR9V0OZk89TQrYwqfjI7BvXAykooHuCTlu
UXqWSf9H4hWW/KPkU7Dr1mPVgeNTy0h1YS23wsfsUmzgQtPy2ZxcC0TjJXUUkuuxmRW2ERGf0sWr
h8Qc5ey7eV6ib0B0C9OxsUqY3KO50b5LkvoHNhzm4DDj/SsBh3krDPlzSxeYs9M5qo1tatvKH4mD
UV4IaxjRKtYr/2FbZN48s4LU2OSBMqzQJPr9LwKX43Ug5L8J2Afm2ZMtzqKz/IKoI4OZ17U8uJdy
8yFeXjoFy7AQun1NC4zQdMx0whYA80o7k1ZnIEdeNr38MEbnK8KRGyY5IQMGC8q8Gisy16K8TPOx
MhRK2YCZC7sXzBOlJciXopVaA3vHBBlrdD+bVF3K7luuUEFYHlY1Y9crr7C3hePMPsRRGQ10xyNz
TyB1oHgD8ZeyIphwfr8WyjjeVgqKnN674uShI9eIlR8/0UltXzicf+a4v+J2NTA/u7GsI/u4VGMn
3rAXc0uUhVDCtMOe126VElK8vRUO2pSa4hKP7EFkkm92oOS8wjmsoa5/46+iV3b6VnhqOvIUPI3d
eYvB2ts4ylqHkAtUBQ1cUUSuFIdCAI2T48M+9ZaP02bl4MWZKA1VQWGrjyQ+b8cX+0syeC/yX3oa
XcM6+X1SjZ3tv0z19H51yc32sWdycq2qPFwsuHqgqYfA3ubd8iDSKpKEd6vWgXLmpcQKFrLPk+xF
yzFmgZIE37udYiVuaFLw9MOo6inT8rE8wfSPRWWq0CVCDWPsJJeVWUFb+ikzOIVYkFQ/tvvPckua
kHYJL++2cBrWBgbpXM6x+lMOrjlM11SIZ1D3NSCeF+Y90LF4keMOor77iRfO1vnpncuok2DqIL3d
L/jcjYvKfnGbnQwlCChHx1FEeCgTmiZUKiAdr1QpBiKwaGEMbzwirFlumVaay1HYttqpUsfWBRli
zFpyw8KxWBl4FFtq0qkIBnENYTRYuQCoH/Kl6sukOOCKHLs/lNj+/rGyTYapkLXeRPxQJdb+yy1y
Cax4hqXi8JpCZsjrFaLNYtEupLO6iBZsouwxRl4umk3T+7M3qtI0KXE4xyvVze90OI5sF6BKWb/k
9cjkR5CmY5Qnrau1cJnOHqfO7iBDik0qxFuQb+UbM4fjbOZBwJWTOUlMIioCEehToLrqJnKFa9M2
hIzoSyZSrC62op2Dz3a5er9QKBqv7jHlfB1WsKgFOIjON/ufkUB0vrqN/UOaboqxBZiYj0lx0zGY
CO4pOIy2pL2BMjEAy7tvACo0bCQDr1fcBkInFbqggbsahbe3rfhMd4YIAmjkep54Ots9OHHbxqH0
LPD5ZBNy+Ky4kUdztLJOPhnY45+1zdMdLSbjCAbfkADwQn6eiFSMvFRtPmLLerPMIB6e+mkO4u7f
ys0Ncy2u8zIdQEHFxBT6RnUfLZ9uxpgmm3Cl+Ue8Ywq5HZIZFrCAM97a84RIPMYrMA+1dlQZkOJI
j78r1OYCX7fV3r1sDTLaMuSH7S2Aoeq9zx6GJD/k/NyneYJPqqhc1ep7hiMik8DBQV+NpDAq9vNx
ssQfaY4CS2bXRLDkdiByTFrKL/ahBAXE7p8BWo7TcVK6fkVAOBTuViSpStJgCUEawDCTO8jB4oTK
LW9SN2bthMuo+aVS08Os9WdsLVAGwX7Y5ywiBSDHwsk0eFZHWdctCkfyFWBdVSYmMvr7i6PZX41N
EXmNpY+vBcO7oyPHomS03ToamuBdpB4K0Pzo10a9FoXFJxb1PslPddfSHs08za+DhjJvaH47QpHu
DCaQFR08a5Fhg99Z1K9ND5w2VyyeVmz2tow5PxW/B24dbDk1/Uu1qCUj7rbgTmalYAtg/MvD3aqy
qjQXiz7MelBm8LjOyQrPTQX7c301tbwHAwVs8i8LAtKdqLbTjMQJzElMlAlCUmlXl1j60o3bZA/A
0x4lJKJBTyR7tyBPpKSfunUi5SttNyHlqDlBaHo00a3B9sasSdUd9JVKO+HWLmJqr0fPQXp+uKNm
5K9FQlEyC7Iqh8basDzWXtuRy457jUCIDXIY9sFVtRW/AHJ6AKt4NVb3d3kreQlqa0+XE7qTJTmW
x3BDFbd6gSfd009awUIMJuK9UwPYy9/wEhxGQyTPjbGcLXugFIgN+EzngIXXMXNejKE8WhjMNQ4z
L74CFJ2lE2yLy2w7dkQdjGMvIHGGI/ETONoDNqPca/dT3vgOgzDB/P8aBL6vHgbjeWBg4GHCrh1o
4/6Jkcx5dUrSBJlRci2l33NPB6uYIZX6cAIygxXxpVVUmZRiVKpIfFSMQQi++MD0Of6Oo6AWmuzq
/6bkoSwX9NOXFbyjDLwPAHels7l1YwpaAskvXkgv4b44XhaTk9AzrN7KHEWXChLyAVAPvu4C0Ak3
ncWTa8iYt07JrLKd7iSoKM4eVB6R+HDK1LzTt2fk2TARad4lvalE1egqAMWunLA5/kcFumgH/295
VxWdG1RGud6X6Pm2/HD9l3VQuBXqCJkx2prXcNPMBOHoFwiET/6U5pARR9l66KHmu6iNL//TvRCp
7CL+Wf61qagUAflOMLCaBuE+HJuXJVWAY+TQrMF9TFr/GXDkEqbF4zb6FX5LUVJkFTLv6+7oJRoo
wMqGi+cp9PqHQdxS5NbKf4M66zgShQApLH1BCtDp6qgHOWeL/eK2zg62GfLRNntt2TKxy8q8gO6Z
ad4UrVVAllVBMk5inDnM0ML0euO0nS+DwFeMN4KdKuPeQHb3w5Q0y0DwjTz3774wV9At1RJNCjFr
Bxy3hhAzODJaubXxy/y3D7J6yVpPmubHRNH5kq7xOlJKyTvhDPNyIE0iwHFptmlndyTrwZlBBQO7
cBVhNBRmY6TYSfj4KiMQyoNJY3oiGxm8oSX98DG3x4gOHJXPdJ9yE7AAMwEWnOiu/zIB+W+MrB6h
2LHfXWYqKRh82Tghv/0e70mPHJh3Xm3CXP/vaKdgBVmgggDyPc7rSQqsoln4tT0nOKUaQIbnS4rR
T+WCEUZU1Zb7OpWWYQI79f+kor1J8u5GZYW0f8FQHDW+hS64eHOap9vKc9oxpEvq8JROHJ2ChL4k
RoDJmwHQxFbA+ghuL5+Ws5iP+c9JsQtxIinVgL4Qw1ZlgV7L6ljMNR/A1x2SXcfMsnDQFGNtTRo1
5Dl9TIC+CmqkfleXmXD7NBLlohEVekC3/F+fq2PzTbqzj9uaXdW3vRcvDGYQdMoqC0UrLnbuuvUV
2ZXNAHKdMmmvSkXKr1mxOk/SiWJUdzFf2AklRRfSP6OgC/ZBKtOAcGTUeM36I4cZfxdgkKGcMq6e
EdY4CFyCcW+yAFrCG31WvXi2T+6L3xm5DVsDUj5dka2hW5q56tWuKLY7mSgtZ6F5+MbicY/qfgnJ
bmz7WZj0nPeWe6HQAnDUeuB74y3qLyDc9LNbHCxTs+ZdfpShhZ1nyBpRx8dQZ6Q8BCTcjH62ubnC
yMIVbBI361bvJs6LC5g8Hp7m8VeNshEz7r/gKZqygR3XeIZKDvxz5jBGQQwOEK7/fr6VQm17QHap
6i/ChjQ2wpXeBDvBXIcAy6Da3DM74luBEsRL47LXMvDIp8jN/y7CTjUKRvy6Mmu0XX2lyp6nyeZF
H6Jq5XZ9yUmgxgRXMxkENl05yg/sb1mEpG2RIfgc9ufFzcg/MNmATxmhueeRl0bpqHzw7NWBIG4v
M38moIlyK6AM3/WLjqM4/rtLhtcpl1TQWJG6BN3JWstvf0gez7rU8KVfkpKMUbXqBxEibFJV4qBz
ymkS4QYbbK5bdxsLDvDgWhsauBtqd2fKZrbrS67q5l5VDvMkWFYcXl3LClbc4N3iX2TwHcSKc8tr
D/sAALn09eizKNewhlJ6OFceJNoW28Ufi4wgxLzIpBT1gAlH2dWfmZSdcJJEv14I/KSD3Kooqz/Z
JaKEEknYY4Ig3Q9D9JGnH64al5VMp1LJkVsKf6YIOVxeozfmqRLH9vLz66JHe6Hm4XDCd2cUfMqN
6+6Kw2zUzRQu9j8JDqPWHvNYBvLNNRO9LApI/f8oGJdaHikCZwY9Iaxsfu+ohWUtgiR9L/3SUq52
eVu6k39Y0SskRwIH3FOL9C8ZaClRT7XM7kl2e7QEXa/vP/Y1cbDmYJRRcUg31I9rQwq5pyoh+zGk
pZ1DPmH0OreU0HCCf4rkM/tCbNxOjz4izRDxrS8jp1SVcYQZCK22JVWdcTPITFIgMXNUxlJQ+SfA
vW9vqKwN8fwKFWNYqdy47d0bPxXfS21lWrLSRQpG6y73mVfGb6orzuy2a3dwXifdfEIBLfDcZQrp
IL43v1yTcfz4zHOhTAU1JknqTp/jicLR48x8n+IeG2plCEYvbKH/K0NY2om8DmB+cpKP2URbAp6y
zlNlR9GjDCW75YArS54K2mhGWUbTaPDqwswAkPcdPh66hefkE4sMoBvOaMoTWMvm5LRmzpLw77dk
Df9QPn9BmrlsBThC1XqnSd99MAcZDSJlltfIHjodbHuKeb+1ie8JJE9pClweX2cD1RZduoUU3+O0
SIGrnab5rPqCqc6rNVXzxcuUWHQCfI1F2xVRfvaVRCNhHj8oB+DlN707S5DBPYf+VoXFP5egSb8h
gHxgWn1XUSvAtXf9XEwEf6ZqiuU+qnOGqqccGOK2uLJcGM5OptTQ/Gz0MSbpJdl6V7Di88Ac89EI
YaZaVx0gSOA42Jv1ZJui8QrBOR+xMGmE4abKokrX/+r/6swwY1tugVvYLkvQJ+rpUQvpBXcxSLf6
3EVtAAAKjouoO7p6+f2+XKIQmaU8h2mo2Y3bMbcclhvsOlq3mACusDKIkTJ9OcdwD+fFArrVx9af
waDg9/BstzYh2mkFHFudmwLzTFSwmsVLoIfoVDBTcFMDBpKdOfJWdbb26vRzi9q6ND7Lv87ymzcn
vBRsd1JV3O3XG+HgVqSmHfNrBvDijKFS61d8BSsjVszP7YfaOZDzY+BNfaja3SrhgRXr65FpmJOz
LMM7YcKpVqePu64YKXno0wLNeP528QG6pa8bhe+jAphe+5hoocdfoSipOFkyB11yxQe5URoS2pCP
j67+NwkLpRiAFRAp7HE6F4Hx8IRmYsF15EgCRhk38E+lZC91u0q57bbw/q/MsqFm1+PXBAz23gBz
20x52cnXcclBxQPPP0WjJGf4eaR3+rANqQ3c5G0dnx0IjBlKbrg++KBuGELSMqiEEzVwf5ZUMR59
I7Smgkj4WKnVTIwfqKecm9oMEEklXYPLhgFS3XS/V/jD225i6yzaQQgHtwv2gCFDFQtfUY876DB9
uZPNMW2yam3JPDEeV0YsmggaFytum0Pf7PQwRaAMQFoaMdy/Y3n4Acdc25/yaloO7awT5M95qcIY
gY0LW6FuaPlYy1n/db6BivhAY8LTfGGYucm0E4Co8luuPylr4qlfqY+Xn3/AL7Cr/b8hUYA8aapm
ZYfZ7l6sJC6EKn8ig5yW2CKdRS3vk4QBVwDQyLDczNq9yKjlzYLxzSNt08+2F3Ifn0dbdM27WWPv
CWx67zd+ToVHRrSKyXJjwMDC2OASjMpFAT65Ne0Am77vtBAAeRLePg3zNwvhSumT+PwG5FfZkLk8
3CzbWi9Fk7Er/KXlU2pNQut2hwhq15Um5CBsLOWa4TBiO6lhc0RDqJQw8JYNtjzqFqJUnhk+ZwLd
lNQmhseMRL+/7XjzgpE1mLJeEYT+oaFz/8P6DmgauXxtDarB+N4AS6sUtGH9j/q+DYQHeAwALGSJ
F3gqOJRPk/HAQoizfZ7zo7Hj2VbQRQF2T38/dUP+DTh4ac5mDbee1WEok/6w5G6PDz49nY1VyuQs
TGXvSUYed8dTYQllkyLlMXeSQHwrTQXgw2VottF0tv7GvnENF/B5Nr8jL3U+GG3wJkVzXSzDwzSd
9HJphtE2WJlkqTCvkzLVZiIrAPxjDMmdbLSXYZVuiszuW0ra/Ol+WBppG+A4jKgt2wB4Lxfs9Inh
ngkvH7A3QCPOiz2n8bqtKVN+zU6PrXzY0MbqiOeoVSDZu5uZCM8oSXonKJ2fPJyoAp5vuezbsyL9
CWf/adWpozo8kLABfgFWfNbggob0LWwOZf3q3BTuYzD+sYAdcwaeOek9HQkQWW+p1efnW8JSYaN4
wspmfECqb7IwsH2UtTLNcg7Rc0m2a3oXETinzz6nHqzuLp3akdqg6Hy8sYBVGPixn2jVXKNQXchP
p8S3EpTvLKa3BZeG7f6nGqHxBEM8tWCpB2tSv85t9I5Yo0hK4cj7x0qdYTQcspEptT01PelHaXGZ
B7svhu/a9lV+T1tOFQrA6EYTXyXkY+vcxYPCyiz13A7u9O0aKHIGfwQ47191ErRvo61oZqI1izqB
G2T1YeWXE93t6HT1imxMX7wsZKO+bH75reIVhpj4JrC12XziodZiD5qfcHHgdKPGpb/gpDW75ddr
qSqwsSBc06NT1UVFVWs8VRdBIYXs/ndPtATNzyMKvxaSDtr9vBUHMYOab6vlVQMb5jWq5TqaK/G3
E7cAE7sHYArlV65xlVwaTUlHjG3VEbJlz1URKzSZs1CDeAT7uzAJyiq1hwnL0mUwF8Q2S8mzlQt1
vb1NV/fXKtbUnNpRTx3U63Duu+UWqB3fnE9j2Z02rLG/u7bhPkrt+kgdqZqUGExSmgfAPUV0ELA6
QCvfeGQ9fAD743ZBJR+fHMh7HPrriU7ENaqslo4hgOL/PASN2OCVqIpqhk9uXpaFWSW9AS1DJwSA
/OYGeRfNK6ihTGMnwdA1R10MzAJqf525LQ5Usm0qlcnJ9toM/4s8Uz4uVE8aAr9QNnCdF7QcDC6g
Lzt/YK/VuwbVi8CvEMHvG6drHujB0RbGDGJc+dKGkUnvi6ON+CcTCl2d3X+RM3gpscYTXk9UFVR+
RuzxhshJoQ9RKzS7VronbnIuU8JqYn6Srv+b3gIhuUCK2qg8lii6DsGrwtSA+XSMMHNP1gHf4ork
M86S1ztSfI3j34lG2VmFGI/QbWby87Cs0z4LXwniH/fDzpF8Mx9w9AfeYHrfQYFOH1NQKCbXjGLl
0BaLDXLVpTdfNzCfCeQnunVDipurlWUEFiUfcqpGLD8qkkSmj9MFoSbETLDBIfQlGH/vNXZs5GF5
m7j1O8w0WCi7EeSRFlVQsivd+8gBPLuz2XadDNOraoPxt0jD5so4lJOnrhLxcnQpPuk5icULlwQ5
XgGA+w/dJq/EzpEKCCkB/yAUKUU1vEb132mfWF3dTQUeB4JclexnUKS1Em4V+m0/87sAm5DgZxWa
P7jwZFoWlQ/nAKy14UECcNxxCZ27IGqhYc1PF7ItgObGMFQaQ196fVVJdE4/qfXvlqn1KYbx5KCp
yrMkP6tZNQBGmg3aGy9Tzt8i0XFP67nedhAHvazS/SRHqFUIyVzX+91Cqv9PkYLvPeN3oJT+FZmt
u5nhl8w/WAMmim6rfKz7FikLw7ouA5uBbdMTqSVTaePb0nsniX8Ohhqu8Gf/WD/hZEFwOvhB/V37
EU9LOMNTlJkOpH3EieeCl7GhyqQqnyPhyFV3rju9vLggnoIICH2CmtT4kWSu+nbWUvasYYYEL7PM
4aCWd/RzMQ/fKo08HJhYW1J5p5Ji0xYRp3gmU6Hsxn9ipXdAFo6F2x4Pt+js/wHo4vSyHhwva+km
fJh6ke7L9MVNe2l8IG8AWF5a9GmStO7JARqSANsjvNkNVIBxHzX81Rjn3hxDQEt3If+0awxYI2Mz
os0+q8kG+GHMwLeKbCes/AxTJhf60c5L35gFBVzAzi5XPZHeLDxSGAJypJxf9m6q4TNWjH1+Iqm6
EfnEbbokUIlO7mTJ0DiZzpnQhygAword8H8bSMCYGN46r47BNanrQLL5Z8soBmchdLc7sIZ4a6nw
DzCHRvlofmGB0fTlUtY13jcBip/9NSbYHEAXSUJGNiljvIXuGvvWRqRcF3OumVAFi2CNVgUDtIzU
RlqGhRjWx4zDd67Pu0FYZxrQL8GpAiUm+dRzneHqHaVlQaMY/EyyLsHHuOkaznWUz/QMJ05HnZy6
r9RR9fIAODbyTal42ujgSLSy4BAcmqnX46N8ud5OWweyHOO4cxTgizw8qzdgQ4j4vx46x3fSV3yg
MTYlCZyBWw2VU29cfaJCZ7gTwX9yYaqUxzOF/aPiYiL+Vb3Bo0j/L7sygkCnaGIjAMweTSrnG4+q
4uNSvkNgx2lTIwXtxr9pRFEJoWYA+/1f4mU7MJFTbJR9C0AUSfK06MsdKj7Xx3z62Ve46Jzc69AR
vEV1/ADi8ZQnSXOZCbDGtr8jHi5Fpcssb3V+5Eay/Aq6/BD4JZ6+zxncq6XwWRPaD96045OWfmqo
uInAhys4LRbzOZkPwJSIKSOIB5xyjoCeXn54VPJT4FFiatAs39B4JwyFoBsZSauWkPB9mEfoGVN7
99CZGOyYHxRtNPrHRkE/tu2LyxqOsBMjjy9TTsl//F2ePv0dWAP++6nT5Q6506MosX+3806Li1GM
3W1bWqqCD0DUjbpcYti0DYVoPiUqgoa6YKnJLs06sgHcBsQd+1YPbuEJTFqIWud11dyIFd0hk0Oj
1mTRUn6+UlPzhoBBx5H14nsKSNXLVD+FsAO3aStq1aJYyAH1E/KOowQ8TApK0g2a5ek4uWhq5/+p
EDk0owknOmepV6WxVvhVB4c18ZiZcQexNNvWFuUWDhnIdRJusTqjdNGZotrTDkEfzt5Y1E3dtRPe
2vpgNW+GrJQVNhpGdwXzWyV5HGVjfoqoCnfd4XYtBhQzkyMjaediVqgBHM9eEccnftkdV3vcULMk
A8iV5GlutWpbmxr0utzARmA52gUbH/ftKzy51y7G1fBFb6H5nKaM1+Fn0dV0CxBVwz3OONiVR1cY
qTsj29tK+USeCex4DwRyF0m9flm2eYwIdiIFAVJUw84PkBw3N55mIol2X7veHNuzwmA4SUrHzFCI
UfKJUtkQ0bngOAAyORHarNSYkKEYSu4fpoXwlQIRKkJPkbZSFFjiSsU+PjGJuy3BvcXxG8bZLH+h
ELyu16JWHP+oncx1yXeUB5+kXyRoYB3CZ2m51gjLGQq0FKGh785j92tmBj1z5gQoB0qVEgli0RUn
/z9SwEDaw9YtUpDZsSMf3BflVcmt4fMLYYAuo/5sItjnrEoe4G4GLIUveWUvlYPsUKXlXQTdqSoJ
HxO6FfWAU9ljyQtzq1jD7G6XVrCttvOqRbPBdqWqErtavJk++MfYKRAVJGZTEVkiHdBNpV+UfTt1
Vd+tg7sVyfeYHeGpEnyG3SC8hj6ZnxyVbhtmO3EMxne3y8bblHdTpZsns1gmzqxXkEd0xUbKXrJw
ebVgcaGzwXU3KyqWDriNyk0H79s4XSKcOj4iBhebYjvb5K2i3Jbz7zuunMqsUXZCcAMHrlBYA4Sf
UHNzLoro3EZKnNJ6nYZ109CZBbM8WO1PX+JcedLr8xS9kpA7/l4iDK5h6a1o83aJBTITHCZ1unPJ
2s4Lyq8TRN1RM2CxEPTayly5C4Ch7oXZoOyYa42xXFYjtSE6pg26RCzYgQahO7DUS2cH0cBV3jDq
urBoxT0uS85IRUGcmDUSkhUbG2NetS941vvpX6MAlFj4OA1xkoOw+NJAsT60kOkiq0e+SEfvIDlw
6RJ+oJNsVNKJGyAK9adRZMDgY+jYslFPLqV73/F5aA5oJjDXW6yX4HNuoJUXKHY6ZITmQI+4CtZM
04r+Rw+H/Aj5b7b4JluVoTs7T9o+PMIQ0LejLOOEa7lXwCJdtNl9IuAkLjSfZnHLutojIzuKpmSf
hEko4uE1zEr0WAaXwyJ5Y1h+S7QGsl2E2Kf6BAAIJsW0VAnVAGBagakce+AV/9R0+Iv+7fIX9iPL
IWioga3ijiAFB1cQlDtsQz8A8ixY23jgvKS6ReBmorfWSd/G4Plxft3AyomoHA4+tzXDacmweI6A
Svj99O0A/oAmkIqZ5A24OFbUue6WZOmbB1P951wCUHbDpTd0tjnDP1+jEh5IjHlB/fLBarKFnfFW
Inm/Od7F2DE2eHFu5etUtkIxQ1ijC1zaBorgz7UcDY7xc3BZKkggrVHKG8uRe20Zm59bRBteYRhy
TWbK/N5Qtt5Wh09lOmK34RPM8v8eL+gyuRduN36dPRITt7xjVShQCdQ/uSviubf5m0qrA1+5Id2s
D7dwVwnzkVH952Dj/N1zYJOYirYP+OlIV8uQ1cuxXUmxZ9k6oHr1ORNqR4EsPIrXQjV7dxYapBQ5
4YbB7XzZcsxJH1x7O0PSzs7rKRSYSpinMQxNWcT8gfLFaiiyxbpy+4TzBV3y3tklDdjiF56WKh7Y
BReCaJnHhhgFqGNnZqJu+wdywLuZU0oEqirTuxd8j/nCBC5eNvuicxaWoFTxEfGq+iQXukw+LcFG
6wzMg4lLb67KTM4f4ejbtFiGL/g+fgNr+e/0EbLLjkCtEfPT93GQYAe6TGzK3RGU4+bg6m4EJElW
YcE1JaH2n8OsdSgGB6gcktHf8E6AZTaBAA31ej/ga0rOXvz0NPuAavUat+azsgoI4w0UsnzWj65K
V/SulnERSpkdFPGVdd+J236g8dtb5b6liMNyQzOksTf9lXHsCQO7IVC5utctxevzx1lAWAdCR68i
R9joGAOTBl13L+QLo77siJvMxMHBOf+KRobrxlbbaPfwt7Wv/axF5xYwBdBWtplZ9eC0h1kM2xe2
VziJ2woXBTwxpmKH9Xvzpm0UEL/1CeEeFcyDQDCVE3oU04Tp4lrO/2+BDRC4b7AgTHldMCvHDvS+
17BdWWBeYc+N1i9z15HaG5K/6LoupV30RVxk5XAW7ji7rzMRGQU0007FCzmbNcXWaggdUbEacXkT
4CXwkiVShsoUuIx5hV55/j6u+TtbP1fUpPBjuTP5huqBF59kQSN1wvSfCUKR17CHiSpD1FXIVvuC
ZN2RbjXgxebHAD/KuPze1r5ijsMOhPNx1UKhlfFbfC9/2JpD0EMkY70mZBzK6hzlNVKk8p1kB1Wh
NsweRDxDmLSFUVWXkIu14MSlFnkL+DHcvYOgRq1W3lPZ1Cfh8E9uu+wallXEtoXPVjOn5HqcCAgz
SiEmCNLiAJ3cs3lMq4CKTvdCP97OHcON8DGeB4qvOTGB0zV9frupsV4tNNf54OhZGmwnn+ilY7y/
aZyzEHRHARWAotx+TVbxkpU7VFk8AuhvoKPDEDIRsxp2ibqzFRnfTPsOiHFJWiTK0OepuTddhyBn
7prYsls2ck5R5KQ0RJAw9xJbuJ6BXdBpEwsMs3FMIL+BFXE86UXMIUd3GaZVwYRLs1eXpHqWl+VW
4S46nkGyGbgeeBJv/v1b23rSaLVy7CzsPvfruks8bFi3Br3WyY9UCURYbcO3fJvYGxizRV6cwO86
62nnGfkKBAD9kOAIrqR4Kg+VW9kdwFx+NMNho5w46+Y/DB3+l+DSdcYHoJgJX0eASXZFGUlDhLDf
zO4KBKAOVr+d1JzVQZgOjhkDtHf1afYWmCPDJQFVt+6134oS/exUU9LW//9XWa8aUt7pGriYdtVY
TjiboMDOkFJZxP2rhrbW0ozKvAOktbvCiWpudurccE1f2Lcm4AJ4pm7THVaz++iFAVTBYw9V1ap7
3PhC2BOxbDsudPY/pD3hvkDo9eXnXkunggL8Vo0STBGeMXRdnRK0c1/LEruOk8L5nBz4ebfi+U1I
HcepntfqFDARsI9K+SVo48f0qGyUZrUZ6w2warxKSuCRc7PPh+qAITRacgUxkjIfg/mDqM47boGL
Zmnb4VtxVarzb36WxpN9cL39OcLlR+b03hsarh9HQGbTjiOalN5OFWAb9AB8zZl+qFQ5XSRxejmF
QhoaeVn9Lmv50kkPe9Js7SOAQZmwbMrEQmHgFI/iAQmWMtsrLCxkJjO76sdl0vcWvucJjhRCR06c
V+nbQBQi3FW6nm1cE8hn6XEUpYL6JTmkY2aEof6scLa3NwMpEm9Wm4rYqZAVZZs1Mk5lGo3N+9vw
wJ+nKd3rOkyCeqBIYDUOy5WUvr76MW3lD8ES5HX41srTG0D4dVPzmxo8c0Xe8FcN2GdnW33p88A/
UGdfQSsMz/YL1ss98LNGvESFUHJz+/SQpoLnlR3SdTz8r9S+MuTQEz/lToT/qt1PA+EMcylQhSSC
lBtCQMVHg5PX+1FpxVayRiWcHGSvFsm5w38a4uw3hoM3mrXzZnIXq3bdp+oG+0gI/oR1xdrSOtCA
pztyqfn2+MRct0eP8LNeo08GUfSwpCLQF1P9/k93P9MsHdtRlbgZ1zEvy5s0xqg72BP71tzUdOix
000/pHUj6PU09eIi46fIqcMfr5xmtjJFg2HHOy/vR6SdZdH8zoRm5hlkewSAcsgVjRNQSlubmZOs
5lLZ4L8Xp2YyPSP7LVXYIgQ9T+DpdmYUA+DoYXKtBX0sDL8z2oscRCcTnMmeDRk1EdnqvDYp3cJF
XzO817GcfrGuOUXSCciqYShpMe5tuvvnsOI1iRqr+uaPp0+buGi/Z9tWIwwVsVrmGb+MscFW9J35
OVkP7JBcI5ekBK588EKNLxGLMV/X2Hj2LL/OqTbCXSBxX4PrOWUARKrzA8vCzxo+W5Bwq4FaBCsB
9UatiFq2FOee+Pe50nX8AW7U/MWzTVIS7FnNhABi7Pj4VdRtIiBCljzsw96iWuvo/7EsDcPIqJHH
jAamTBTPCoAwPAsWc9KeLaYisvnQb5jg08nc8/IyxnlljEWGLKPgktRSd/yvHfWCkU4L4JW51TuZ
iqMEwADvSNTmU8oeHi5x5OUCL3xrspv4Tb3bs01VIQxQwuyw+ogurKCsaDXdmAptze2rZqjCNKs4
UHWTpOCQo7sMAa5J1AfCspd5nmp8nzrHhJpZM4rfIZZk6t1xCkMMRFOaqQtQOm9brD7GUK+cKObM
OqQ65eiQZb8gja0fjZpj/NDO3m0+OkLLtZIVb8jZYINreNFyHuKnN+K0kazijsujRZNPBdt1Evu0
bRxr1U2rtrMDOPd0d/d256psbC7E0kLTfPIIhnBAGuii9EAzOhFQBJ4Ey7Hf8eZCcwAomdJDKjKj
juuCMBDTrOau3FyedYEljvxf/+Q/TntK8H02lls3mMtRoKQe0IF7LV+wNKPSRoWzJW3aPXO5rPOD
eaCdnOyUbUNBxiCm4gGUqSNDpLbmYuCb22Mrx4YAetAGr4x2YUX/+uXTD9HFZnspkAnQUSkAKRMh
phVvm7JhW5nnxJVlbGWFAjGIYc0dBuNMCDfKqqcAKTmeagcCyCyEMYlrYLqZidLyHw3a8akjXdF3
UnE2hJqt+eE+sLLkHUiR44B8MJ+V9ZMG1wrengKmDF+y4zDxTWFLB+B2AGU/mAbqslSsIO9oVQlB
gpUYKlFemhQIBGERwmbpz4rELOIzHHQxhkCxQ+A4ykBGGpSYFsh0v2jn11/iz50Td0DekFbyMy0i
43DnUl9Gxq2Z/IYIof1w1d30B7S6Rvetd9qajdEuZt31/zb93byLKXFjEL9X0AcgxwYQ8Ajv7/fs
NJmp7FQ/f64hnhk4gjCRDgCcc6ijAgV8SWk+2If2W/Li1MsZGQBaZFAAqBKw2OIDyISATDfHRVVd
EaKRqYyvr+QhGmXWStESjO6bRVjS4ehEOeATzGwrh1f3bgErV6dOk9qaHwQas11dRsdleTlCLATk
heIhVu+StyU6gShKCrrrWyAeZtpuWRVIyTsHJQgAnegpqbQzyT1pfXhcTRLfPCSU/4rQWZNUyo+y
lzeV5QBTSTKV0ENiHSMGg5cLHfYOs1mwmMOYkj1meM7nztP/SQJGvsjVxXZPokzYtx/ADZovI1G3
DrtkFVTI0ag8hVewY4yDRT12BLpwZhcnf2MZxSHAC08L7570+oHE77sTvKVwxfZoHdP/opi+XrEW
ZGWKmfNwaKw5r2maZI4vI6kfsn4YvY9Ei137kvXxgFfixcWEKsCRC3UkqkUfL+/nFrFtSV0VUDU+
jI9hOyACIH9LHD6ry91Dn7k2G36Q2tXAgU4OBElbLORTT3ETZHEk6VpPDUfP3B75C7jr5uwhA99U
K9+g257UEK6h4t/SMwlqKAaXVV28uByE8GE7ljauSA/JkzAB1OPWXRx8EcF47R/QEgZONAjdETPC
fsiZmZdZIS+oowc+xR0RKKYGjgRaZ1SWO9ST/PLIrg2IDyphS6D2zgZqtAjZV/RmsNGSr7qbsj5n
GRqUvunV6a6phVTbd0nVZ6mL73Y4nnfbNUHE7CxoHuSxiDyCTUVWmPCAwXRIos8d1CesC94xc3oF
pX6x1B0pptpXrbHoKKW4FFs5sf9fS4cfew3x5XABAzcgzBDCRVDeVQwDTIJ6zNw0Ipp9SzfupMW1
VAG/Mb7DTOrZOpxXcb7zvZz/bz/exz/93Fbn0aXzAaWli68hSngTEWSm2iErdHINEiGLKnF7d4C6
kGPI+sjakShU+fIuDdpPzziCmuntCuyTsdUiffJdiIOgjAvxWey3IRJqQaFWMRiCCFV4CoHPagWv
OVFckSm5lfD8CtvAIbDjBxfkTKfruhf6Ju/ZDlO0M/msiUc+Z2eSTpN5QN//P7Cr9nuOCij9NuSZ
bxwZrm89zwNxeAKbLn4/nCa7DOK6TdxYQZK9MoXMzOXavysKXBmcKfyAchqvHhjObxgwtELunHh+
rnglmHyD/zP61vH5JJOgcKF5WMVm29cCC6/GIvsPbqQGJuS1jRl8XP6aDraSoc8NtEk8HEfLU89r
vBiLI5d1OsCGP3fS55FqUBTTWyFCJDmywd53Yw4AcfYmZvS0UFUz+USsVy3M5v3HwZQ+OhNE/WjG
AM+bQ+jQarWaMZh9sxsUP36sAMLgOV/+Oqb6STlHbM5NRFPgqLzWr/cyrIczrRIl4CBtywD9qlvn
mfyuAhLRy9hikNcE8VtQMakLGxhzMNNClASuElCZq0g0IsyhNqbknnsZysHqkLC2GAgexLJh+Qyc
50cSjP9U8EUecOCouZYP+V5hlKHqu11gXnEzJF6rbxs7rLrfB2sryzdzy06WOMvhj/1CJiFjHo2l
BoUn+zc7xLEJHryxBycdetVRWAV64ljhh7XU//LNHcxYzPI8WlWDLwhqsCHum1D+nxUkSPOKvUrO
DntB21vlU/WEr3hQKoC5YnfYAhkrJIUEle7IFBF3B/WiHpDfI6xLX2+cgnBIcZHtJw9CMWFpIuEV
pNSwloG7euVrkrMNYbhUGK+i4GEjMMruTvMhe9W0OoRyOcCGMOyZlU0o1c9F3XWlHnBpu41kVkYX
E8mp+g9A8mmzxqQAcvWzk4silGkhJCalBkTqbCOgV7eUNL5N/2OnIKMTMPmPiv7yR8BUhpWlHEKO
17isI8OI1i/DdySJtkDfFCqokE0KYNbd4xhjNMriRYkeZF9ok6TR4pFyWiuWMi4yWh330Er96Wz0
Ku03AHcvX+AeelbHXcDqSrKvZfwPIvTs/mbLp/Bk94zg1vlN0TC5AGBnTO3Evnb551emeoLzmUR6
CeNjAwxTESCYKKbGvaHZfhHuONJzEMoimFrimN4gwpfcYUIgbaLqVPqp8fVboDWoLTnUrg3Ng+r+
qgoK7yNdbyxgxSN634BPaGOITMVDzAq1qHer1GtYZbCnfEqxzBerEyrdVDRVglk0tDBV5eMlJsBp
tqZOV/UOt76Q6HtkV0kC6pqDdtoKmKzyEM12rXdZ/LZ5OdY7MXcnBfjokLvM5PvIUL3Eoeh76mYC
CJ5HlpyyICfrcBNpOScUmXZ7htGc+2Ga/wpVmm/YoDWZoJwutiHPC1p9Jy9Rc/jq4O2c1DxpjYUE
ttQGBx45zU6MgFhojUfF7O9EtL8AJxSl6VTg/YHl1VG9bDobWrN9QY/H/vJfMPQBOWt1Bd5A4dNc
jKUMlpVVu3nh1zlr83poh+SpIwC+DUgr6Fjg0jIWw1Jza9LSAkhx9a9Q/Wr+LAjXWWdx948lxe+/
Go5/3313l71x1bLB4lk3YqzSgeHDdwI0xijeY/EROfLVHe3lZiFJ+drhh7fG8FHlBi5dTJu+6BEG
9myF8fHzpuG5kIccYiCsGusUSKHck0ssfdQEYE8JtEzxMTTY/9Fe5MOA5ml5ZwIPsuWPvttRlQYf
k4cO+lFpkTjT6lncJtZTxLigT9zq+uhMU6IvLGGWwc4UmegsDBONkqoH1K9Ai9FBE+fNrmVuRjgR
MkJDPZcQdN8F0o99p2J1MWLHJ31XgdD0UwAcs1nyYynkyO1dVLAkPAZUp8r0zQzswhAOx4qFH8QW
+wTIXc+JWEFIIuCpSv9A3rZ70h3vIxk5Cz6o5v7ptBBueMnFQNY8189KGlzY+lIqD2GR5zqjAG2U
nUOKeu6zeyvHtKYRNqYeEoQauAzpoFBGhmnBzC6QkWWDFaDTSR/UVvRqLAbQSXDqkQ/58Iw0sGVM
iWqppqeEdjmSez+nwMLjHRLiPiCyoMryVU5KSAYsMQp9HA7syc/t8VFCRIunn2kG/JhKTM1/V9Z2
+Op/ldQ9q8vw+M93o/ZCEJUYm4y2ys/zgWKYp+/LJth0n1EjOtrAh4pQmXnr2Wx13DhT5NLPpY1o
dCh7TCg88HjvB9GMTEIGA2GZ9E0N1zpn6MjpeNjD/X6xtohFSf615FANUZPwTfQJYRBooxTotsvA
ZVZLcSuEGuAWmTBYfBk02FurAFNAPFnWHNCXl0z0h8jUD3neDdstXvgEqS4XIUge9lYSAAs2sWZ+
LuxYDzdAxQ8j6njLBhkcxayXYyS51ar7dCp6pg349NJRXY+t01ine+eU4lt+yo/v5SgTWMnoatab
Kxd9XAEY9fAwuG54CgwL2HyPxRn+cBqfblc4BLiKWbLJuOGyshtR8iQ/Cqs1qFy6jIna9yodWJo5
TYN7FfjxRIaagHj3y/kFtIrOJE4ZEac7L/0lA6xwCHZc7qDrxOCIGk+LagbNDTuDler8oTW0z6hl
Kr/4KwV/tDFyskBSQrpxbD+u8Lm3ApeEpkQdfewwUvxVYIh9R6h4EcdzIn4KkQPVPNts+goTN5Qo
jq22yFx2dCw1S+XehIrKRqX2HNyDpUw/gHMcL+D+r5kKEpsohpJImT/VNh9WHMs69nR4AL9CSGPs
Mi/dvozwv8lWkFnZUFuiPdwod3bbuMAj9uWGsalL1R/fZS/+VLE0U8PoZW9XFXMT47QBcBRjRZUo
pg+P2CJsWzZsOdkK+CriyFH3YdLvHdjXBTjbULSkHbrwqLCmKEtNSyw5fmjLKi37dIPADVVuLtzI
re4gellQ2zq3J/Yvo8QVKJVh7K7CnKY67uk3GQohwz4lunh7SOWxF45603GsPwtE5R/9U+9M/0cC
sElx42uQLw6dYP03QTyTc+TR4GAX0fz62cjj2Dg+vLe2/cUwKx4Toc22Ju/uYJUQV4Y1xVgTycbK
PG3TqCVlPr3zuTv7wXxkbZDUlwsvU6RzvziwtOzKCQ+/PLqTHmDT8RvY+wTfIj9cvM+xjT+UDFYC
3JaT2ry8haL7kWyv9OgKuzEHcSCD65t76O1+6p6dLGthiAcswVniwjhyR5hrEvvN/c/ciWaOhJdW
oLkiExVs/cYyfcgTZfOYbQ7hZ5NtZMgRSUehHeOphh+xvsQoTxk1f25X/0hOUgnShGc426tvXIVh
E5/sPjMyUsSADKGqIL4TVkkQO9DUZ3bPcHq4ZSQfQTuDXnv8WvVlao8hdYapIFRMYs+pL80gkp/p
0pUOBI8taj2PO8suB2GIMioqy7blF8fwWd8jINFyxpTPAfzcFNj9Q2jxBkD56yr6Ka5jvXYy0K+Q
XosZud0KknJnhnqGB4uf9XBdHhY5zm3rjhMeWIROTu6WaqzbCN4iNbbBgzxpLVxFYzp1bCkV3xKn
RjYCP0OStYN/oHx0F4heFejTs5z3aMsn61phZZDTnUJ4rMR8FTypXGlmB0UUXIyTClWgx8M0XoWW
hlKa86677anDIIYbJuSQ82EdwHgAVPdJV1ekJaWkOmuBkCCtuxnQ8iCsZ+eSDiwq/h9ZEdsASmWh
bt4XcoNFlWZdT1JF4RtXoSCsDCnx9lgWJFmufg3YOPYH2wLn9W7fQIRMegVP1bmE3PkXxc+MAUZ/
uB27JCnuDuyYKIO0yutQXW95ZgJeNcHHTTqzAqf5GWTLycDFAfniyXJMvevvcefU7YY5FkF+4Oqe
XAJsO8lEc8MXQugXLMkjNn3v3b9fV5cGmTISfexcyEESxOZyBW+bXDwsw5MH/Uel/3QqOSzPvL7T
z53h+w3pg83NsaCJih4xTAJvA27yTS3I8wcjihUZuY4CRRXupgm2wxD4UsXW0el1Lvg9zUxCbs3L
k0jRK42k/oDlwLTnSCcElk0vSVlYQzcZ4ODNcvjNXz/56KH8wFda5JZB+ZB24Y05GAg5Df9YY1gM
ywg4TDwmFa2m6SFZKmEdWFKy534dYQgHpsn5ijxDzrb1epWJTHU/s6fY12e7+MZnzqCllrEFU7dI
YLWzjhckDokPd955KP8gsKzMLQTijBzeEc0020jdcFtCVIfBEi6EG9vZEWOpEHVXMGOh9eD4LfxU
fgNTI/PppocZW5wjf6tQEa/Mai+8I1AUovVjuIz1QlcUePGAPi5podMU559uXavXbUYlTk6kblLf
ha2LsubhhHMxaE6pGfw3mLcmav34W/NuaeUXwYabpKjXvgMS/kC3JbJX5dQpphIFvYDHXQpAw2Al
7nOAn4qd02aEfdjQKcAeb0o3RCOhY1k6sWy0I6IN1kg5zx+UCwdH7cVNv0BQPkaEuQl3V2FSlqO7
PdbX6vJ1FInQQrQGczXoF5O5rgEtcD3hUMFYZT0Rz8GXyxGT/vVVgjlsaMzXYi0yYJZwHEp5stcW
Pmi1Fxx8WONGekc+D3Y5E+Zhft+WMun4RvgMDdofC3Q8PSXaA0EDMZ7iDjZzwtVGqpsfG8uoIHQD
7YYwZ4uQzD5J678GmoFOP9XoW6OJ0ySNo2LH4QFsF8RMl93HNZ/HcYHWWQOgAoX1b5vTejs+VLKf
UCocr3W8TYpS6cOUoATKSUHGOOojZErLiNm99xCaVaO4Z6pqXtSF1nhIZO/uc5BdccPg5egcmTwi
fYhmZJCjz3xeQeNTR+02JtYBtOUhn3dhlfuNCX49rb6LWS1IMPbFEhQWa/iGrHJgL9PtPDvy8MSp
9ynGH9GMCd1zMpBIy2g7MqPBzNcOEoC78FCqPrdAEI7ECPEe3eYuJYPlfOBmKZvtyXjs8oYyBsTA
rO+xXx0L0iA/9JZrQ9LTSmdCE+PS7/SNcB3FZ5JNwsYJ+I6PsxrDJOACnxLmrrmTLPgm1K8znVLb
4fkm2YQpTl6TuWZZdVWS3xePkZ/sNy3CbIONR+y2+W08rHU0QxBYPwztsSyjw5eEUm4Iv5UU7ebP
pgJb4II10ZrD3FughEnWU4Y6LGPd43yMUA7UT8WTObVXR6lybcPmutdyAm8LXyws40C37547ZUOy
qhUsE5Z3EEeGx5eqpMOJYoh+PwUF3yNR70+ev5dLNMKnK8llrM8ZWEEDrGW4d71RfXFRdwx63y5R
7mlila1dgkDeY/CYxAmNb5xz0YuNZah79LCfjXtLm6EDcdBVXWNztOLn0pqQXLo+QZdpJ7kERP/5
CK6FkArdS0YlqKs8Hkwdpq78m1cfYgcAkE9T5cswj1xrecocM333IxNpoW91TARWOp0KjRBz+w2s
Y7IZ+weGHf1fpydCK01VQtrnHKgQoqRX2+/16ML3kNUcpmTMG4AyKAWRI0K2gSilWNXXlqGBYhMW
OLYpriDn5y5vcI5a03GRC9YLoA9y1bQuAhk45Z6rRD8P2PqdFSWlSXb0LZp66BQMSy9WsVF3Sxvg
Cu+jk+3my0D9xFlk8ejx1EqOfBM4J3Giir+Y5y76/XS791sae8qpSfmObA29XBg4Ow37LvrCFTCl
PGR+Jw2t4/phK1KkuaqroqEq0Dfw5+QqREdrcVUO+zoAJfDtPtKHRMmE9PLmmre7fJCLBoQODxoZ
cxzVgI+g64VxwTj2Yq2n6WWDif6JMdJ8DCQE1rFyjMLlpUYBXzW8EQTRJds3ljKDsMVtA+7Iq/xd
khdeZy3gu++2VSW92qk+n3nj8LxG9ng0i1UzoLUtPOek4UHv74lwoJW/YGGayvym6HalJNksiX7H
Q2HIHKv9ixxCzGLVvzcAAFGnb6mkSQbP4vHA36t+TnmwEIdLKYKYgptmJBYj6VteqTb/+3zLqbQa
5cyHOgxvCGa8B4TbPDEYA6lOCuhdRV/Fs/pUaE+mtKJYOVgMkJvWPwD1YN8LuzMNfIHG53tNNTpz
oACeXRH8WHwG2/k3stXXNtQufBCxxZuAPirfpEmUlA4QhkCdBNIvy94TqNIMWnk9uQ44Mbk/zfn0
wc4QvA+HRiUNnbcZUI8NScfNEmqRqKK3shZjeHUDQTRz1og+4QkHTsZjUEArwgMeo/Mj3+3Ze1wb
o0EbmOX2B0G/W32GNEPDnr+x12Rn80cR5JnIu79yz5NtHtYwD9D3bjQMRarzB2yS53KBosf12sWa
MGSUvEhc8VjX9GV9L00iDELDM3NroaY5kRhpo/vPl6FYgMgZwccD44M7k5xBPAMNOpHTdZKq4jOc
EL0a9elWV6O9V5RFdvRZSR6wJtc8k6RZq9bZQ9UbpkBD/rrT4DwwZ7fUYrEPqSPWWDTYdrhrGdd/
uYhNOc3SRv5lwT9vSNhA9OtKMG+saZeYxb+VyTPbVPkOux3WdGPItM09/0JX0mQJfXiTxMj9Ge5p
hRXQ10s0Dwro+A6GnBQ9Bke5X4KkJCeCnEaEbFtnlMYEY8/OrPoesokFTsHhuqUioJjNWcnszjRZ
1LQ8SkIMxGRFe32SURL5tc7xBnwW43niSCZ0I5OVNEjeggFB9AVEIxI0e1bF7gH6ddR+/zUftsu/
bEB3ZQ3Lh1jM6YDqp5FLbl2U4lHwQSu+BdzsY4jZTkXxUrELpKEk/1VumR96r4vY6xo+9MuUEGQe
/0A+5JUbk6WN5z1FL5wMeveaNSf2DZr1orz4GCIuNpvQ1uKrq3JeQZzpGDd6F/+kJMGWVfJgNXln
wwBtBoFMoS9h5CrborEVFfBzrzNRoOp1oz0hZx3vUn2yYWyWak7hlmmBZWOF//nJKCXwP/Denzsp
i5K9t6fy72NQdipzp5ul9fI+wtyjSWLav0KLbGKMWHTnvg8psfJ4FyaLVOTKbo5cXmNnSJkAyw57
V9Ak1i80Kc20dN6p2NN7zfWKO3L7DRcZg++2w1acEUDrmPxTDJ6VIJL5Lg/sQdVo1h83oCTnwx4m
9bvEtozyf4mYeU1xqqrnZNkNxa1wzd0pQOJJDhUJI55YT+SdC6+xc/1uEXkbvCtwE+5OZyyk2zvE
WMidcWrLhNc/C75+m6zO81MJAytZ8X2wE2lko4LtCKu7pqFpqaM1x7UV62zTKLgFTfH211lv87Ov
sZYPqyM+dMCtdB8VUqa3/dDMpgY/7pAwFdRxkPBhhGYMMpBrEu3DM7mNLx8isbseQr5Sx2rjplmj
TV9T559nWkBuvXKvpygPwIoXB86n66XzqOh1MJoNkFBrNHc0Yi2MfYs1dgKXDK9Wc0k/K+AkqWhg
lKcbZ4v/ILX4L2Yevg4eIIDURSFOtdoG/yMiijvLiZAMfSpeIVi4yysiFbQVL5UiiBP4muimmrQp
rhpW1xuUD2PriNKBHfTIodlZS2Xka8I6bmRjEadACI6uNfLw8uJ2JVxPqtfmkAyQSTDOZvwSz9Aa
RILJAxrw8DIwweQf7HSO/PGBcZu9Bfx0U6EzDiOPr1bMv5hei5olnIU56+KDw7sVEh69zCSvD146
KOGgCsuIPx4F7dj7wERyRfmik2J0myglNipZyLGsgHll7x6cR/i+4W7Hu6Qq62PErOmtP85K9uFd
B+8qO4CmZcLnGnHbLmR7uxih1Md7syN6d6fJikXWJE+xCTsVJTTsqGKsZ/GDvxDyG9An3UfI9C/D
+FK5yYg+CdXGAivOheFKDYYqnmAJ+7q0nHVRQ3wKvac5+5gnq01CAZ2YZqidlxA98aDGmwMDGXrL
mCxICV4IsLCV7xGPT+Nh/en7c99/rxCF4C4Nsdp3VQDIsKE7h5b9k6Jza4w7gwQTKrFIt3v/sUa7
9rusiJDHtQGoPdZpsc7hstD1usYm39DXUL1PmpxjEynNdxoeaehZ0VBIrfbecUvbIoBMXIUwBafJ
o3IpQIT9yOrrxH9sWyoJ808YETNXShR+kK7556X0xBk1KS2qj7ubi1SHvo1zoAqFnFH8LaZYC7Km
U/0bbGORlNexnjev2YgKWp5uyhPiOcnuFwJZxYrB9PdDgF/MzvKSeTN696HhEKMN5gYoguycuYde
2tplGPuJBdk3YvXApjI8hsdKGZr2pYhlren9Ctlx9+R/S+atxEzcJUuhbm2F2swnni8WxtS4Whms
jVzKdw6rjdulVBKKXp9kizp7zAeIEAYc8rjjSGbl52G+RFrCvJGIiW4slyvquR3lItUhClWPSQg7
A5k+mlJVZ5+l3I5wTKvdpX5Wt73ewjgth48Ug0N/1GGvw+qtNzcTuxuF2k7oE3KFvAEE2oOLOQrW
jx1bo3b/Njim9wZdNyB4Vpwuc+XH4gWGlkqiuozQMbQsvi0GBkuJeEBOo4xcCBvhPoVaI0n8ptal
wWwq45cBhHIPr3IKwRuAd2D4ZQxnlM0LW+WlSnaBqPvaVtEae/WjhJ8VdyZMb7n3cTTHwwpGbV/A
QzFG13P/mrZGWn5u7Z/BXcZvLVFScM4o9DmAdyZA5AViRTE6N9s7z3djKEIap00dDE/c1724CC1C
aHg32KbqjOwBSHTENlESV9psGNe3fCvpLRskJ9gLm/gmA2KhDzAMDIJkpYigmHiicMw4vrzUB0o0
k7kvOuhg3nf3AM4jLLc3iix9T2PNZFrWd7hjRnQj99TJduMIUDhhZ1tJaPVmCKqUkAZG8eBWx9Oa
id5NNLnb2uxNxRPDzKibBP/BmLBKNLhtJ3vPOQ7vgFpG8i+Oo+TdXU5tW2DIXMiHOzXD/yd7y6MO
1uE8R+t+oh77IDUp0a7gk87TDkXVFSgXHdggBpkSXCzuP1bFrDjSr1JnCW/R5u/5AExFiAWgzYuH
mWcw2661F1etoMOgPG4Iox5BkJpAaHjAdqX86iJu20Xhat39krdHRMpx5n8w8QvZDGeyZnVD7P7h
IyC1uFaTciTRc2jBdY7nzhF35EHGEplmfnRmGbDQFDVydTrKMP+uw2GY5MrwW+j/upluehV+pT4q
i4vSIWexyElZZob3jwV9s5ZX1l9s2YGiidy3qxr9EXa1zw+aC0wSd/Y08mYqH6N3w1E+Xe4Bwg1K
rxnwscj5IxIjlEH16kvT/K0mg0fWBsf2H4OM0aUiB+KYC0vS95BohVPDEME5txkPhREjK9GrhV4J
zM1RmxF4YjmpCBWJJvLoWAqtvn1zVyWq9P8awRAO+Tp9jJJJnTZ5pHpQDmin5pGn4X28idknxQO1
JZ2FEzl2VMfs4799DMgtXyPwvvdBuWBAbIZr17TiCrHLVPS7L87XQqNx4FgeiZT7d0BDDzKEV187
//RzvNBr+4U5krkYGp4nN+Gmt/ozwC8O87v6L6FtOrnzjRROcdY3p7S5RTH2vADqrxJKeDh2HDcu
NauZPMP/aJXqc1e93wZxvj61YvE3d8O3YEqK+FAUjRZcauh+2B11B12la3WladvXeqffS0UyRPOM
N3QEN2ZS3St4ev+fF7fqNewNNow/TlKmN1tqTqEPA4IlW2okE1s0Z/flLAKEmq0E27VR2k4R/FkQ
OeBpuKncyfgClRMk7gvNlz+afAsAxbNvKpeKR0cVte2tKbcUBS5zyn0iwQGljB280OaoB9cFE64D
5BR6JIBwI1GH6eozr9lKlvOPt8f5d6aA0R7DGS9Lg/LY4qQeKR9QX/btrTCmAPxSDm/zTzumugCZ
/a5OPWIPufSLpxn/C3Ltg4MjqCvIXgF97vUKJLFOapeSStt2orgmEFEGlJxVM+MSmeOZ/nXG3IwW
ZbwCk96fv8gjdrKJq3B4kPkC2hRHzpbbVOswx6AKG9bLmNi0Qu+kHsg8sBniLhZpdpeLDBAXsG9Z
/K0hA5riO9vru0IcmkWzi1eL7ERZJTc6juA3GBMLXu6pePuDDa03RXet0sd157M+02YTgZIGFtby
ukRkvJFgoWleEfCLuxDjozQifbzJe+GebukXYEX8+jNwv3kLNu0yrXqOQJcj2nLHWBxnMLnBjc1/
49YS3qi9Gv4sn6A0xrUk5xzji/wDrld2QpVk86SUPi/7IySAkcMXfrRqHGU8T3Nkdl/XYonQpR0V
/xoCBbHIrxmBYs8shxHM+ZkXqqJafA22fWUCTqB8str4qNyL+PpzL0WglMXdTIedeW0eoXSWNFT3
Ku0vvZ9i8ts+5Eqslj8qpgqMe0ynVmyxgXdP1IPEGVBNWFPXc+3d9dv9mzdjLKK3U/Yjp2X8WHzU
5M9HLcXNWEoHG5+/ONvMD+deRtnz9ExpJoKPyIiaaYrepNbhuYLyauQNxQ0bFzIlXte7rr1AX9i6
0t8IAn3LWPQ6cuxaw8cIegcH9pC4xtMg+RX8LA3ovsZEPeF2zIaG0XtRolqDIVaTNG4hzj4knaUe
r0ZqKQfvkAq2cVpWlQkdE/Y7j+l+EjyxwKyxOIzxf7T5xpaB3nvrr9+MyMif75Hn7yr79kGzI6Kv
dv8YP2zGP7PQ3LS1P2M/6QjDTMFT3yoV44eYlCpolE5+omta5Ml0OzYEj9WwoQcEnYxMlJ9nv0FX
FOAM7xqfYp047BA0kA6aIECyZ/WwFR+Ksic+gTF8WNU+VoLFez4w/bAR0yH/oZTD1C5vHhsSQ6mr
NtK0KeptizTuIbG2MWbG22URPH7juaeq2k/ttadyUn+V/KrUkFtw2ILt3qvesTTSL/sP2AYeXxnH
lpTooP1Tr9AND4hLJn6367mOb0IfkAHf/h9vlqCpZm/V8tNPcXBPjNdiBLy5Ov6g6BhYJ5K4VHh1
Zty60+CY0orNErmc9YWpptofBGQ9Qj0VosIHd/EIqgbGyO7d20u+RYAIoaNPfPDnqFsiMVj1v1TT
CPSHyUZG1sy4MxukUZ4qkUsiS06FwAvcLnj7DRLSxOASZi0q1qX1JrteIwQ50IojVQdseW4qhFxc
mX+i5SEU1/ljffC9I72g3L+aiLPh5Gc2MoRggJCYiESHpE+ss+h+9elzLnGjHORHKoLd/nw3nRcG
UOhqzVf9zPwuFv2sj2ZmBZcDzvXA2Lpd0G7twed7ISVqFv0lbb6jayhXfk22it4yy9thou89eHb5
qR3soWPuGQ+ryeXgAvB0YQChNbGw+UomD3t4LwEdfQVa5NYL+EYvwNqAYYGBErxIWusMPBDwgcYW
Hlsv8vK1B8/uc2ClyOzGTgNh7/DXMVrbyXZY07axtUtNca5TWGhnPH/rm/XGznk7ijrxbsntylsG
seS2ZSk01r+tXMhORthVaoN3upfTqQk1Mdj4NNHl6EQAP0iTkfdR+qWmbbKQ3F7aP+VvmDxQB8WS
P6K5Q12i186tUzMjzkdbyHhrgwjl1Gom9hTeX4Pbkv73maQU+4SOrL0MNWEn7sNeYj2P7BdPDLCT
jtXqFXydzhropUnO9Jp3M7+3GRwRmU/qGezDF7BtNc4Ivvzjs/Av8/q0fpOw4O3sJlTKFJ5c9j0s
uK0962C9dx3n9Dy97R0zNkRLzYgwlOP8poiRTXbISu4CzENaza7rckqO219cpufWNMl764cAB/N4
UCHEjYv94s8YFhUA0oo63cS3bPp9V3O7w7FKvSEeTE3SZTOH/bNJzcgZ0L3tyW/5rJc5jOPVqUvo
1NGTaGKGR7+ZgO+hH6fHqgehhQXsQLlSlA/N/AmOv9tbAOOqlValdim0uXfJZjkCGkbkY9DXJqI/
0+ZgC5vokIfKY3an5C+/BKogVaoLl7oC9yBaf8uTJm1jaf4zq1O6u9xjoXIpqsJAyLUE2YTsAX6H
SPHesoNxgPZKHFvf8hJQntHWZbRw4q+tCgJy3Mgw3ZTOSwA41zK5LiY8pSwDWP4pz/N4QbysvAip
YExyoS3fnX2/ynCd2NttguD4PRt8gh2buTHf//mqx4zc4Sw/sATyv5qJO6B3Jana3cooOyrepxzC
d75qWRsxgxNehS/MYJMYxEynw3jGTS3pmhRBYtgJpitBgbbCFxrumf/Rq9hB2IDKKs1iIY5aj1jz
dlfvPHGkTMPyFNoGgyXOULvII/tfdnFsAfoP5DkgnC0BZJ0xsLF2JoYpPDwuPTvQkQXH5S7A4FWH
OA/2kunDNh9g/Hnmjp1rc8C2kKalntiM/aYv4VKi06v718bufnUsEuzDhVD7je9vCn9bGpcasMt6
3PfvrR0wqsBAx1/ttOXX7o/J4zcaVrU1dBXQgfwgkZQ1+eL26vcyx+1r6gqax3tshU5tgzuAW7AB
N//fQd4udJeEV3fDHeyenZbcRic5aF1WYo+TPZ5o4U1zLyWQ7uX11ybXsQce7Ow5CWU57l+Rn/G+
Rjr4Sredc3MSuHXzNuqozGHk15zDml+ucdR21yN0V6Vig5IJcURRaAVJinqbQ6t6K6kHF3yTAO6D
SUDzTR+ByKXYme9XGm+OEZ+hjXVGf1Ftvy7mcn83HETtHHfJDEJGGFc+0m8+m+LIaNoHTDxc9awv
Q07GZoRSmaaWSQc4XfPGzw6j/5mmfeWAMpqimmrVErDf6/fhF8R1vxEQsvlUNoQ3qotOGsMOtbmV
LqzIXgkunYDV1ZEoxYN5/pse11RLZPOtE7dCYFmYMqSaIIHp3SPt8XfOa87ugjeT4E+MlaXQ7Wpd
padtfZjG2oKoKRGEVnonsWDVzecw2YI/ezhFU5BDcvXIv9lFBt22lvploOUvPPn9bLEdzxbzJrnQ
JyIhx/oKbqmxWX0ck7DpP42xZdkrr4KGq2FhNaLSNXmgTLDVeoZg2zxc/kzlz3ACRU2mLALs2pv4
SEFUURTX434Q0D3SSc8MOU3no2Yt6asUUHplKZybm9cYNGZda/tWqTtvxOnmK4+d0Zcc6gVxUugX
3tbOX1WrBsL0VeCkkrnCO3W9IlV/GCYSRyMm7hHg7WFzzawlDh6EdwPSfmBrvflqZxHU8KRlLj/F
Jk3gHkd95jx+vEGJvMbsCy2FpWDrPQhBdudzWYcjqwQnagAskQeOnBhSoVLZNxtoDgKrqsKocy5z
4WNjX8YTJW5g5moF9V+hhz4nD7m7LApOA3nYjcr+dQpDjYs5pDv9qL0hA+JA1iNfo+Xvk5h5AT9v
sjnjZUZWB8WSju0Y9xBnjGEpFnbZhGIHuhoMkHcGy7zt+FPtfJb8yTdNCdEXpMC+yZRWfs54Ykwp
s4DHPKazuQ+RBWuf8uHj3zHiKskPLpto6e+wzN6ZCVwvrOQR6H8dH2Of99SuFDKd2waIa9HSSaIn
+GSOKt3gvEOP7xqURv5PJVe/9WcMRInYC5ELDhXaTjAphrtLNMOBUm2k8VhqI6ubLqqXoHJiFCIE
AvMoGqok1adgsgCAuoVNMeJUHLm2Bjw8YArH+SMe2Kfs9srBeTLXGapEOjZPvvBMKT/fcL2Pg1Ba
fcaf5p1dtrTu+UrTPmBy53lvYa7GFs2+fIRZ/xZGpgr9OAB7e91TUgD3XDnXwYvdEEYZfNYEFUIp
3+Iz1o29hzqBz9TyoaUoplszEAmWNKxSeAkFmjqr1gQ9FkVzfHlFTIx7aKDo45jCKnh8Obm7evMV
FCzOsAu3mxovtGRoduHLOEg4Bo2AhNqW8WtNKxfDzj1jVPECnBqJ0zCaQJSVUVKMwsGEJvkxrJRQ
XKBk7Jmm2aY7pCcmDQ9DmnwNYb2+MnCHKindoTzVfoDVBuJzKKdoA+xag8lb5LfDh9ak1mE1jhck
DvOb0H8PeZlUzCRtuZUovQgu1wu169k3x9kdPtdrCUeVMFZmOvlR6LI3Sy6QOTNPITONog7Zc6GN
eVR8LFYt6CopDxS73hLGnMo5QIUgFrIaHjsgzme+zm6lxY9EYPababzHoqg+f9U+yOuGvv1c8i/U
1OfZsZQnEzhNGVYUtU7uB4KgFltnTlG8WoyFwYLEegWnVhySvJCpX0CutTUQ36bc/6DfFvm+rBnJ
Iq35RKFDmdeUsXvsZ4biT3AtAwTW/SLRSLIKU+qVhZK0W48nqknDwzdUuSVVRSlgZHwiCyvKKzV8
vZ5m5VuNBOC+8V3HqiFdCt8BhXKUU6DlD2z13DU4y+Bg6nYRz9S615jqnKqe4ngo4zd3CHKBmFH1
PrY/HzPqumYmiizrcTV/2o+UcrNT9nSI1pwrGepbzGPXm5llgYkS0D88i63IsGZqfE613cNk5L5V
8D9DsINyOaW0DMbtEyihgoWLYL120K90DVcSHBYmc01uVC59PfRPS8QNA7MBxx0XN1vlj+fsRAFq
AbGlSiC/js/2brBkQ8hDf4MnGfuYElcfhdkrF7ORPgZ0DNDmWc7Gw0M8I7qP2UhejZRWr0uOQjHM
/tOz4HRtNQFCz6HsRoYxqUzX4RE7BFQ+JR9HPQrP8boequGCRZ+Nc7xr6cDwg1i1ATdT5m9s6Dmo
n2gnS6XLeBXYZ8M8RE6pLWnpHuFzArIE+E+X/YQTUXmKIoML0F8Qv2OOiUsma+xzkyBo1UTO8OFB
kqpe18MaTb41+uYwkUqW2Sr8U0UNLdJJXHJPjOB9Y3AOsX4YtEQbd8ruJ43fD4PzkRfYLE8G/oov
ZcxJZDPBtJV5DeRWAcdv5EWRsz8tyOZiEGosOrq0fXyI1XCcmQirb35BvRvVsL2w43OIy9+Z9Ssz
qSs1YJP4PsfdvqZ0jKTxDpYjCNSIQZ+SVaSRWgnBE+8BwPOj0hFwP9ztMn9chn5iADMo6FHb5GuS
GVpvaOOcnc/ZHyLTc5eAQeMvbUv2Y4GOyxIh/w7C537J20hWB/567gXdangr6SiAcWLM2caeFK4f
u5AdvUYDbXbPFy9YAseXMIWAA+qA+r6RJVYVSXw8wdq4c4HGCOynVxCrXl7yFGinw1X3XJS49DSX
Ip0aoad8A9Z5wmWGSoFaUZfN2S9//10qwF20lNGfhpuvhen9SFjU1gaEVihOA7rtGrg2mREro8w7
pbI42iCsesfVuvC0W+3GCFfJBE6ID9LQXldYGqL1FPyzKRjKGQQaCWQIWoKPx4VnSacGvTpSIZvV
884Z4Ia2c23BiTWIEG92RwvUpAwsriwRQpiF7neGEy2Mpf7u4YILKUGvcnv4dPFPN7LF8NFvPdq4
GDq+tNWs+apd5yHbIGe4wDQyYMh5gOqiYyX+H6Sqtnh83ZJ+mFelBVwSz4NkzZ+5Oi2Dfs45YYMl
UDA59umu5uqCEiNv7G0L0iMEURuymh7Ga6wKgsFpY1iR4Tc8l4z8WAeMnTCrUtNlI21VSXRwtdAb
m13BrVdHgizzIowpvFsCAY/r65GXQ1EY4FGFDG7MLPbT1sAUqRqpazh/urCTJrExCne9QgRD06HS
YsQurdp/8VRq2InKBqlGPRlQ7zDfgpGZCLqndiebkZC8gfZvkKFlF8oD4hgifn39Ryc+Lt4b0E4V
90xLz/YHs2c7Jb0R+pSh811YA82yDSd+/c7yct8UxXshS4bIUr4/z3KtsX7BflbRZofZ2k/skj1M
rOR3NYTVCVVGDIAE4cxOSh9685UGN1TxOfJ2Gd92fmpvYGTXDnD5rkvbxSq7Kt70cvtW/H06ZSLZ
OZ8ZS/hDYM/hXIDg6iwtBw3Jxzvvz+ZqR1PsRiNI6OPYduomDB+kKQ1iMOfpuxf5paftHJ1tG3Wi
ao7deQM53I/irI9JOLPIePlW1OBhdogspZNR8XTYdPmxTr44YXar8WJ2bcCHG9hnoranX7XT+VZm
RbdXxrgbkiRp0sroCPfuenPKuPGyErEsxmQfmh6QeqxH6cVxC7rYlqh8b9T+iSpo1sY523jeOqUG
cwuEksJ9b8flHUnW+vivWzYJgXzQS7IV2UVNxLbgY+nubjSSIqN3zcyMKvntXqRewvbyGQzFsMYZ
yLM2CU+iN2p+A71SwoLJBn6NaaCR1JZZaDxDSijxt3RkALlU6aexRxnLg4otS9iZIyIzj8oqU0rm
g22l9BW2RpR+V1i03KY5BDjHMczh/wtuwWjKeiRfoNhz5/XMbL5XQxK2xkuBrev56MQXkiC71CJS
3qUIHo1RhnM1gyQyTRwgNNKGM+h6qZ/15gxpn6oRzFowm/NGyMJxrB6gVtQDNZ8N3SSGmOnCV3qV
VHnzHwiB7POmuaa82DRYaKurAhIjbZuVi1chsQJcUhfGk9CfdhWk6Dmr3kYV4CLaLUXNBJVzHYls
WEV2IQZrPdgawrZyRrjOd+y1Cq0IZfVZ6WOfvMY3oKart8kLd3jxjuxa32tvFx4Oc4wSSun/JVsS
pLA2IkPLPEXXEhihKIiJ0uQYxGMJmYZP3SnXLCDpGCLhpjcDj0c/Qp4zY9vgYiQMUD8Pi4AJckeP
j1GDSnMvZA4u4WWvLnPfTa+DYPYJStzCM7HhwtTec7HyjbhejoSDFXS1XXTbjy7ZOPpBbz1xXctQ
e3MEBwtfvKxs57pAcylAGsUy9zgJELrobmlTa+ic1Tq1dyRrWK/veTqmxl7z4j0Hj2pqI8K/1PEL
hdOGkyX3UhIiQzFml3kvth7Zvhcj25kfeuextT8qCVuSptBJ9+Lq7uSNw5vvjp9+yhfM5+WQ90tT
Bh+e6lURbx3MzjdecSBk376xo5XkWS65rKtXIF3ZYa1xrSdFcrMF1rGKk/qledWr5y3cgVGpln8q
lCVC7RKl9MkXxXamyPH+IISxl7krOxtF+CJWtJdysgO2wstRh6rPQMJEE/ddHDT24jhqeCpHzYyA
NWJEDwG/5rACwLlKDpBuMGxH57mkZgRNDpKr3wEO8aFUZP7iofXBrAbVJeplFmzz1edG6FB6qsbX
hm5FFLTwHe6uA270+FGkX2GlfROdiKL9Z9N02+FoA4hF0CGyPgs3KrUeTbucgZ5Ubon/DZI4Upus
2/c9J19j6h4ypb97F23qYQN/OeMS1d63X+BI0Qn8kjgaKuDp5DgeNLu4/fYOrXjMW4xDSnxM0f2h
M9lG+14s/mgCKsEtweI9lt6ysFMI1XEUmktMbUMfmby9g3kaairHxeYA+LERVwuzl3Qvbs02HMUg
ZR/txk/MBbs7APDkJk2p9soOLOS4EfWmYav4R2YhE9OD/sEkckQ1yEZThf3V9gLGPLH2LmmjlPbL
o9lzu5eu2l18wpZfGeA/G52ZTJUeWpeLrtEihPxR5u50LllfVuhkVPCFSCIZzb6KgSJHg6tCz0aV
mxazIWpwYjzeAXMmG9WFzpmaBS9p/d0lVqfcXOYCQx0iAT9/pa1/guzlFf+VDvPAg98beCf4UYep
99bQrJzqlF16MtNCTyZMZ251+0jBLB37RcrzhQJ7T7SYk0Ryo/TLqyVs5FZboc1ZZOrvoi75NeLH
AA+SaKDFDO8K9iriBEDe6vTxoWkFXIM+1hpIWzCq+pRkBjn8lFEn/ARZiKjiMTEKSf73goEQcHcE
WOWdVd+sJzfLwUqBF47rVvMNHOT+hnPP2ETS8rd+oH8tvvX1NHU7G9oWZ9sco2qFyP1OLoorsftX
EuQZWlikSTOqnB475XeSfrQSnC4rYujH3d16i/r6z2a2i6iRQqIGLGURl6PTVQiaJzERYNjv2Hjm
hxXQE2UIlZrEyhuIFVOXtmSdp08WTGRgjkstd0X7IpvLhxPbDQKjNGWfawO9We0YTW71Vn8rjeqI
io56YQ1Okp81I+WIXSxnxPhBd9JUDjK0d6DG1qefKT3p+sFEBy1/MVby3f/vEq5LPBY7inB6ICVC
0gn3bLtsfX2R3Pz2YYUGOVdKPCAVsskEQLci2sBBHe0jiQoDN9KSixnYJxlXoVLu8VwLu9B9+p3n
fqerBellK4SbvPFTLfNp4RFWbGxwlOwD1B1jcjH3a9+fMnxJ3w0abI5S+VlvlL9lxTh0eg3L6DA4
HPrj5ntBXxphM6GVMbUSH2Ll7Oda62eqTgYIPeH3B1Gvp455VSCbhAeiGay5r+wKceyDstpAMoI/
59+KvEIFrRr6Y3yNncl4JwuMSe22IyI03Qz/LgT1oS1Zzu95tq4JoT8lU9y2z8/f0Fcnbe5JKvJf
CC8jAFmjXEtKSeqevxUetGnIHPZ07toZe6Nsn8wJKy5rQD2zjVN+vxv7aq5gzmkZLlS62sTkPXjh
GwWNbr9Y5/msG2kae+3NdNr3EKS0EJR9P2WclGUO5z/gYSRHlMxDqIH319D7c7qHE79Xk4N1gGh9
DhNVX2a9Rp0JbCWNeMZ3Js4bS/V6sUd9WBMH4wb1/7Xxs5Of094BtIr6EmnB278gMHNT+orIlYD3
WX5UGHrfIaZFF9PxgxN8gkq9hxjwibdTiG3qeHVP0Cd9Vu4YDPx9XNcLrL81iAhvhOhVjTfbtfW0
cB4XwHFUQyC1pGA6+04t2/SeNgGxLhPffNOaZdeJtrvrQg9w8qqkLVbeux1Khftk1x2qjgUz1MDf
/vfD2AfCQ45u5YTrBal2CD/aelFxg4QrHBG9O0l40B/VbYEIN37aSoF0MS5AQEuolHDg507ju0jW
9rqFpXiToWfHNloXcwuZb7mnXWoxNLHriYbO/GSsGaAGmDM/iUyTsz2O9/NNktx8ZyVYMlNzivyS
EbxI+6jhrnY76QARJlnwSE0ecaL6oA/ZNzOjWUhL66qZIgSija/o4KPXKhWAI6RhowrzNbM1pr75
+D13XyjGH7FofkONdt2PPU3jHmkI/oOgxyVRpTDln9SPHrr+vWr1omMV5Cv6oUqsD2viGQlB0mTh
JGFfks1ChwmNTmU9JlLVBJjcmEIxfNsR5M+JmbZdBlrkw1Olr2GIX0SIrWZmVNSBXTbTGknGi/YQ
KTpdrVBViqHZ+Cx4z2Oq5WjMwH39AKA98XiDwpQf8HEXCi5bI4NCUs0AKxyhgP9w+Q7dmi39O0XC
g3xOH1VJVHyny8dvJKrD9ZpEuErmK3Fm6gHB4bv3Etntujp0U0m6i7lRNeXVF6mFFnGfx7tDl/Bn
MUq2E826kQU4GA7Z/roC64E3LX8t5LJ7/hAhugNSTaFp7wl93d/Zimipu+GTxF+Jp6ODB4pCniyD
Wxg9t+MN6hxZVRU5CYYqtVJwdqw8Ey0CuUeMoyE/mIgQ8lXBTZiscaRBd96XDhp3Vj0IYpK15qew
WAZuCB+q2sZymwP357x6CGl14NjsWouxHMFsA174mQF7EPWWlbhBnX5GfdyMKqpWxz4GUntG3iav
rewuChmjUVFerw3HsOrWNzSrDvOZJpMuxjQu3gywD8pkt6lLDka1L7O5pwNzQxlXZfclqp5Jn329
2dlmLL/KX1YZZ68U42o7H5a6c9uC65EtoeYHKbkpOSdIaAmuOvM0qYf+Df1M2wDGnEu/gD3IZsB6
lcXpnyFhB1DNbKGEGnaN2l2rNHPJSHYC3yHgAyErLnwSKqteG0i6p4QmgXfnVMP5MXnHWGc5o6t6
/rpIbB7CLM6fV+j+R+kZJsDK/9pptBPTAUHaMe5CQF3qvF6To0c7W9+hnft0NpDbZd3iVSxNJTY3
0+9VhkIJsDfNF6DkJEjozQGyzCp/KZ+gA5OiktuslcZ9tm2ClEvWV3YUrZ7BaeuTMEZzL8yH13JT
BiNbMQjDQd5pp4ZQkJkZH3bHtwFzGMYdbXRlSstfTJpUFFsH6MZe3zOH3R/m4v6O/Hi3+7O9ninG
z7GqnkdmMCM1IBUHSw8UsQdkxJRLTYUx0Cm7R+6YFwacnOxpd88nDX4pt1iPo4d29I2pKNlwzBZN
I0sC79eFUkCMh/qpmQ1alaadaWryhaHCUobhio1H43DCaM9q9HQ0VCFYlUBqSerwo73veY6m2cKY
+pV63aiLtKcFE9YGncoBJols1AVv76k+wkm8b2MKMPaALRHP0SxNiXUXfYKA4kpKiY/HwKRA+IXw
qNK9UXL0lp+Qccq/jmCiL50FdhaQVyS94zJBbeQPaUK6cnY/lx9rUhKZMXN9YopEe3EfU4AcXuVP
X3ZKBdBQkdcmo66tDDOVesfFxYDc6UqIwPLdcOwRliJt7mwpT5wGEhB9AVc5QHjs+2gVie8+BOHo
YNcSvUsXSiDWmKm+GmzHmjKYHRka4vtxMft6ANIz14VmXSh73mao3YDpNhbq9WumkX9poD2FKC2P
1W7Pwg+2Bsw9/TZTdTDMscBbWKIZJ3WOR6c9YRrsdfKuqHSra13UZpOtgTFbMciN4ZOakJGjVRGf
BlBx+S7kdYrQuBku+79l/Oh5IzcVX05nX9e/Kjw+I5ZMjzrInEQkovuVEUnZH7DOLgIhJ8n5vONE
sXn5IDhlr6aOjZnbxCnnXJIvJc0kG8gun5MVDLKU3gp6SoW/VADk9QfY0UxbQOqqFqd/ulpx5h9/
AvsfeSJnkHYc0j3TCFMNMpzBkGrVCQ4YHaJWPYBxYu9ucRN+83iVmjkzyXNx92vgvxTiS/aaz5CO
1WimGQLo3eCjv++AZSHaCQxMmT8/o5xkMUubLgixU5mgmbf9kjV83ysPN/LA5wB/z+xtjxwbx1oW
C0BG2PiXIghB14n/WJXySpnWP6KQXneFG75lXGblvOFmxDZz7FRlfA+sTsNXwkcQdyJ6DZTrH3eO
fzhMgN0eog1xOy20BHdDwlMi7KOJu8/HrjqHwguOA4eQotGe55snVWZP4RFhyZWTiXgLPm64cDjC
BYr6uZja9sHXxNRCtUVwVFGHSL7NPtQstvJZ2cWVDOP76Pyg0ZVHZTafvp7cujnoInLUYnxUbHhT
H1plXb1GzaULbTjSiP/MSEdWRxV8axMxMuMqkCCCgCrYkzL97csOw4fu1giA0lUJDVpem5Dvnd87
mD5137Wm8lUpR1Rj5QR9E207Ty50rd8NbaY6gE9Lu5PuFf7TyyFW4RHtejdYEL4oKikLY25HNd+N
emBxx8AUZT7O4ywEVbeflUlpJn5mpeY5BqFRizCxbcLzt7VpIiP8ytTDLvMkbWGqvy7k2OUpVIOT
vqASjDxjRDDUj2neVHpzxPOCDxl/ooSwiIT7UeewGHddm/44jpbImNULnlRyWy5n9wttyhMKJMnV
CEuCdyCxM/8ZedaShqAR7sGLwAdXk1D9UQzxBN8oYdo2tF2eUDD/65QAl5PeDx92yfXcXjMOz9Mo
zdKW0fgimTtpKHoXyjXlorPCJEvP7zu5Vyhi2UkH7Wxo22JKa0UPipbJcUvXO1B3V/qfVKD+MpmC
y+1RULlLbwcqLvfRj8Ai3fXbiHwSD3ps55c54Ft9p0qqjY4boiwk8C0BljMgvgsuHdLPKOBdeZa2
7lz910XdPzSoBQZdg/XQpT56Eqnr+cSiyky1b5YkV8Yk+HdllyPfaTZGBtMIeITqSUCis5kY0P8m
I95TrE/AY63DoP+3KjBsqg+unX72PKSA+JDZgKb1k5zObtjs2+ZlflndBQ8UJO9GURFlpL7tk9hD
8Hu6RgFuWuAnGLJC/SSLDDHgppef0XN41nJf+fIvhw8MDlbv8fZ31kpotQI+gheWJHRTrfO5gaMM
HvpOkk6lJ6KUizxoBbgwRxvi7kgjyo2cjL7uJYEm4epgjyHO8TC/DzqJDQlU7/FbfCErRT7j9lRt
Uyxe8NRMuT+zUp/KIrfTSr9e27DlOkUhZg3klO/Q29PDtYGug9Tz8/8hSXuSkFgDmj006jeAmdb+
qXzcpVY9PGLAFQ97xnu+P5otCe9xfe0m6IqGBn6WVpEq6kpXLoESqCKX3r0lXFNajvDTOISfVos9
mc6mH9dgy8alZrahBZMvRJFCw4m5NDvTpdC6yVlGQ53moIqzdhbQHsicN3DMUNL2kEK9274T9SvC
IlSLNbxA8HeCqpgATcBXN2PeggTYP9PO7ZIFA9S0tV3v5kgtoYbcquRJvAOKyXQVly+6svO1lY+o
Ca11DcMnB19oGbTDy4ksFYbdHejn6+9uKkh5lNYy9lYROtdx1+wFk7lNv+eiGHBawrltuxC6UaaC
7WVsAH1aQCDXqYjBwvxSzA7k1s+4iqtf+6MK+4B1DosL2IemF1C0e3At838roC9xA3flVqDw9DA3
PTFPbZNghpOFObdf5G+x4iALofiPAtJ1O1z/vEAN9cYK0a/hv5E3XJgXzWdApAzzuhuy3ZKhJ1r7
qDFGBWRXy8wQsVSUlazYlurZNRCw3qGiAT/846wIvvLpoWLKhj1xcU/aqTyjqvnocXX+RS8j25Ie
IQ4iNY1hBvVfbflSORXgrtwfBLil89lCV3rUy5ICcrdqJt8rDLJzWpf3iL33lCvGaiKd1N8snGQn
p4/3sOFmNpsli779oke3gTocsQy4uCq1Zxpt9pDUeTRsFgilMP38aVunxOHedY/rCb3Aa+q06x8U
ES0hk1tTCwIbJ2a5Zvpe+zmNovBxO+cYcGR6fuZ58fLEaeEWEVeE1VD3wlAMIrqQEFqySkghvtWv
njdbl28WVy9HaKouyuaY5ArN8kn9pOnNXZIKntf6eYhVtRlgnBBh+0PEOafBGRcYJCL0Pzc/ui8R
pS7noiV3P5I67Ll+4zwhGrBeJx3WAhMqGShF4+cSACyMTjRxQ0U+3vMNXMVwYtpr0oIE37ryCgys
nZbZHnCcz4xHncR/0Qs26yOTCCRu0VSidET/oD1Coxzq1EWWJ7vJ1X7SrvLTsVhMynBA12l0zgW0
EUXTStaMrj8ZIRYt7RGIX8De8v+Q/pAEfVanV6dpcvrwRoXB2QaWeY933McsHhltMv3xfZkkGfqx
8xqUGB531Zh+Tcvlhe2VdeWEgrCt7z0fQmi05TZP+i4xAeks9GyMq7ISM1X6rwHIEH0aJDGEOjvt
XRKlVL1BDStK8T1nb+6cNBqsOIUw6qOvft/n8QlGJWFK9z1Zk/Zw2e0rKPIzCI54vCT/CcdryIFN
sUZUdcEbNpySvXNWRFKYrK+tiaaxhdEqPCSHDeYwNG1SrhUpOAJojvfJN7I0bVvuliEaTRp6IOio
vvpXKyBY0VL3xZn95vwaidot2OvQ9jC2dL5IzruuOBrEzNK9ul+XxASNC1+q24Bm3GzHpYdYNqc4
ChF5rjqdn1yDR4Ck1SATT5FJpRz4XPdqHdqA9nUg6f/KEAlHHyV9JG4RE2SheF+zBxho/XCwviw4
OqkRH3x5ARRnIFWsFqMB4mI3YTEo1nxIdlrH42O8XgTX9UlnX6R//coi9ivuTooChs4kqZTqPMoI
QdZ085RUDWV0LBxOBhJdi8WQfRMTZ6M3NuGxMeEYD1dygbcBx/ItPoXhNyXLA2N+9PnDI9J0/2gZ
KJDKkp53ZZ6kKykqTTUA13xvCz2zJ70ShLihd70dAW6lePwPhXVswtmFBWTlIFyRzHgTGNK+VR3R
YScEGRj8il53qrURrMyyFis57WAUDwQA2gRXrFH2atEJXsyfnjdeB1w8wbMb+h1AhpcxfjIV85KQ
BYOyxvkXGdofs/0IS5AMR+y8wjQ2O9BJYmbdbxBkQk8nXes3UrT7cdPv4zNAKIhOn4b1KToR5Xil
h92dwthMa3Kw5A4p481Hqh09C1IEnDK7tUU+14jc1gx0Stjk8iv+/pqINUNzrQ4j/SFlYPP2vo3j
g5JA8lY5HSVoZx9BzR7oli/sZgjASaMx+v1Q8DB3SnxsNcoWJNNK5U9ChnGNrucDAsuuXvxHXgh2
kNcMHVI/bjg3mjWaP3HVChVpwn06bNn8goC/S+sqGOgYD0T2+DwqSdfKgda/tb4zY6N1ZsCVQ0F+
sYv+o6v/MnkdgoX41uT5V4DNr/VBktzcfg4Je4lmZUGoM0G72dVfeIdEje/Ms7M1KRdkA71zJsLb
Z+p9JSTFgMfUdirm6aC6sSlMiKP1fxSZaAcTZHgOeAUkNCbeMNQelpLEHSb4+Xzig1JG4J6LweHx
ECPw+luSta+ENCWw8HGx+FiajCGCzsWfovzj8nO0BQazhF+vGN8DfjaG1HlzRjkTsDKAX3vQa2qn
QkeCfb3ELYUyyYBAEtAG/msdhGoXxAExS7z0hV50qpXEJgPZ8fn1nZOT/r2zGWRnjLCphh67GBhJ
S0M5jPTsIDChkpWpavB8YQIXLucWgm75b8nb5AKvEcJMdgY1DUoED7EHj4717hFDzvmSR5UEXrCN
b5FapqObC+tgCyUKG5V7VotVBMjoa36h5TZmQKoXdCtpJnT4hzzHvKZMrQz6mkLPo2Eoz4JO3yRm
Y1nOm37yymarb07U2Hn438xgOH328CQxq9USWT39C37X/y2YyQfSSpy5e4f64rr5o57CTaxKvAIt
vb6Pe/t9TDwE/tYTaUQ8UZx7rvIpde/NvK3wUNyLfbbKRjjO/13jz54K30RlKxOv9iVDyFL8DBDt
nEjQPgnISAgu7gfaDEzY+Imvj0arbxp1rgHY7Vy07aLwi5KGcvEm1qqMlLTfHwoQni6oZjGNj3pg
HlWi2ycudj7wbIHpCRzN2jYWRDFhUttGikson2XhiulLd+0RwA2kQEZy6IfgpuyNCkW75gpTHWva
LgPou8G1B5/t5skzcVvZ6RMwEnI/GfmP6FF5asofN3xRrRbuYscO1XrzRx1Bx1u0RYhrkf03LyMx
CMcNcgFhulfAjP+DfVFtcR2ndYnbKycTGuXSxARXlVHnVmbToeXF6sWisVPW0LqHpQ5o2Fi9LywC
tO9AMcM0pCql4/quiszqB982251UgY5fZZLy1wsD7g6oFAme5dbZbEqM3bx+m3inzu2i3pn5kenV
xP6Z6dPZCo85LS0NnMQ1wnNKe83sQdAC2ZJhTBMai0X8I1y+YF3mliOflRDFOLVRKaO5NCqYOo+o
dgUVbDpVzd9/hsZSqsGTtXrT4yAy3uP9SwNIoGHLKAMa4OATq0WbQbE4JZoB5HkklsgQYAxLJe4s
k72Fy+xncQes4giQT/hrW9+LL6fq1o2IWeq+AcqCWr9LdEdkXGhywAD9lHus2GdKDqO/Bh408SF9
ZERO/YS5lmSI2ltWcbNulnkcQ9sdV0T9EqAs6J7j0T8IzQRiJy3VRsBcJZDgyhZFEYhJduBuG7Dv
zb8TdcfDDwNW5uFeUd4vqlg/XUG2EneaBmPxBowhMBkLNmEZzOTDZ0jeR0nJGC5Wvw4+LJ931QVa
W70POu8zLWWzYVGwVpAJRYRtSCBZ5F87/dlc93J0UfVU2Vt4xoIPnNp4KY5wxQB2dYFslxHZbOEz
hD1uEGZ1otnBumEx9FdI2G8JS3+mL1hSYf9GTDsslLZNco1ubMl3CjqQ+myhI9KLT2dvYwcqOJDj
QXRX+iHRKFVcaPdNrqYPsxNRpVgn50pr6TB9YAzMQ++57+KFAkBnwls6p1DD6fVOnal8UXhobCON
qPmAtqJinV66KWbLIFLBC/3S+ODZWBBp34MSRuEkM73+TA+0to/ZEDezLXrUH+sWRxZiH2Vx6qlz
nOCMMMRhShJdit5Hz/CzOmDieHEUBqcch+PnyLb4BSUOWnMNt/8LXOPLfWOdJPG1HJGeNopYQFJx
sRntvSumXXkITmO+FNVyV9masmLmINL0K/PIypAkdVac0X/PCCiMQuAIjYb0HrjZAwWBQxNHaUq2
yxCJoOxOtOwnrvcc5Z6lkDdB5VhTJKL6Ht/ke/iixINO/+MeeI5Q6V9H9gkVlaTIMy058e98dlLt
v0Kvhzj9iq4N3whZvskKmzw+fWvkl+SvbFVau0oPSzu/dalC+P0IGSZrb7d0YOFdbhLtTNucx5Po
CCdDF8qXbZT4AEsDln/pcZCrNgIT67JKbx90vE1YcubRTXQe1ozFtT9mEg16GKETz1pa6FxKSnYP
3VnBdfA7yQAcjQu+TlxZ3oc//srUGtxQeMk3IVvknCjkrvLEc98HZC/wXkZrOXtUyLromqLBwMGz
oAg1oG5C7/BUcjfqjmKIEHlQ5bA7B/mHvdf4bnV5VKTaXHoJHK/pHD3y8OKyga/84gmgCOGOvgv9
IhYTYzpCqeIFOT85H/s+9aTLGYnmodqW1+QcvV0ixiA/1FjTn8ZX7u2QjSBHuPWhgPTFLhNWKSdL
z0YMmfebYqKghi+iTvhWlFgdNypH/0QI28nBlAwpl96goNavLQAymEp/EbrwP5tc8jsPh1qpuQ1U
LQFLcX0D68+i0NZh1wkfecijyMrH43eEC1GJ09+6iwM0+c1nNHp/CB/exFOhMeF5Bp/kECfcn8Ca
4fO2ehSJ4keXhI5LP4k7PG8PXa3cB0DmMzzPex8/Nd3d8cfTPFtMK/yPyyJBSYf3eGo1iNf4RzAx
pTB01Ys3kk6Jw61So07bENtll8d1guXMIavV5PHRTvp9vspZWAGAzypN0m34gP5P79G9d/oy761W
W0PeLqofV94dpPvYPNJmw/eJz9jnWkonlEOBQaxiH2eReAlBnK9s3k6col0iVEpFRudGEN918tf3
3BK3c6MN1z5B0hLZsRvNyqBqoe7ehj6TMsmA+lzWZOcFWUbavnwO57wdUmPPL3/ldsA7TMeqLkb8
jxcM1RMS89DH15BI3a4LF0pQe7aoF0T9x96Jo4Du6QeAkq5srGTlPW4+O0byVmhmbjcFBL1hhsh0
YaNVJYsm0wdG2Gux7+ncxlDAnakbQjt81JOdWBNoh++lz4R4lv6jJ5am+c40MlvhLWDA732VMuSd
I1/WXZvG1H8be9N6TcjpQj7AusQq3OUYudq2TXHr84eMieD/3kCnOqM+ottn+EM7evIYas+Etdep
k1O1XKY6dtp5f4xv5NHRNKDRgCgMG0aAONYcGr05jwK4Jk6qPCJK3CN/dMnGysPyywk3xRSEFyjM
1ly925ldWAUm5zloRcvKl/1/c3k+9cqjfE1Tvj6kOU2dzRkE/FRjBQFg/1cdukb5biPBUakTYxD/
41KoiCFbFCf0FJz7U0OHTcyDzWP60yJrEqIv8S1RTbexdXMmgbeJdE5moCXXc3vpNAswjgjIag08
Wue60uxidMZ61sGXKzurD0BcVB1BHyHVkURvBPtZI2xTR9aePkKzkTOYFAWAX2BgeZjWvtUoYcCh
jfkUdktJNYJpZ897pWjgHPzwo2NWX67aq6uIbnAQhjm4Re6RJrK425cFtGuk5NcCDFXjpzRaGjSN
TTtJIlIdlbt6uMSRBCtX9ug4+4dDgLzYd6qX9Ga73B3CsDOw8a5KFOnQZ3o0i6RAn/3T0RsKXiI0
hdZGEph7B8QxonkAw6ZkTbT1QHvEoRaG+AUs862sNzbWszkYo9DvZv7Rmaguffu2hY0pw23SVnVN
V9cge+cwyEhfLhI66wN+PCOkCkBAsM7ZRLGoFz3H9MjeOfaIXOWSjWk09JwU7r3H3WiHITDj0DhQ
0n4IimrvPk0JUYWtue3iC04HzcpTiCxaGzjVF1zOHJwW7J3cnGdISXUBHuS/4Tq5gSJSwKZOZFoj
UAB/5/kIK7Di8OC5PjV4Z7lvJMSW8nZ4Nc3Jhouj392oSyxeL9GJt/kC6vXv+trXul99GvNdWBMo
rLdPt4D2PU1H8MSCd0wVAobh/8WOK/h41ai2QMrGIwL2v2iTuILBQN8N2PqGBu+U0bJE5+3D/Qar
bmdihPQWRa00FoeB8uw890c77ZF9Zwl7Q61HYPF/d/0AKWsrQ3k4LasAScrGw0LzcMNVltPbC0rS
sIoEeVBrRItb+mVIYyC7UcqqYNffvDU2qDmv8GEW9WEIbdh6u+uFNb89jnHhUhiDG9LO0SMAmRsc
LTgdb+/h/oz6ih7z9G9l9J9lYpXLxKS7DTP0ym0/38OEs5w5H+hIsEXCXkn7SQ6F2A9oggL338dq
S7lTI5oVtG7f8WKWk1TnlMh0wSztiw/zD+iYUABA/oxlRDzqhggYM8WC6xh9Rd4zrb1M/SJIKroo
vGikyeKp87eDxzVeGh1ziSvHmxlBVNB2EAJ95HMKphF0ViWLWGju/wCpN8W+Y9Y1VBR+jXNzLWxA
QK0wKui5UqHYso1UMfwHJlBvdNfDDXkxqNeeO1uiMS7cUjHM1p98eePf6g5CzWhkQ4JFMOW0qSHm
YJODkf2hH/52oxIelzCqjFZQWZrXWIeHyvgqu7kPoV5u3VS+4GFahCyt8welZnbR76l67hbVZYMb
VMjAfEuw8sdhf3v3CCfEG/3ixRt7NTDZwkHFPA7hRskRcdpOYZqbo0/Ty624WUEchXBa2Xsor4iX
aFBwwi5UwVrXNs73cz8jLoAYK/aUin0nC99wBMxa0p4vU9CmMDL4c7dURJb3khsYwCpTTX0qBOfA
69gJaTK62ZyCWm0IP28WgB3LYPvjHOnQPMmFYW+Zv483wkHmlN0TCIC6InppcdLfPJ1YgHILeBdE
fYo48Bwzgo6Za002DDOm89e3O8h1CeazsRVxci7QXuH1e+UWHN0Tx1NKqPXRjs+//H+V5f18r6fe
8k37IUmw23oXAYGEZ0dA/Q8o6GvFeVGca+0RdTHQz1GKd/FRuYor7eeAULTF1AfQGJjZm7eotO0o
Pjkyb5j5ZK6h7VwOEmOncYndc9UUBuzXeULK2AzZjM4ijLrhLxH6unG9mvaxI7+42h+l/PcZMoUg
2UZSMgPaTJBBkBxlHYbc5lmGceRZMjGVGM4rnwiqmEXNFhDwCbeA83U5xxaLopkVjUjXJ9AIxndi
5RQ4Kl8DVtwBRfozO1Z+DheYXqgrFbM98oJN0i8rHrZhnDrxZJzNwKXjY4xMJp5pHiHiGTslBahl
XGs3UAgngzQdbrv1dQ9z8o3qjdrKRHfvZb15AZCc9jv4Kr/evDFjGaL30S1VeQpVO18TfeE+8wZQ
zcuPlqChP7tUT2O8ssjBhcA4rQwTqVed+Sb9N5GV2GwWdU2sCc1SHNKaXevvhgZVggYOqBiB6bnw
+vcgUP1QBVZ8CXarmZxWZhOOt5vCODBG3eX/bQGa3yhJ+5zVuwgdezlbJHt9xE2vV7yIguIJbDlD
YsP4l9st9/Wy8zcl9Xx4GD8UFfpoDliUYz8F25XlhN3l6bd+EN63BAyvx1mTIoDJi9EjYEWcsEgg
UBegJ5qStEdhiqEL68YSJGUZynY4xf/W6oGVb05XIXFgZfBpqZNPHfbPlaEKSdI7o/QM95n8Cvk9
Q4gC0zKe5tetbpBX/mPMwaWJPesgUmuSqVO4Iwfde925trbu0IrhH4cUmC1UBdvFOThT1DvXEBe9
2UXTNEtaLdCwYbBqILV+JeNaXd9gncq8naPwOA32FbgWYGU6+265FNqd7TU2Rghwkf2nin2kf+T+
0UUG1W3otbjz8yK5ay0Y2rAJrA2B2wYErrwde/uin+uPegQOTxejT81q2lvWCt4ZfaBjh+V9DJQu
wNSoaJo2ymKCCHowTBNPMDUqxIwy0aIifICWf6y1KuEeQx4EPaJDZqOimUZVHP6s984MHlgwihKK
Q8SygyZT1ROR2S616jUSU7nasTPvzLTErH+Q6nxgBidmxMgtda+DZS5+yCbAiA7z/aft69ib8Zus
xGFvKnRC25Q0dAAbb0b/m8QmXOxPOOdej5GSo39TqDB6+zVdSoP7PtrY8Uy4HCzgwUpvfvp5F4hS
VcsPKV0sHWyD4yEGv9j8aWSDoBBAaBXRWMf4lrfFKWvR5On7xqYACejQfqNd6kyHy07ZaRHT87Xx
3kyhNkg5z8LtDNfNjjnfneHJ+lNV9i0OkX2nqRJTFPCR69sE2BO9d9mW4c2g5tJlrVpa7xq7o3G9
Bcmp+jiD/TyoTk4QdvriK6Tcu+8sRTHvCvUbwMcqDs1QhQv+hv3Dg9v940n4ZPMU6HVf/018J+l5
DcLkhk3OXiNths4Zgh3WTjnn1tBb9kSfGkDXf4bxhIyVX4DEVxyN9W0eGxAG9aiQSqcMii0zAJdN
N4QuZ+Z4EY8uLgRilLrC2qEmVlmVPmgqZ69qUyU55kjJ3lWTfqGdlVivML5hi83/R1TMQnRr7uzl
2PTuYMpky4XsYxZgtIu44dwaM+LRnZOJDvgBqYKJYivmsJ0je5Aa8ERduZBVfYHeEtNusRgy2Mm5
LFmBZkwC4jUphwQNL9NBXCWjitKVOyapU/JWcbPVuV/aWW3AqivRwdZutuAHQP8+166biH4nHHnf
ir4R8fap5yqauwzOtKm+etp1pfX810W1+WPOGK82bPeYuorNtEWdlJX5VH1iPzdgmoBDVp4H40pY
0qXBh9uORWMQe0FqMVeHoC34Vg+za32y7SiCAStzqinTyVIvyc8eE1zy/Efa8PEIXZE2cRs2QZA0
78Sn8cRSI4An9EN1JdhcQWqS2OsyJYFscu57RwXOP8AgIextwKuTAovtBZb2LLnrB7oAISsPl9Cq
6/i7HrQh6KYPX67CMIUsZR5wHFRh64Wqhb4+DKSvhEB6uw7wNw7TCaKAHBw7C2oxyyI4TeRi2Sc4
DjGOS5crlcG0XJ5uEPZhB8OWZHlveaFTVF8zbKkspedbLQPLGFTgm8cfZY79H/jCpT38+1cJOV75
FYnL/e5S5H56awE73pEIa2WcrFTEX3LSeMyNi/EX+hRUJBI7ENLAHJJnEG8aTE6CUfTs4HYtrDU3
lky9Rpugh/eeK5++1YQ3GGpKwDUiufBV0JhDr1TtlMuqBtoLHaR6Jx/HqPQ3zRPhKrVUw2LUoLSz
DbkEWBBUm8P4uqmGgyUvyjeycG5g+oEvb6P+onEZcZpZxe8P/Zo+QerHgUfDsB6Ipz9rHM6gqbzV
KS2r7mcIBBrmHalnSW0Qp2/81dyKehvLE9zvWbYwru4vKbzDr5qxedHcHvf6s3rsKdc6mrz/0syB
3HFgEihjo5zx9vVO+X4ccJ/InbzuzTNLfuPOpBSl9hbmNxwky7e5zHdWwsUa+sNsQix4VwHXo7In
dTTmkj5NBp0ORKhOhtN2f0p8iKfPTajfFLoGpKODY8STKjovyxR4vR5RlNBfhcYrQs5GaL6ZIRhx
1ZDbLadKi3NuH+DHnaw68l+s3+6dcTLFFtimZSkFz6YvXFNaq6WPEis0wbhPoybuNr2Ah01oXkiJ
r7d7eqYNhEyuBZUzljMfDBXQ0UIAkICRh+js+Uuo5edklskIq595ADrs3mVq6mWl1qLTDoFHJtrb
7FGZv2D79LFlzWyvddrsrNjD0hd3Hf8NZWxkZpwu0WfOWb/sPSVUp8FqaoAEb10INZSVy+ru8bth
EnjXyg5Bxfzc2YSq7IxJy+RYGU8KezPPpS2m/6gLIRicnl/PdVuNW4388emGuiduBpRSLwfRgHi2
o7wMFAwA5UrsE4RDLqbNZeKd++3mDDyX2vy5pFp4BOysNrrTLNiubA3EGyj+faPXCsHRCNGO7+7R
GohoIH5BSJyMWLZGXpz/rYMxAWI/ujajJUzZed25dwvadwQdQSBtJBWNhkgUh24zWad+79jkxKHJ
D0K3GKQCjXmpRe1jOMxZmuRJr4uZPEzs6UzVJW6n0vYlXbJQxfaU25n0uJ+9+6tSIZryA6FuZRhC
WGF6L6G1RQZebOROl1bgSjBoCwCpa2XwFZpoxE3CbFaAOy61/8Mjr159YsjUWUfhJvURCvpLF7CP
WbyrhcL1K2oSIeM5w6ZNA8m5e2Znr8qSb5a3SVBhmqOJ8GAnv3s1LO7Wd2gfdyMngK4hIp1ZbdyU
SKFuMv0iIj/mlHj2LMQDwBaT6kSwxHIiJXulVK6S8BtVEAfF8339BIsXRjVjEdNrPPEcvIXgWtlB
2BmQ/8B2x1uhSd5a04qYRp13PexzNzQtFl6rgKFFg9j+3lW5A6SVNGytxa9pds1odzmhyuwgG30T
wXM+7Mr5P3AVLmcTaur48cNgmpeaYluMbFPcm0VFbT+wNP5zbGB2+Q8gu3gJjwfDYRBREHbUS2PN
ZbDpV8vkEpNUaG7A2Lvis87JkAfMGWyhFLqUNP0cy4NwdQ9X0scs9czmtODukOKeGxMuSj6EA4PF
NJzB5UXeyGqx5dyuXho/Fu8osxRqb9qIomMLotaPPotOzDkV7eZcmE2tr9IF3G4L5PT339ukIBXS
Ui2PKHsjKOE2bC5wefahAUvRkchkBLTr7SxSeDMEX3b9WI+/b45IZpwxEJA0a9YkpQQ/g+NaWR73
2jl5uf7FItYEX5iKjasvuxuOnobGRUspuuh9GMNC30/Sg/WrBuVwFQtZXYSH2h5kEEfSE0VAYRDG
ZwDz+EhqHraCpdmoFX1MNKkpl5zvNw/7JjjZoJWim5qruyGvJ9/zGf8fPMrofJbYFjVhtCFbUe+h
rqU6IQD2xWpENIFHRrOFuOL6UR1Z+OiGH016ahG5g+6ck2HUV5waQ5+4Rcdxd8zBwcXQPSmtPDfs
qr82cCnronfQF2YCwO5dB3r+wGMQXOOmiNAnZUZ6j5DoDKu9PhEfSQdeUqYgtUT6qj5M34qj23pU
qDntwDk17y+n6KFRpDBbdcN5robkoOlPPxtDGurJjOWj+NTFhhYxsndJ1u/wLzwnOSSAE/DT65Nm
FyxW5sJ10gNGd2+fLrpqo/911yY+9syDkLlPpapl5JY3LpCtuWRxnUOGOIitRgwK1Q2IZ0ZppLXw
qoS7KozMjktYLe0H1Ru/n6lifkFrC1f1p82slTq4SKIjZ0y5L4XYdmcPobfheMQ5kb/u4Y+mBDso
ogob+jqCN1XuO3NaL/o7s49kgVmNwQggbX+eGT+uQY7eilzI5eGbIRo03XYpDa/vPN9KUu9+zVqh
6nqRzCUSqdq0+BkTycpiD+g2LyMWToN/kuyRxCzowTnSPJQqqBUyo23OYlBj2KjkbMwfoPioTV2m
uqTAu/1yKb8Txb9ip1awPivj3GfJNOAmEX8WogWpg6fKfwwQgrk9TCxMQP0dfvFXANGC3loRkSnQ
7gjSClKFjjUriIuJQx9s13PS7RyuRjRks7SDprHMPQ9LjICT3eQQmdTSLa2V+9Qf6GYmFBnAAwFr
xG+sDF/lRQbHbT1F6mZ+83e6sKRxkjlhVI+SCC4Vxs5zD9ZKIaYL+hjmETMlls9+Afjyrfm2Bgnd
pYnSyVyxtWSHN1h4A53Sgl8UPFsOh1YvYMcadjnPyA63LhOkaDuLZd9fZeAflIHSkAvZ1/KtBeFd
CBLmG1Yt9VMdShVMZDIJvtmEx54mYeTx9RP/mE+wG1LwTP3jqiR/hC8pVIU9aqic21fVzsqg+GqV
tsM5uoqk9u5xlh6U5CHPza/ccAq4Cq5ysQZPvMkFv8gzlcMmEV4Wj7Wk+vEdeYzfO0CNfvp8hOfn
cDfjMRgdWsGYXGG2anIDgUAAyRjty1DmbFhPmOaWFajFgOwiPiTB2AhFkCm2nA87CBJFsmpqiJyI
B5YAI9afkFlH9VtPVBognB+dJjSQX+BUnLyLqNelBa996P/t6R8wgQlkeDpmNGpaNIezuno8vCs/
JE43dzmFMm3VFIeIHzZheRwSy2g2xbdMTZyFVw1jDpDBKhgMjzChUpAsFCMmu9SrlOZh1X3HJf2+
NuIyo0kxIoXgcdrO0B7Sxr+p9LdZobEVoFfWmWCHXe35XcdMvCSMnMLm2uXPZJM7bYnKH0Ih8zXB
l/1//V4YPjuoqFWzigXoEEUzBIZdDHLUWjWbG/kMVt5Q8TLHy5/r6Ab5Z4QyXCDlnFqbCt7S1Bbm
QoBcPm7HSuHrkc1v5d14Bs00tVaUiYij0rSQA4sIa+saJWSBy2eaNRAyQ7aLn54tyLhkv+oTKpyz
CC983OrMr3AwZxVTyM2ofj/0l7tKS+KVoNxK0KU7ogA5l7dSNHCc1oBsHslVVDRtHfgNq3OuExk4
gwrn2DetpBRk9UqvtTRplIX2OHq8XUzEF74+RfYh8V02WQ3xRjbqJjRdqv7vmDz8u/EjAO7GxqPc
qpgbedlSlrza1oUFfqWAgblEamaH5pQKAj2GPuHvuGIqcfyVAtsmitiK0qw9dRNfYjzbPng/5hKk
ID15HZ3bHsv0T6KNQGI5XW375+9IZncdVcEYwB0iP8n/PJ0tQWIJEGCH7fQn15SVKsuaX9YXZY9V
m8I11684d5FkoI7SpjxG7n1X1RgTxJv61MUwUQi6QocbZSdZHhbLagX6qaUjJtW1RfYMZSTSbs46
YDSe5bUKfhujVC+qgWEvIF3EONljexCvaEbA7egLDZrbLbYOusx91pjiA7dtIfsckN0fj2cZJkTn
BR44182tQsxJ2DYQP1rdPI16cADkpBg6MmqAe2HEg46QVB1lur3pLXJX43rqjhma4fzOl6jmSSFg
XQq0xCqeEpKl95csZyafB2lywfvnCagNK0NLO3bym3iu4UKMnpInRqyNwcGurRmdfed8zTPKPZBW
Nf5+aFT+MKZc7WHIjkJi7yIv9ByZvnOcWPTNYV+Z/HNl6biFfGR7xFdGArrKFsNMsXwbkzxPQgIX
LjrtPPMDe+SkkDDF3RsXGM8CqnqZKtZxD5BPU9OTGLDuMzZjkuqu1Bjj/yEU93/tATq3SWADt5yH
ctvQfjM6YGrmr4NE2hFbnC7A0rsCJs4QHcNdhBFHkqKUs5//S9bgTFRJFjbyc3d2YfVeHYbhqzCa
0GJ+w7HZB0N6nPsxjDmvjXTuqmvqDgxmM4noFahEs0tcChBxNPw1CFlTnnsy7NdfwGkPOdJ5PNNQ
jkJ418m6aP3ad9hhyWrEcK8uoYPRg8qxYm9gLAE/3dTBuDbOdmwjJp6OSqrUk57nNbWutZvyYN3G
3qO98FT6PZ/aTjE5u2ROglThCTFOjPCD07OEChaYOXl+BzzvH2w9ZOJXBgmjXZSJoZf9Z+TORyjW
MPLFLAS0UZcjL8pODgOt6/yfrWoahMVwPSvjETdhEHotKalKq5HW8EYNqMIWduDEnlgnSKd7rax1
eB/BSRHuCA7zzGrOGvQltbcgGVWhPjlVcbZKl3lMCUreDHCGR0dY1BxzbzOKM7wsKgMcrGqfn1lK
M/zyxkbbCkHoQldg6arpmEiquy6XHIM2qNMy1A4YA+U+BtWv2+do7OJAGVrjGbaXL5fARkRt+b6N
nwkogUzKzXzuiDabr1JIZYsqr8r/O6HdZcBTi8iI2gcq6fv/Og5cCpRqQ2nfCVqsURcE0uSb3jnv
ydR0CeIUt14EimRd7GxqKnZvg4HKE6aa6pQl+WJM3c1yai0hQXkA5fP18zpeq9371p0TCSfFMxFr
oqFARk/x+UB67ygRvay5+O0/yIUCefKbpQFufl8Grhp+KCGCbsfdYmgPpK+ygfYYguSNeCJlgEue
cYq3czvf5s1fv7fNLNHsLgX/Me35wDQkVWJgI996a7zQdwrZdhzb/cjsK+GuUGL19IpCnDEFkNqN
/JFpU8xEs6eY4RXU5xoHsgdhMDsYk/TXO7cUhZ1PFyTJL3+O0I13fF2XBq7UZ8JIXbtgn2uBrT97
5dIRSE3cH+fzwkcwYMv7DRr7UnoEVChASdr8THzSYYFgTxof74myrdBd8e9xPhfS/QLXE5DuiatD
RUPj6EsPA0S69HIoDeJB3DmcY9nVJiorJlnaQu6OP+lN+ca7XxwIXAxR0XQCnOvSAY8SQKBw/5aM
KC8cS5hsw+9GJ9DEhOQByM3mtR1v1Q+MlGJOvmWhNLY9Oj4rJt8vtGCp4jnnjOwoqlWCnCAnuCtj
I9I5wka2JS2rhcixSlN2CIsMt9m1zrUKenbhebvaKSh4VDdRjjryH4hvUcmnylio5nRY/g9Wm4G9
/oaYyeNXPw63l0xLjC/wyH1dWjIijhmbW0VUviNwBNd5k8v7Czo+AF8zif7O+iqbvXlCfzS/UH/x
9S79qC6tvTFWZaRUH++5eJR2vQp8eu104/Yqiv03iFLi07qUD5Qazk2Nb4YG2KnDbuVnVGA5Dg3W
myx1+IPl5WU307Vrc/HZRjhJ4m4Zdcodi138ElPJsbJAdqUWxl41B1AsaWYYKK2O68niOaPzkSoI
a2pDNoXWjjWHOBluF9rtSwX4hVsXYeQpGQaDyAAo6F2ahoIfvlvQGzgsrOIBdB3S18dE8i6FpKnU
Z0jkcXm58mW3k2k0K+mct2W/CLYkzWhK01S0Lsml+HNwHSgtZruZvNS/eo1TGz1SR9WgHsYg8JMa
x7rIm1Q4kKsUcHoR+gav2phgfNamuVs84LYZAL6fuMQBYylX2oEYqs0dMArFdZL+zdRWZC7g5hKn
3t/e2kLI7GaCRJbfmH+N5bEsZ8Qf2pjhWTIm7ihG2JHXHFCfgIHEFuZJtwPpcP/bayxgNB833mfA
BGyUbHBwqvkqLK2QaG6fi/fv/JCNkWaXLOmoeIOr8ayObal9jyuMyyNSnHcFRUafymcn9t+UCiAW
IUYRd1YrR/8ylXAWM29WJNoBDtagkyZF7IdybFNVyT49llVrW8GktaE03lBThnmVdcmFLf6aFyFs
Jkea1SeaCKejJxAaG2YOFBnjiHzN1JAR3FgQrh+zoJlIksMxD0jcq28LVlmoKSauZWi2M1x9c3qh
NpA6QOuYohbxczixx72vLe5mPwBUHew1Lcz1o7/NmYyJXlkLaY2SjbpT9Sdh08HujEzp6S0MlIyR
dRCI1Ii/Pk2I1QauwYye6ChWLdIwOGWgJQM/vP6rm2ydZRv8kut/5hQhPucP6BIoUl0ud1q3y90P
WJgKYXgYRO5nvDoleFDT0byr9RhzNaMrFpt1mXIHuxqhtYHop+g3fUrUMEQmQlarJyHUXHAwoGBM
+p8RpLJqU6NQMYfZ1eiWCXtREBICWDv9HrtgBP041R3xiLrE1dr0V87OhTjRJrxLpcpmWVDpWKjX
K0wZsvHkMozarOLJFIDcWhjSn2nazH/ROu5MRFj/rJlAshKQQyNBrfy1ux6j87SGFeQC0shV4Dg+
WvDXHfKqYUAV4hiUBlEbXJnmgRiOQaBONgDIHsogMTLm1GdXTIwWr03YYmsEh0te1XcY2QVg4wxP
yaA83yIHpi7T99sgCx55UAUi+1vM/GY2Tk+jZvpFEKTu5Y8VGmgu5qPLSAv+83p3wSKlwPJWx1fo
pSfIZXvCC1jpHdnzkFL06iL+lzAB8d2dmLvSQcu86Y1xBW+8EPLf9axKjFS76cO7SO6Owh+GCpUl
ub1c/MqNaUwm3AAZrhFzMXeChyB9nSRQ7vtaMfjLGChqU8svqsvwfHZ9diuCGNEw0as1yX3VjFkI
7Z44NvWaZMDsP0aaLSxFTaZ7LiNMAyuCH75zTotmIMQL/k48RIAQ/ndBUOHo5MuvAdwbnE44ZQ3N
FMuJ4NLD1cY7VWvyJ+pDk1/icTHrTb+pxaSk5imjjQtyqGz+aI9VW70xeHh2Y+nDu+s6hHSIDqaY
ryr1uRrbi9PI62yrdymg8z81Q6ijGSiXoc1qVL3J2i0KwsB3KCvRBIc87wqVfVufB/Fm5yLKUWz7
R9Jei3XjCqJOzEi6C5EC3GaxYcwIqdxcuhf524LDeAwRlkh2k32MSmbuEMdCC7zRZ1r+pP9uNCR0
SaqTqQE4cWn3pembBj+GvNXm7+Ka3CnzaVGF9V9dvsXLd//BrZjGr5OhOHtG76cCmCY2oZifhWa5
Z/ozOOknbx7uUvTMb4efPsasGQ2dE/DMr6hBHldfgESR6HWfDNGBqLER8n5iAV0TmT7bk6o2149C
FqHOcNAMVX9SDU0sXpP7lBwcPkOvS62HqinzsbwYxpplhqP09r36dnEhEz6oa8KrGcRFowgwj7wO
c6JXnlXWwKXR6q5UJCeqZAM5Trk4gB1D+Ek5NYJQvN8GsrvWwNJPBE4KJqduekZPDeVNDg0iNpvi
cHYVxuk+SdpnrRSKcP+LVID5HGcRm16FDE5CJbPuXWQTeDIEIE8VAnb+CyK/Rm+7ediorR/ZoN7S
/BDRqdBzyW9uPnlSKPpnI78iyayHn5/wVLKT+7d5aUVGOkZSoKQMZZHLs+Xo6mObhnuReFZaNqEc
dk48njupCdWi4A8szOtB5UesGbIE45iJzic6uwSoun8Wn8J9CTElwKxEPrTscZIjTEIoHWY5Br3q
6DyNhktz1ZNOUcOVyl4jxMo528myRoqhf/WjKF+AdYLFrB999jwzrq0b96GkaqofYQAIeIRTPR7N
gSxW1T28pW4f8LHUP4h6fpU0FveOHH+7wFxr+x/i4zF6iZ1wJp29dvOqY7tXuYWumS3rjGTMXyLY
DK0vLHeIQEkva5pS6UQyvtbvxaas+KnqOnTu+/TWeyG+kClF0S5g+iZ+gcaBQgrFDT9nRyVsVwQU
8VrXk04/Si3wG2QbEvyUSpMqsMID3HLx+dJJFnTbsl1biD/5yh2lD252suU4dpJrzn6qMHi8Fcbp
7oVd3vXSqs5neO2n4Xcb2aF8e9GIGkmK4cHGEm2AFcW6g/44e0Aneco5cZddhxGyfzDyVAG8W33k
w7d4HK4LeR8QIKmhiWC4aqc0JDyecbl0iEIkh+M52oC8W/sBFfHuH47PFXOx57qFd943UDpFiMzx
eUwBjJhw/BQ0qf1TWiSEsuwglsf3oKu7xG7Tr4SjbaQKowC2AIzaZngv0Ie13ZbS5qYbA2QJ6Czq
Uy6QMs8EWAvPs/R5Am6zMFxwEJyeCCDGoTWARamT4O8Ilc09k6AMv147oq4RouJJW8BJ6271YMr+
I0pd9q5V662xv/0OrwX+3GsS/CjSfN3OdZdXzh89H0QZHANENyt4lMh5q4weGzjSMpTDZfMB2uFw
jVKeo5M6APKpd0VhzTcWn62rccEvPIZOQP9YP7PuU1QqyEP1ozVqx014PoLvlmM5ngVXLyyETtCV
c6TZJ8rA4jxn64SSsUhesYanyit/GZ7W0TKuoFKzf6oeoy7NSIpI3QAPKOh8s0lqhlrSxk2Gdzgm
dMwAB94y85yrzwOQrJ7nmJqB3INPBoxD25qHQbLzno2onRfT3GsV4Er8O39rSVxn1QGVBBJ9AgyI
V8mskKh2SF9rkVpqKCRKr1YuPOlmvFpz2trTRla1jG1jJ3Q+MSEaiBguvrmCJiruICVSPZaarWEY
QdrS7QlZE2TkA1MBV1UeCGi1+E4L3e+QLPiLV/QZas1m5YATo/AT/rDMoSKNd0q4GTKURR9cLrkf
jTWiyuNp74drlt6B3FtHRpLQPnGGIRMrO2FdwWyoE3bFD88y3WJbf8ggnWnGCg/NFclo0gYxrKul
U1Ya/HQXsUNH53EJ6T3CMn40Zesz/8UbZfvh+6rh/4iJLG/PBKqg/cBObULRIPICZ3Zd+kqKJhvz
qU1p0Ch0D7wT7hkxVxISQzk6/wLSsOQT8xd+OCieJDtXXT8xMFaWZU/Db6VsQkwu52+VQDN5hskr
uny05k6k2ktqJYu4fgv5OH33nQEa0uf4rxkMMQQXjzh5ARASA0miEFX1RvZe+soiAb1LIY9nmPBY
QW7nCFPpTJxOnHE3Cvh3PhClSHESapSpPMIFJ1K+ewvW6FUIatmEDmD3EligWmEAYlvwwEufsqZl
mK1chbBXwwh5XmL/GBZ84y6Hjnv9t4l7NKr/MJ4uucpYBEc6BDxLnm0wJy2aiHAZaq6cswTQHeQy
h07cnvUE4ppfig6UYbhLUEQNsA6KxtfMQmiJIFCqyuAOFcfQ6kPSZqoTgzB8PeNwADMKZBxvM3he
iylDvzpJiuct/r19QMCAuzv6hjlq3urWG4eMcSfRH/d9hJvmDUlTWJvRLMdKNbCp2AN8aAzPEuE9
fPmWvzw14ZnouCxWqMZauXUb2nLi9pBYMh31COWRNnYIzVjDo7GGXI3XRqP1Qap44LCnohFE1Z66
gS87aARiGE4EqKNfJEWL1hv2Aoki0NW5+fYxog3t1YePy7lXaY7dd737tq4xGEveoUDYqR0LA+oC
pCVpGphaQHxN+tgusHh7WomocMSyDDRl/CpZyH5hLfUSMLYLtQvdF12IuKSdH6UyjoZ0Bfe4B37J
sVp3rKAIKuEHUd002efqb1kCdGpErrqu6goY9MekjKb7O4kVsADhMW40IBZcglFGOBAl/Mu0/JLe
hmoULlqMAKh8qBmvVnTD3cEkyFfTP+UWYna9EVFc6RJ4736sce54sYbHClVqWhXmQ4H3qWV4vdcS
vb51+Y/TdxG+jWifPpgWYiTxkwtIW6uid9HzNK0RYS2c4wbmxT4uvhqjucq6Ee79EpZkKUWIdap/
rQEmFmk0CXrz7bY6ivmRudmZeliL/05zJnSSh2qf2ss8M22AosWBGTolJmM1tYyPXg6TAFn/IQaK
/cTpNJWpyeKvYLC7bbkzaNs9d/bu01LhL2p0oZn8M6JOxHgVH6RGk6v7aVJXT4aJvLK4ZmYVDFHI
psHGYPMbWZhNRcelac2JezbDWurRJ02JWDOg0dMSb1SOTCSKdn5NZyijda3SA7FlcdkB0SUXcwTn
D8AJYyuqFi+MR6BOW1FaTdbXdsjeWq0vdQ+NinYJjQlP4kiGAPr9aV/U7AW7G+Pa1smGEigAgN/Y
AvXzpKfjFqccsCF725s5b9fBQ8iu+JuqHix6QDmiW9dMCXywbJCzZ+AZW74Gfg7O5PKTfdFddcB7
pIEOr5xvnxyFLH3/WHjDp0EI0VW5l1M1F7x2YsJ5wO2XJLzZ+h1yueoyGBKXbOqKvjYocWx+ItqJ
n0/NAlH/fDwyZcWh900+0FZldSsgo7ZkbCaq3xB5BVBZqHgh6cu7Bo6G+2yKOWPTIMWeFWyows3T
P+w1Up/smy/l/pY8GaVKT/D3ujin6ne9uMghKBiK/nT2LSDv8VrVOj0xB5FElVlH7XmS4LdhkU1L
SbHKeCbPcurjrILxx2VWeFxOAqJsV7wR+JF9bkup7CfAZKJMumUsJULsXauRjWjnFbOPeXCLlaUT
MDMKIDMGOO+82Fkvr2pNWUcmG2tyrQXVj2/gwtOWLSmrT1NMv7Vc/le2g0hF4Zbu0nUWqnl/Di77
BOc6BhlLU14qkM8VKn0r+gb/2fpG/HV61eO8WzJJ2nvcsAVQHvg2QS2mDYqWlLn5D9bADtMOqwdF
WZS/D3LCGsmxmNi+qfRbQRo8wtXwOcDeNduRBm7xOqiamMegI6QCtd/gNJ+yhuFg0fy/WbdPueNy
QAyzUtEWOvgihmtlWOoA9Q9NbhsHNqL3DaY/hFKlqiQnayBPTdzCOm0ZXO5xElPYRJASdJLFG4k1
4dZB1b0Jjsz5tKFTl1WHpDa0K8rjqQrNXIgd4YPbb12uCCJftGLm/iyxMTonwyrkyL3hbZRUoep+
FdMekGLL5bLFTRb+qNab3d9HkGHf6FV9yVLhlOApi7rtgnNGPROra1HpNl/dNRRZMSPTaM29nGDY
0tZa6oYYx+he3jd/NwnCH7cPRNrTljVrMrgtz6+qtEbZRaHafyESzqwZCMUK5PDBRHEyk96Da84x
4VIyDuGI2gpNAqclIfjqP/Qp+pk+vXjvawpmh38iRVULKqt2oWFrmnUi7VmMnY4sYAM/D2u8RJ8l
8Rt3IRu75I1TTq0nR8aa23Ern213jtT4maQFVVkYSd6JqXEtAprL+uAAYGRcUpQQsT6vtbUl2FhC
7SHQIDIcf+LbdRyBr/j/dBYZJNuYvo+GWUZ2S+PC/s6D5PjaBxgfnkxw8hpSYg3Xe3WNC0ofCnin
iIk700P7ly2XybJPumQYuGJcbwI67blq2QR3VEBIcSQR2d4/D/CUI+xtmRmGPLwYAZ6Ow6jPunPt
PfGC/7cwSLvlFrzMtPfoYh641UR0S02y9x59MaH+Z/cEjKDzaLqoODOZVpVJSI/I0BFnEuZ6U6PB
gJGnJfzYtGnxaf+C9LcvyQJLKlbhqg60Iite6QhhSMwGjRVSB66ozgVaazh55s8oVCoqettI4q65
TMv7xIbn355jsl4iGMbfyTtIfHE1wx6FKyEJMOokTtqAQ9AQNaaBQnaWUzhXqn5QIjHNTMgFwgP9
t2jOD1+H4eHwBhwVAksgSgtld0OSGgubDNOGaOCVcQuauE2lPdl+MaNKmx4Q9eMThzoevPgM3mld
7+J9Q9ive3BLHLbzxG7b0z4nVIADh7eI2/eT4ZPUrRi/BgIarrWGkrpSBsd9uWtq889T0jcmPbXI
atSuqZWQglooO+TXkyh07P42pTRpOPBzeFkqOGhLsL4jtClEfvDl4LF4AE353KAcxqUduWSSS9l5
JtGXF5+RDgqWPjTBXH29CyqgE1u1jRDWA3fQo6e/mhHrAb0swwtyg7KH5wxtHh8wQNcuWd7LbOkp
7dwHTPLAf1OfUy+ChjvVVzdzSzXGvUpLMgty0yZcKVZsTzkE6A9IAmDY3eNmKGvfDIDxVvZVVrYU
Jt6JAvqDb5DRSdpw+B++nt/L+qazzd3tMoxsiJDiwrWCa4IsT1Q8Ca4nxlkHI5Xr4da2smS0VFwl
UVw9y/HzGr36x/rNj+OhfeWdqNLQBA5e/1NF5Mstb6D5x6irBOKmG8Ni2Sy+LSmz9umGT7ZsWKzA
qA8HUFXxxPxrHMPovqdP9XCMKamIsDOQQVajpopR+MYhk8/hTrHxXguQOxyfbyL3GOewXp4DKyN6
/5OLpUrXrBI1L1a6DR0WDwXiqkZtco2JD6BaEOczwqKXNVEtvVJUlW/xLIMBx2YMECEw2qT/q6pS
1ezsnz1fkwPCEsfkXYS+D7kmuOikRwkfr3JFBa7iuoWwXDCuXJ62VEpSfYP9Y8Dw7Auj4PasqWK6
2zftDx6RLvXL749LFjFG6z6ONFpYhHfhI7OuadSTy/YWHzkwy3VWLbwHBkEAFjOYe699swz+R3Ki
O+NHF9yBDcfv4NDlas0F47q8VG1zo6vrffO8hnJVQlrDlXD1l6a0+D0nrzy1g7VdXlk9PoI8JTXt
nEU+neggyJk8N0zXq1j86LyvMNftBvVF3DdDe3O8KM695TL24KrsNZNuWbIGQb5D1XI8Ak++ZY4W
VU+mewJcQMlxUFn4LvhgGfHwoRgLVSx9zEXieEY+F3LumjDwNESeXcyBEYpwJjsoMhEZec0CtGaS
PuJP4M+qEI4BhvuKwfnEdGGCm8r2PNPloqsNcD0Ah8Up5wqXDWYH7DREIjK0puEialfm4Bvmdtuj
+xZKeAYUfn0q7xKcKOYyAqQZdIiv306pQXEqW+l1f7J3tE5tfRGi/if7hivINIUBLlNYuVJNk6xc
ywpzNUXqnAZrW4yiGaQzG1fz9+F8iJ8IPMCT8i/HL9NuE1EBwvMvfSScOa+JpY0k4oakYf2rFbCO
X5FU9AlmIOZ7ynwE+gYdoIMki5Wjt0ejZlqYASKC4Cmuw+6Eey+LPXBBSWpbjfMSEdEfmbJdMSnY
0tZfK2Q4mrtHfcx1WSjrV1OUYbznMUU6FCG0rkWXwrRPUWZ3BWlaITXjHbKkes+cXo63FueFrOsC
CfNa0u1D93DIx/x3sXx6NlaTXztQPxMGJhoNk7eGyRQqXkbqjiZZHu0Y4GkvyWFUNtOMWjQftiIY
cJCXbuKhUKIivqyv54OV75YOy/+O1CCQVEiOi3RwNjPjKDfBEaGOE7Pt6Ek8+HwUXqEPCapJg5/u
7c9hXhL52duhpzgBQyEQm4wIP+1C4QVYnT9r2TUsY1bmTeXm1fgE8QANTEx7eZetbNwSAQdED+E5
wRLoHaiNhJJlwH38PZaVNywv2cCeniEdraQvjPYyij+Kihmm+P57P1G3jy5nL0FS9E/k8NL/eniK
I15MN3CsSiuNDG1OK8D11/paGO0C1YtdpuYITwsS5o4UtZ7HY0njyMrXERPRg3sqW6EjU2PFlGKZ
8ghLkTmGAFGlkjBLg/zdy9U4MH89yjy/f5hgyFkqK6K5GVmYyV3mnIRJGig9DyvC4OwxSSt5L3iG
mCk0T4yYoSL/gYMMtsyeroxF0bkFTEi3GE34uk0bpLriGPtOxETZlCZmNenJOfYdMwR1dYnSe2ZS
pYp1yJHNn1HRyBHXc7rs9EuD5jebqk34Etstd1Nj0em/lQLjVQUnb4IlSYuYz/QkYt8AenEx9iWd
SwlNKmgSTnnDc2PK5bTZojn25ZK3M4HhQ6vTfb/GY4UZupzLIZ/DsUcSemjYgMKDJfPxSal+geEd
IuMmUbvPV4vX+7/p7i0fOmnPnGw6++L5EjLPbs4TS8EtVQ0yugVibGlw50OL9VwITRVG0M2TsmyT
4ujygsPmkPdO3JpEyZtxbZVbDvFmLVWLYWGjjVSy+cOXeogBw0ZCpWHDrHLsChx6yXUhGd5BOZbV
tSJg7FFSbGqiEMKdevfBUfzOqDMDEtmYms5F3zIv9UYzhEcKpG1b2npXxhkUibGAfdyHJ8dE33gU
Lq4VzveSMbKSfM14oUj00GMWf5Ay2x5N9wvKLPA19xVb0lhsaucZPJ89iVn9feMq8EWsZljFlGhf
fzZqdoMiJIl/JBtvm1x/l84Seylvid5gT3T4jm1dAMga6V1kjvRo6W0p/XVg/EgY66pDhXrOYv1S
JzK22mzzGSexn3iUStKNA9eIsNwoccqfNhe5gKpwZn4cZHzGqtJ0MYhtuNIcd2+Qm4j6+0hnfklR
eptFSR868RNntR6ohExLV1tdOxhUSc466y6/b/JVjHF2hPKoRepdUZbr4SQVYYRnS7brZ2HcqDZZ
zrLJOxte1tT6DhvE56cc+CDKKLbKxghxtfuNQ+uumJaWIc1tcdiX0vPhySUrW0PsBYrwLeO1ODPw
msQtATcF7QcJ0H1GuC8PCYuEaYSE2UKDROV3RxHfvCqgPz+8apM0qwOxsntnNgqTT3tvUUU5YdAZ
YoLUOyc+6rDldGefD2qbtuUAoKhCVF0pzGC7f8mT3U9bWPBBwGoU+KFDSct1e+PHW/+Bvu6sRsnn
8yV9dszBjXcILPkK/cnJ2tlsuak2Pf65MQsYrVjocBFGY/+SIipwI4F9G/h2sRJiIemdcd7/VjRm
Fy+9yS3e1WwclsFUwES8YuHzAfZQe3tXnak/i88Y9AlNNoCvAZlGlgOgAtg8hOXosGRDsUdZf1pk
Jap20lUWh14WFYlTA7NmzffEzmQ5jeB8fs8BEnizMvzmmodvPi2MeS+FMcqLcoOzxz8+Tx0uN78N
yvT/NuOqOGwVCxPLc0IUyfvXvf/QhvHm5toyeceVjq0O6jZ6hYjENvysF0mfqIBnmKfHE1BA1A01
8uJeKNbfcmHbDlM/sgZhNcLvNu/x122WWBDJFMkUd7QVtX2D3mYOO6pvbAVrk+GJDciyfrEAZNgF
HOWc/NkchSuDET9m34OGyrdkMEPONFIUDPLTZp74y2CRf6jTuMibRdz/XYsr4CYWFaY0z5hRYX+8
4pLUxJl6eyP6xV4VTP48YWNrzEkmyzIdNq0f7KI7IAMl96e90o4yzvO0VwDXI82bXJosy0FG2BfE
gjNzpcVcaE6GZkQAtYXqD9ttHBO8WbUheTf1qgGmL93voHPS2gdQkUJgczJdoOXAz4Nl01kZWpDl
58XTQAmFRynjMu+m1Ein6mJuZaMQssGa4KLNhyHbmBL98G28hqZueP55yvCrlieFtTE+OcVpPN1M
o9RlKJqUNJhG7Pyf+ktTGtVPHcp3+uJP2nROAliq1uv0/oyHZRGIMPAXO124d9RiPnncWlyXOG2R
V+0/cQ3CCg23GLu0w8TSP+CEzJWjR+kuPZ4XRFvEz4zt5rfYxkvlgF8XYqW/x7GLkn2OYXx/JHqN
VQ9ywOgWlNqkMtw9XFROJZxZZ7eCfswIRJ2C0tdFI29D/jyFutkQXNIRKkKVSe0AhN+GxdxnNjkO
hkExEqTGxx4OG45BJWFuM3WH8n0i/DFZqppQ/vivjsL9sMDHucAm6aWnCeLWk0Xoht2cRhvFv59x
M6gSAzlPov4C4/n+eqNGJcGJ7NFk+djd5vS5OvnwTNUB0cKCKrFk9oEdF1hF0dmvSuDgmY1Clv5G
nXGBBHZKnOt8JsY7znw+XFma3yyo5ibgGSSM44iRXnYwYMNO6azmjbIS1n7cMaDS7tDYmXw6pIwm
7vcchC19O5ziGYgB1zRp9lNipDnKjxN0rFqCCnfinUiC4OKMzVtTpmWETLmZxIwKRBkBq1HbNLbV
WmGtrG1Zf+k41XodPEl+6r0fzRnvxoULWjjyA0N2vob/BPFtH1wr/9z2unqanJtuFvCHbG03Dfyx
6XvF3KgTX/OaFxafrBGKmxuesIcYOzT6oX8ca5jcpP+ZZo48/Y5AdMkTqosQSZLYdi0onf4AUfqC
0N3vcSnGJMvKkdIFVVK85RCAQX0DeP1FZINFLcMh2GgiYFd9DjnzRXD/t18pegGbePnJVl9nKDqE
/6bHst553ZlcUcZHjVOxjvhhF4EO1YnNPJkV06M/SVxnyiTz8C9lkrR1FwHVlfahsEuAZjS+RkE9
AxBLLzhPbPkEZ/MOcwAIJAL4lWP9MVayBhD9RFqR/ET3PiGkFRygNaqR1Udy40wbtZFHivxgmkyr
OgoyE1d1e60MK57B2yGY2O57ZVU0XJMwJ49EFK5YP2dErr5iDjbzlMCO5StNjNzdPBiBrDH0qIRl
bmzKI+JXKl4NZz6IWaRsBS8FKfb48S58xDAwsjdDOPDTHWru3r1CYAgBigX6cdfwvevu+wi48Gjb
gmvgHOUNjWnVrA4rhdKvU9KJfWPX1UT3NOcIKunVCLfhKwtsavz8EwgU09Wiv/QUjDfmLpSiwvPL
iW4gt7LtmlxcCG0sfCP+7TwtlcDDn0dt2lK8OiqcZc1vAjHAOZlztc8ENqN7IFCNS7fcmeDQGW8k
Es2KeaS5h4ohA6JDF9BXf3Ro3v9acR0cvKDfDC0zaEuTNbglmrI7GYFuR1/zMFeqlOYHmQm6HR8I
RVw8ZdIfiK/qeWaTyX2k94JRr5iOsVFCoi0XI3VHOi0r5TUVS4VLjaogub6rVG35aHwgFvP3mqWH
k4bS2DgouLvaqVkCYJt/RTh88UIrrAXX0v5zek/wALjpAwyHHx8cpeNVVnsXlsHyz5jnpHwcbwyF
JNt2h7wjNChMXFJbFe4FTZihaplQmoW11eugZos6oEXhvnd2VGsmmgtOST6mLrWUpNtfff6J7LNg
YJ/B9IlWCSjilckh5UJhzWG8AXx2T3ku8U7yE/M9boezy9Na1HUFYx0eHQAVVk1+ytpCn+SWGbEu
Dh8PnxTtAnBRhg59wNIU/NedS0hCiuE/ysc6e5LeAC8+BCV55RyzG5IAEFDDAuil6Oei3jsE1T3n
fD0PjD9p3V7bE75hSAm9z/QXlEtC7IPoNv63DeoPJvCEBgk3NOQuFz6o16uM+YPaZe3RIFGYAZcu
h8Qe4tAE8zV59BB/D55PjWnhJmtkd6L83aBkdBFNGdRVPKgUOWAaOZbsbNYOc3bOjbCP9vKmxlPa
+4iaM0AY2U7UmWqd/zqUD3iEA5UjpyOrUf4NYFB2QeXfxlR3fRB+3KqWbfczuTOsLQJ+HIebeamc
Ut0TNuv8FQUYDzaJV8VzV9fau9KtP0c5BnEmWgNNsP/innZzowQl/td9z+75dIP7wMzFGNzih5el
1lWZ8oaLFwE3urlEMQbfxvoyRgie8+vfPzHF54v+yy64mz4IyvDEpHdRpON98M7S4joj/JGFiWrL
kC0Vz5e22N5iPIxbpd8irn9Xh1xdXQPtEo0dDeMxBegvkwm17vWWXjpvBfjriRRs4Cei7B5z2jvf
KPBkMT7rHX0BwhDoGa0hZOIgAKs/NCaRlAAp8EHDx4Y/gNrr9Smx9AmlylIJeIrDJgyEulD79IEk
5dVQlZfoqX60tm1rjdvFg6k2mIUMuqgEjPcWp0yJ71W1peXqEarFpnqpMAX6amdKqMmrV9yVRkyr
NQVHt6HVmldpYGU5DE7FfAPLgWpaH6Co3GTNEg1gBT0gFEDgmZO967iFPOb3cPfxIuIuQPiLEf5T
FV8EyXN217jKjpeulHWRz120Zc4nMZS9ftCC7sb/tTMCKWxenn5/i7Ya+LbKBEla2E3h06JAC9y8
n7I9rj46qLf28eAJHVKvSZWuQAAyVMgH4edS+81Q1edHINygLYqvBYKwOXMUhiaZoWUdlMtpD1g9
UV2Fc8XgU+SSPJOD6+jwvZnbgdYOZqPQ+P6A3nyf83c1IOhkrLd00fIqiCYMyjWwXSFvZPwt+2r6
ZgT20WYFfuy5EdbXMq0dzJpZGQ4QZcXcbCqsA71qXV1ROGRy63PvuLJ99gH3DHM4SQcdGjgHFLPh
gCFJ1WRvm46shMs0boCQ20nagPNDLZ8eEcLa2W1olENHdDbGsqc30z7cglvvTlcS1Ot4YuNMm4Z/
fC9DX/4a0DX6zOWwcHaF4Q04q9YP2t897IpoIg3eZ5XWCO57L1WOhtG80lRtBK3tYKgTABmhsWQJ
BvYkJSZnsfu8IddDWZNnO0LWmgLKY7P+6XdZKNKOGl5/QJtTR/2Lr50D55jRYVqn/vXzaek1K+jH
4AmXvsKsoFtnA7UnT0fuShITnE2T9XlVuJ4ACK388zZnYtCLKHilJ+LAyG1YvyRYK5hNmSIErAYg
YiMqD1wT0qIvnN9LO/FaRsVPPUJzIPoo/6sUnMogp9pfHzx2FH7n4Jm4qWmxEcXBmZTLrHOyLKRm
cZOsdNugC6uXbxjL6YCb4M1L4+d13m2TiypySOAccnvUq4paYxtizhFeelUEYXNMOlsEuSIRk+1M
LhOSQ4PR8DqkEIvH4kgR9qiXdYw4vUpx4BTKPNsTev7ZKe0U8ylzf9SQa8AbkKVgIiCEyG4g33Gg
J1AkdYhXQt12nmFxvHNUVDfiViSyTCa4fZCxSFN4Fyi/vCrOsKNp7w6M42x+V9/fcdP1pVWoGRog
qBe7PPbwCQmelWiwqik3fMwGQDdrM67KuO2lDhS7IagiBX/NstDQEjpe850NWgtlKaMKiUTUDZIH
Q8LB1edcgB9+NouLnsZfqJZtm4nM3rztxA2rwjbh9lZR+CQbWYsQezBeHuLBcfdw0lui5+V2Q7yH
GSkopZi+fHGUmTSAPUmynX9MrYca0eAL01ZEMZTLlFu7kiRIJCb9bq9dM5S27DHogsqyOf0SfXeJ
oRaF0syRNrI1sY7CcQie7iWSsxWrFMoe2TJHBfE+NMy35v1hSDb4HI9nyaUI0IEyFn3DpkiZcn2d
vnCiYf8UeUlKzkJK6CsiUSTzqr6TN0/f4t/R/4xoWcyDX1LWYDuq1WTmEKC4eMDyjYd/WyGh4CxT
uPckSHxUwp+FFcXHUzMqqUJ8OXSexRu0ykgOj1FWpjvw2uJjIHfy9ySUMyRWy2Q/UqxzakWBNleT
eX+Md16bkzzcoc2rMNvA1Z0U5TYEAk+QoxbX9nyZPGhFm1KSURszl/uISnu3thygSMSW4Anm2S5k
ztbEkQYyXQI8e93zuwut1AO0batf2LvlP/AvRAWwooiJr6nUDF+HyW+6DLsysHH8O0g5Por3Q8xg
wQxFQ9ahWBEFq6gtmIiwkiZR3wVU/xneTEaaKlhuh/qu06OrjzIiHctVObeAUIwoo+7diuceA+bX
gGmgwq8tnFyfdRZi9r0rpEtYW1JOgJOwFXjwSSPjZdwB9R2Lsc/rsx1KA9SRIsvQXvoN658rWCVk
mqHPPpSH/vYpgE+JynkkKSpFuPoE5+/qn0PseSXyrUay0gPxfA5Vp0ksu+wLFLmjgYDpAtT0FEyb
IFFgAn7zpZLaSgkgELpU5zxBDPthqvAKHJqR6IUVBBQBU1UHspmxTc1IMx0wbow5zQX11fAwMVTt
DkafPcpFQD0fhEi0RJ7eg36O6NfC4Qf2ojOfa5GxsGO0epsJPoyq9n4NAyo5AG5AAH1DYmHOC1Pl
cUkXzzTHpgeIrEVNzycAo2ripsLjhCT6b7c4jxkMXBljKziblaZo8AzrRes4vGPUm6Fp9jTNWhLe
6tDbG8Bed60ClColmB22Rd0QeEpupEo0u+bhUMzlmPUq0rPQn4W+ICrSK2zgWsdHBnJqA7pFUdMD
DTHrqZ62JBrQ1Q7+5+TsmOps1zSNYumDrPRrP/j+k5N1wmzAnApzoPXtmUaq/x6aDvhlwiOOvjUF
kRiTNMBR/8Yjji/N0fHNGYVzhGpCqDnntt49afptVd48otBBTwl9nij51BMiyhoHNo/aBWVHdn5b
z1q0vN+2DAEcsJK74N7pb9boTDlZClelUJlE+qstgqhXrw18ViwPU1G54FYmTSSnPeQ97P+UaXQJ
0RXSeyfUgPMIjoevfrX6hEs39jB+W9X2pOf2VAXOR1j4atyrANlQwBLVLeTZekD9RRv+or/ubO49
q7QrhpINPv4hNJQqy61+2oEJkEV0gqtllATxyOqZVdg31SJMJF/RNsGnoHtnJ2bVaPkfNY/GIPXI
2driMOh8EgQFIRnJbayyjn1GhdvC7QViPrwC5uotWJ3YYP7WQJJ9E0rAQ2EWob2eYLWrYSqtpnu4
jgg1Ap/NiBrAT0AodxHHbOiFhrujFUY4VVclYCFgTr0jl3tJz51mkr/ejMzmE7aROpXxA6zDJxFG
fz7r6e4xHsuHnQnbrPjG05hEJc0rYWGmxKvIyyPQHCk5ZaSEVw+RnXx+2wSnUIWOD+grQrD462ED
D4nJIv8Lf5vHIT0YMJFMiBX/Ep3JV0rjq3LtHpKpgb49lJl4Bekl9df9RhNeCF6Pk5mr1ZN9Pr28
I0weOAnP2ti+l/fPdsf15j+V81Wk7AS7vEVKivAmspSAvY+ZT2nDyQokHPyIA+Vzcdc/ZYcPJyTC
cYxA8c5ZNJOyQGCevijpJE+lZc3EYZHo9ooNFQ16u4pYg1qDAthGKnRPK6G6Tvbv3IjHkiHOfoOm
aLQMkFGdie78gw4EphbJElglTihkoV+niasfc9RPWnblw+wEr4sjdJGzRr4DgVUZuWFFdKA48JkQ
kueCyVCy2YJxkEZo13iyvq+t4SRxpeK5Wsw5ZNrPqCLVe10poRKrlOMSgK9n6rgUbMjwdrHph067
c1WRs9919926wYeLp/TZ8qQNaBXQZYAWvK5aWFVV9pbKXWOwX0IN/in0hGwLhOlTVIgkSZ0msH2d
rdzDCJLyG1BMa2Q1Pt0Xg8F36C3HlW6VR70A2WLIsBNPDjF6cGqru3NvgHy+ymYURWuVaSBgpoeZ
WjJJ3zaqAv7UoG72wzyUxJeOB0FkKVm/S4g02HpTnWvshnSa5/XLKZE54AthNUSR4vhatKxvOCIo
zW9m38jRhKPM4iWrig7nzZPOyLE8MEeqOQdqsKIhZuEUm+uJDcekivdf3xEsh6Qr+7Hj8eZj3e9B
LC3E1bSU6nZxpZ4oiYBVVvT4pIwEtpvawciAdTmjlGiSAuWz4i8zhtTwlsKcCAdCHpTniT1bbWEh
0A4almrsPiA7x17DGAe2T0XtEgcHPPzj+HjUCp2Bc0Rk0pimh8OQViJAGB1LvwiiKBAxrcV1m6c0
H0v+L++Gp57luSb1BPlSQ6OHUCC6t7Cs9T0Fk+irG38ET8rRg5iTslSvkOyEL1MZRPUrjBJGcRdK
kCR413ySR0b3nm658VB41bzBSYb79BwpbYy9wTXm0mr0GZ4jTv+3KfRoWN7Ocr4cMeMG2VnHSwP0
QIXtPKoUzNw3ZnOv3RVV2+eZKwiwCoc2SrR7tLaKA311+gX6l2VWMuaH6NPNpQ8BdcuOMhW010eR
2lqGeb4fmKfwQ2HGGnp1yUOBhk9i7PonHxGCjLf08LSaHY8tb/lI6NKPXZ5p/D3E8x5NeVImRNP5
FS9HuA0SVV8qCt9IRPWRPDmt+sK+FLgmJO4KFEBAHr7jS1jnG/VVwU/AMQd20LyQt7BFBO35lF5/
k0zS56sxGRxrzypw9CsJ3e7OH9NrPdrNkie3TYva8Ku92CUXw9WsMoNTgebubnSP/hydgQVNN0rB
6fuTUQ/ZMFFftNwofp03Ct/UMbsyGO1lg6q5ARUaMQ0piNP/cWgE4AZwMoaLUjDuZcF6v4tAD+W0
tt21OrQuvkgao/T7Mg/DiCpRiCEusiwJHjJn/85BjELTG4VmMmNsRx1MpK25k2ynWJJsMlQhXdHE
Jd+K5JmiVv5LmkH+5DO7aSyigwzBl+JDdV23x0qqEHdM4kDioXxZ6NjFXHZw5UYgX/S4R4Fd8qCh
6S/irViuhd5WJiNEvcOECMGnFM2f8GcOP1baOzBMQGhvnJgbfRo2VbmpXRHSsKSg0f9rELj78qUg
w4REpSoihwmz2K090ItV1g53+ihmJEFCkUyPorQrrqo+RfmpToyVFQtSPCs4TwxP18QxVLgWeqoi
WKafn+/nEH5tKPAtitfYaEhqljwWhB2nunDS3rb5N6MfybbjwleUpZHw75UwDmgE189xqXMv6X1g
thg05R3B7uRo937QiO397yd7CcN19QasqpGNrjT1HChE9wAPaVr7z1QSw3Ndv8uW3rZBjmA6QJNN
QdY85D+0Ohc8hv2k2eNFakRfz/xDBFtHRFczIGaQKg0x6KR53k53nm7/Y2qOJR1v4js2ML1/qiPC
az9OEWNJZL9HktPkmI5NiWM2mlZkfGURWxXDnZw9oI9eJXbE/DjjizbqU2h7HavgizJhuCBrSrHQ
NUwP6Ji2HbYwPVBn19gpvOiw5cilU2nweQCJPvfTfMzzoxAdKhecveA0YFQ1zUOVLyVQIMkWj8ID
lyH5bcow8zMXOhFU87f2LXPRCApsCl/8rCTld4zmDBODftXXS1UPbJPTxrECjCfK965asTQF5wuT
IITUBULTM7jNtnAJbwERoF6kI2UPWCV1ogxJ8d2hDAoS53HmbO5+q/nk+58NZLZnH5+MBKRb5R8S
tSSHHFprRmiD7T7oGjfeiABkce2OjRufWcF9U8VZHRc3+ExvMPKlkk/iu0Mt+i9ur3iKPZx+yRav
m/+DaSTCmI/kRHNmtyEKAOcBzeYu8sKqSj5lLHM2HxOGx9oJbZFxEcbtreNbF5ZVU9utE8s8kpiO
cbAD4S92Lqb7ti7cEVm+7bUIlr5B9Ic4is4nc9fhwVLU3ViUXvNCHQn0ylDpsGq/L96Y1tgwxh57
4v2XYqIddllFBViRK21uF83ulq9CFGnyteQTh1wx7XqQMQ6lS7v4Z1skpKHu0qMH16/+tP5qeY0Q
PVDbegPMShact5+//5dqW1E8ymYzdUjb2hBcpD622CQg2wAb6ZyXbFlYp6GJT5SsYnDULNLvgb1c
aTgafLZIcvBBnaroJUd7qK967yin1fzIPiuTkbQzCC/kls68eWro3H49TTs1IzP5/2dOG/LBl4ud
+AAbgPorGCPDwvOujJFPOUjN/KiNwlPuk+Tin0bel2EvyGW++93GEAFda1tNqDPI91SJhSHcs/U+
Uenjg+JTP7EFFG4pWRbSh5e+ZjJe6B3sWZJvXa/09JwpO4STJo9XcaMY5yCcTaUX4CxVy/1v//ny
avwCEn9IqyHeQ3soB0+c0wGDRV4sfivPb9gbiT6dMijwH5t/iT3BkvBk3T0m8SkZUoEBt9YoFTF8
smP/D3HXDuJGS2s6/d4tq30tBTPH1V88Zf9cwLLi+y7mQX65onRePglwuIYAyvN3pQB8mYfN39x6
Mbb9OzP5S7Bfw14Xw6Hhlq1yTUZR5m5iqTq42ZXD1YPIQb9lNdkcZglScFTaM8UPuieWoH9m6T76
L16ZhFWukvkPHjx8s6e1Ic2rUixF6tj4+O3p3l+CoqyxWjNqdUKPRBtU5nT9iMWvQ2d2QA4I030R
OzM26a4zUiZwCRf1V19pQ/n92yns/cGxZrMUErVxrDgcM+2ikE11maBFKw2SUIVeq9R1a9/JE59E
IFoe3SNix7ffVCd3rcpTuHrHRe6Qh5RgJv8GjzJN7EKHMTQ8MzJtkNnSwn25zaryIzO9zx6kpGyl
7IXgClnZeGSjrM66zUlHjFCoh/M4DVmaHzE65LAHEOUR/CFrbheHHSzWaxQQdlUkbKjAvBHUo1TH
TQz+DxjnnPvrxwRjuaICiFYjhqzLd+YeK0GYmJqCXqyB6Zlq/2lPwzxFQZsi/g+PLdaBwpGyAXBP
kG5ZNlJMuXEp27x83Uf3sFgR32TRxC6k1MnsQnP6MwQILqLaiO0JNZmmCj/klro1I2uGCGh2yRgi
dQO43oTqcBJBo87ys9A6E+zqmJ5xcVgNuRg5SIWnJRtYz3uqnGM3AiSZfM1SJfknQVCaD8Qx1haD
VFneTc520o4dypGvQiOPO8+94f96wyd5DfYF/vGNRys3gH7oYC+Kl9G1j3KVfpDPqrwPNu7zMWho
GHKttLpGo63W5NWfpA4rROVeY32T5PuSvrp6DBnLsf7T4NSTk79XM8SR8J/yPLiSWK1HU5o2IVtR
mQ9GoYYyliBdpeXoRSnUj1b86hZZa/8m9sJGfz5dR08+ccIxHriVQ9JkOgPL+IoR62IImJzpxTRP
2YAqF/6kBjtkSpLjp05+TjzQPKL7W2uRQpT0GqEuXmB9l7de3/vQ6Xrq/8v8OhL7hAgWod/NwY4n
ot9vgrWsGOVhzBp7FwLtOV+KPzcWDYKVSSvvBnUpk1r+JNU6Y1F7GBnijoJNd/HIYj5wmO69Vg/S
2dxii61SJj76PeKrxiQy6/a4ZGy5q4Le92QgjoCV8o49qBi/2U20GDeoie2guNqti+2bjLGapfl+
IN8Enx1HMWQyBRoJa25D8YQHZBHCn1LimARQjP7n5Zljgdk59c0yqS7QTRmIdRkvZWouZMRpHe7P
Rqvqv3QmACCxD5di/0p9wRQCi2LgTB4Xl+UCtEDkT31C7JgXAkY91MMUsR6CGQRnmVDqnvYQtTOW
J8/WFRxpqEYmC8nUMdFXLoi8yIS9/lwoQCqCN2GgtXePEOL5fjV5m4eT7nTUNo0EtKXL9kL3lw7Z
lY4yMp5ihky44KqMifU3wDrZRx3wyGfxjzf91HBuuojO0AkNc94xSKyZJm7G1t10GssVerfArGvB
R/FDuaxtb+j5NDAo6Ku46JXtG4r0+WwV207x6XQTGarkd+MHu1d5F3dTRi3E/7LiCmKxlm+u+GEW
sTILBnzpiBI7iqEtaKiWvcJu8qfkYhqg7gzrLBc50OeTPboUrzvLpp2nwiQR3/VxGy5Pg1/UKuzG
/cfoX3Ela3+rf22qyYfHIPSsgAMo2zcghaPDtwGUkoK5u9wkYVv88xZyGDovWc0KxDEb85PY0eTD
uMEplVwn4tVC65osewbAeUNricibhINlV+YGnmLpI8J+gT4JmCZgjaO51z8LvsfOhDOAtVqqLnOJ
Rsjufaw/pNwV8BbyRR6LyRWJo4F4OYVX97KjlYnKA/QpssXzcCxdYsC7nSBzEoKGFrTLxHR7yAsY
OE9bCsDnNpWOTmDOAqr5XvoQv73EZohLt4mQF4B2bC2+ixkzxVgT4M1nQughY3DRu453y8dVukY7
7FDdUTy+0ZFSsDe2RoCOGPQYWlgbMXG7GppXtVdsKjnPtZf/pKNlvMmi99oQQTw5gI+hy5pxuNtQ
8P3sygHPQNci7cxhM99iyhSK80rQXyKpntL5wund3ZXzpIQQNgYTL5XDxi9Q0RrDr3cXwZFH9+vi
ppDYBTqPkdcRjoeUT3T74V5C/MuwX5Y/WzK5Kmr1TtR4QqnkekvSWx4g64a8tD30o4oiF8C3Huy6
rb0M/dUrIkPrE0ArNFGlyhzJosYfQlDIRibRWUYzuVRZQIe/6IX1RRF0qHU7bvx0yN3Mkq/cuCiB
MfizxDGElerlfrYFXqLenKtUKMe3oJOP6y5uDFnlfDYSKEuwUhdGBC1B1kYc7gkuF3lusDEJWIQS
BqY2bhtuYjbAw8jf95cySKPEIv8+smng8qGbraR8vBX4XM+S/90R3byHKlk7MZmUOkFNa81ymBpb
nakbP5pR35CU+WUJQkZzLG32Xb9oZk7TsBiGuLI+C5ZhdaXFaUwCXLC9G71tmT1QycoOiw1HMn9G
qAuTd7dyZtFl1CRXmvxNxpD6D0Ek8LRHNnze/i09tiF7HH8MIo/dHW9aBkAQgfJ2a4QfMIztFUr1
CWenzfYZ9gVzzbjtI2EEMyykAVnoaHGRK26yyTM2LUTruhQxk/iLX5dMiswbsYU5zsRCOGX+opAk
BjinpP9kvmQEAodWwQpU3bo0FkdhcXlRtw601ZZcA+GOkND9kymPwoGyAEizQOQ0KDXhPZTUngz3
Mur09/A0pmZfuVb3dYalN2tNiB37m3arKKxzlmKRp9vArA1dyAgCTQNBJn5wZIVgApngkZE0VX+b
pdpDreqf5W4ZDQZmDkrm2BvMJvj2NKBLR6miUWA7O1vFiwPN+NGVacaARNwfKT4VPzYZuyDzKu8c
DY4jz5bv+33NkegcYwVvkxsGa/SADq/F3CmT0e4RJWdgibjE0Hs79X1TCSmIiRkYfiFmjFkSSisS
MWrq2aINKDydb8xcWWzKHHgx96weo9U0bqrOE3AiMRehcYOj5ozcF5+YzNbCdEjhwdRi8kQxbQlA
pIhGPyeKm4RDO6MZeI0wCO+2HWBlgB2iFOO8CxZ7Wv07JR9lMK4W1+J0nBqNeDqPDoUWlESMUqCu
PHY8X5UU4JlSB3cI/SOHv6JsjI7wsqY8LLyemp/13frA/sh4SMEkFiV4mNaXQKK033l1fdv1ayvh
PHOfVuKUyjTdAfy5aQDwFcd6fTwjLdbUb7wNEGIcOwMF5gf/DymFJ4JrUv5Ehb3fxuHu41i/KcJB
CF8LMkoJ/tKy+QXWJ+Se1jpDNxeI6psJKyl2IU5Lyceo7PaUbvLeA2spf8wFPeFFE32LhZYHWLQh
pKQnp36rjQoikTUTybyUq9JyifomjncNQb64CbrKztm5YV6nWue/XD0T7+HWn7SWw+GaqBEHta0h
6BL1UrgNPsxxCTfpVeVWR9A7sWSp5XSj6fbgAybQnQrvPG890d/VInf6Z1ZRr/Y2q8Uxj3WJgNjh
GJqq5RcJOrDGCgYs1scq7ivE3yCwsSzq8J8xe6QXV5NBm1Kf6jvruZCUIb5csuI5jIc14sm4zbkG
EhGn1C7MsZ5X85aoBT0go7SJGj09jt3uWS7K8PMudok5876b8Bk7PXwKre0byPnr8MJo5AM7knKk
HHrOJ1Zhykxk0p1NjL8VlbScKuZJuGZi65+jTc1WgDEdcmcgS7AvIn8w1qytFrUL846l1Zn+QVy/
GivuSNFRaYfUhkJafBoSLD832ZfGTkKdeae55qHKTt4dqYkRJiMi4zE8B7TVaJ0E8ySNH9sOnhem
SPzdDEohhQBOG7TvWuvOWaPfzU3yF1bMDfw7Va7PRFoPE0Z4ieBYrysIgBhJAg6to236kvlK+2B9
sghbsM3UDV3VQYI+WGR/g2TmmxgoIN6o6WrZpnIxxDpCX2Hx15F1Z9exOq3dpKEFOvuwO6zqM+5x
UvbvG7HdAOLqGYdjs2dGTKEnDOlWIxPAm+7YvCtwRIVDgRDc2VbRguXWIjqws0b4waf+GD7sFI7S
G2TLwOZt0zl1lCgFBAuS2EOU8ykbZZZ3WfoMrbCCaFPNwpztgOHR4YWkVgIX+MKZKsG4VepmEUSi
OBEJ96bG46Z+m57oZOKrHoKei24d3FhK09iNtrzEJXMwLXIexnS9qLfH/ykiU/iMHutPwuzxvH/M
+qnwdEkVyaPrZiRQlK6HqZuvGGdUwORNAMEPGZhpc8Gz+YNLnjomHqC11/e2dDVfc3FYy7E/jbw2
fjWP4HxQs6UZeLQgFm1+RFkWT0jrGb1MZdMZrOFT/vUmS3QxN+rNT+iqC+8LlP4apTENUH27qinZ
v53w4nwMTSGwyVJLh+utGNqtOt5EGSBm4ygUPoTRLE46W2ETeBykGou3zT8+v8T/8rofUVoboYEM
KVjAFyXa8weZ6mwnhhaf6tC0BYa7QM4fH0qfEyzEct0HGtNInbK3JCYwmSX5epDk4hWnq7oigiuC
UQpdBZVF2I/BkCBv33D47AQgFlEnMuzkS0FBo1YyrhwFie5EM5El5lKPVgN8UohR5n5x3D9Vryje
Lb8QSem9vEjx0FVA6Qo33DCltib3zqaShQMxN0Xy5D0EDLICrk5RTZJ/fhKKDCS0rdq84/C9jI4v
5j95BbI3f2RiQx2sd0O2ebFVRrKolLw5ag3Iijl4AwS7UV2PWtk2OGrWTcf9t6IPX7s7x+r+gncL
iZZGkNb7VG7sMBSEoOKcS3BVlCLO6FLSTXutryVJ6mLmcAaAAjJM2s+IzJwEbi1dy+EMldy85N2Q
5nLbzBoWfMSLqTYnlu/fqtJ1HLl1t9WJzzbQ8PgdymPMKXSkBfGkuXxGNpgTC+9Qm872ZYLOTlnz
x5eWPqs909fIm1gofEfS9RCGy2YPTalaeMcJi5n91qLXbqgcJXshJE0nlBqZVCG3RKlk1Y5GhUCa
NKwnc0GsV20TPGTCY4EW3v9Ezmd5yM/1lT6Q3eyQJFgklZWJ1aKvBEhY+9rWn/j69EtslxFZOhC/
B8RykH4nbgzhrU+xFqLnne1oEr7qyccTWHMpmlLQb9I0RvloDb0gVlSQ2ZbiNlfHV1zyUo4ifauK
UILfGQaJgSLfs0urdmLbG2OHMS310LTa6nq6oDxAolffLj4GKz6hfDJ86oc+9U4Q03Lk6N+l7cZZ
jc8uAgLf9PFIlbofU/jyIc5UKd7EUQIuXPP/nyC/SwNorjKWDgcW9yFcAqDQckNBBKrk2BSn0kbC
OXgx9B2C0XmgQxZK3jq5jm578abfJm9nTEJ3cB86+6kmuXzHMz0OJ21bNcxIk7IlaolqDLSYmaYZ
fO4TJ/AciLEI4qx36W3iV/2tBvhJ5fI+QjYhsDkj4tFuart+3v4TrMIxz9RvnkC7FsJDPGmwSDY6
NGMAeFOPwRP1UPrYmNoXnNoJBNtYPHwtsgR6TI1WVlrO0nHQiQKbuwn3TJvvRdB+cink2PS8vaHV
xYILtTHbLaHxPJ7mb/41eRq13tzcKb7eLewskfqX4oCzUcfYnWQqRCR8hoqYWwgnUKEjIayAS9tI
x8mVMEdhGCmL3i/qvTAFcUfrCSoEZf34s9Ov5poZLSCh/SKXf/+b9vRmbKpaxONL+BUtRAmbQiRw
6yke270B5AjH0rXlBLa+F4ebEMm+svfSYTnXHU7OknGtY5KK0KcQBiR75fLGdtsTOPY2SfaztTEZ
kVdd0bpvOMBJhWuJIuUXUZ2OvurCaSgBx2oubkVoKQed6EvJTfWcW37XUaYNJUxtHL5FCRvBOo7J
5BC0pcTbwEk8FHwYqYZz4XrZ6lR5JI+wUmmDBLBZugibI3uRFj0s9wTkHPFrk32oQUwW9f2E5hte
sJN/8QiXowtRpvuNf6JqXmJMKp3B8AeE6HRNYmGCZglZ/xQiGPlR77+o92crom/A0uwzkgLlL4U0
1BEvVsomvUck26+X7a+gGruwNV1WQuR6+e8lEKQNLIrinKrZ7RgryXjrpLl0P3MSGoSoMnG8TUBR
8KHzRiLELG0d7iGJ4+HdGAGOfTPJapArRhBhTZ6Orsv12FWGVA9OhoEPwtfCbAKNZWar7pM6cuOL
TTG1HvOUjb07qa5NvO1EFe02/J429qwwRiReGiC3dGEviIgB4DIUzmHfpdWveRuXaW1W6Scuo3Ce
hTYE11edFg8w1493OTHEM6OQrUoFl14keEhRGkzXi5p17m7u71aK2w2ML2Wyp1m9Go2m8M0xNN4x
3ErekS/0gr3hT1qne2s7YX8Dv2udIefYzjLOtlYMzZ6+d9Eqgqjo1+Xl0XBQ8kDMB8GHgZ74rRe2
yeMOJtn28zENTGY8ZjwE9fh/OoptzIcOhUWm9u5OUPt8lK8U8joRwfJdSEOPCnjAB61DR6VHgq5N
n6NiXNwks+EtBBF1oF6BaQ+f6b2TMpPWxoLlacjOdOnlIyHYxKCsCfn4VC0A+bGRzG3EItVpCVIa
ikvYvllqxLJCqFpw+bB2Cf8s8xONoiLtKiGRdzrMALWtfxbg1hfHqGzOUC7oF79cxm58Zdq+Xu7Q
9c+CWty5bqaFR+SuroTYh86nJCIiNpq4VOj6assEEAcA0dDGJsM6MebaoZ7czx6TkDd3BZU1cVej
KXGEGXfxb3LIdjkg6SqKKTRxQ2/tlqj+tDVlpXg84qtzrB7MHusMa8vOqdFxP7twIjZJEm05Rhnz
QsSUEuRayLPLbmV8LRd4/u43sZOEtbaQkt78A2e1HapJZa8a+DT4ZQSqV5JuvxI7vIkleQv0pe7K
iM7QV+zOTwQRh89rcpPykeEuPTAWrd2UibUUDcryN6X1lIB6ZgWjtWVorOE3t2H2ZinxPF9hqU7F
tv8MPayHCD9JGNaG+dR5/oTiPA43UwSfwInUsGfmsoGsNVcBDUjlSG0PjGq1FJBfoKpdKUTF2IRM
qdjf9/CQiu0rpzD9i5Qsj1AUbAg3SniiLflLY2nUWKvE9yQhouNUHqZdhCxuA6MNzuB8yFiNg0/x
dT68MUS2qasEQPEk0la6aBOBwbKdmu7J5kQNQsDAOpulWypRlN4b16pD8npEivzF3/RtVioP5/wT
H8zu4cSVZlLan9rUb3pAKxh/m+M3+lawjCS5nAV6VfSEH3TbHRiRvrelvkYo08S7FuKt7b6mQFn4
GYEBP024STc9QgkCT7PpI9KlEJO5D1y+Tuy8TPTbToV/29JyknlEMj9b/fkT84gdhlghXIDCxTef
qmeif7CHKJR+NZE4EDECeIm7uzFpTaN/Dqa2NnUo+oYuUblwrRn9+US0qczIyh3agPFoUelL/uQG
005zMjHqGR71VmePT5jgTE/7BErPMvZkeBD0sut7U+/mG81Hsk3wI1dxpaFininR/XvR5kyAjcdT
kyHJIAw3GQzPpB7gVo6qgv10bcdnB8sXcjnqfwtN/OPlEhe7l+uhWzenOm/5HSRFjbpsIDJ7VkNJ
1KwSxeJbfJ+NxbCMNJrwaJLTKhiHskPUeTEEqyXgRq92KflTWsAXVgZo06TSkTzZVGhJhd8OoSJ5
ex2v9iAB4ArMSnaO7wTz9Td8qezeOyOtRhygH2KQXKPo8eUt7mgrM1x6MjsLMVmMVWgb5qkbPZUz
68jAQ6LPXe5nYuL6bIcgMtXujF0rfpNzPFmNGJpnAm+gJEpvkBx3cWNu8WElvuHGeYdrctxMTKzK
aRS9eTUlCxhjYDedRN1pfu4ffPdOw4gvyWDLY8hpbfVCCYBEYVlADUSt+63eQOvn4o6y97Te6ix/
CWlQLfLQtD8Iudqm5kA35zAQoqZKknjq3r7F+YHlNe08k1Wj4Qw7j58y1Ho7X/MvdYUJz6ObZHFQ
XFBrIX86fyAA7oBbs9MrZH8MimXWGKkR0uP7+pM0Uevhqf73uH375KTmtYW++PZMyho/vhzefEHi
PC7NIpOS7HxMXZrphEEDLtb4R/EY4FUdirWX4xzJjs5cej0x4lwGILZ8ka613TUg8LWrJcr4DG5p
SLT0zBaagqJKfo7ZklayUslNd5WKIPKC9Qr8tvc1sA2PuXy+ll+RFw5KzXQo0RuIJzcNUbmG3u3x
ujwU5WIRyf0INqHfcO3VcsGBUyM0fNg8J9zmqwJxUpqIJdOUfAJhWutQTVhURjFlaWUE9nFVoOS0
ZK4qjh7ijvh9Ak268zEdMDVS00iidHQKVZIZmNd7KvFdRib9Bu0BdXL/JQc5aAm5kkLUUMp3kb7H
rdBnkT4t8K8GIfRorWolU8CJ9eR7CYYeSivEUCfHoBAJJrHVZDn0xZ6C8z15bhQAOcrYPA+TRbIo
N+wYbzDaOHeCMhvjsyzKWHo05os8M21bPi9EWigfkc6/sdxYZ7T7zn2XYXK6p9o95F09Un1pIjwu
RIUnRjz1+yAT+PS1K/cSE8tc6Hbsnz+o4vRQPts13SGowTnaYnwHhR0kw9wO9j8EqZq2Usm9sv+0
qA+PJxSyxVKrpSgQj4p9ZPPG4lPDv7l+MBOR+rh++ZT8fsQJWAQfyoQz/fHP8ICDSsjN8YjuvzRp
j0S3UQ4KT2O6C4AwCGWFDmwyKqW3T9Wo3RNdOeHudN+dgge/j/kRmPw4hVqlDJKwTOXZemp/CIA0
K/8W5h767ZpKwyWZ0VErEXJ/2gUwbcXx/ewVJbDIHeIfbSvYldDveQ4wv4iQIufYToRXP4p4VkWv
QSkMENU5q9jMdO0NwHTF/T9oDT8u2ZpsK3DNmBhAkTpTXml0IhSoqn4di40xQzhSppiuVOfsWNS9
FmrULSIo3eaCrT0AXJahQWti77c7wTUOVUTiZyP5uswhPhQ/0D7cgHuir7nyL3SU65dxFbO2kUvn
aXkJbrj73ef2nrwQOp3c4/LbBri79MXnCpyS+HrY4BPOHFN/gABbKKL2tcUM0zsqt/vgau9LIo8w
bGrHHfb9UfDN9FvchT6IBUWpGv1c3fgNxdt5s2YVcn+lF/5ZLW6O7dwakb2aL20L0GroIc/Kc6Yh
2iGLtBBF0au11NhnRwf+I41jvYbJ3oC48TiypKH7bI4XPVN9iowcwquyetsvJ9dL5G/9TN7z9HxJ
h6DRfWZlbcqyrFPocDlfGxytqTlpw1cFfyhoTR4tWvr1tJ0DZLkwCH+ySOg0Cc8BsZUDehfxgVt7
975a+iM9rKCHLNs0VDni2j9WIyMvwJzOr7PQF1J5SAA2E+e6b51Zg3WJsvpiyrvFWh9sAED3L/8G
gRakducX5jD+xRIKB+gcbOnZmQ8Hvr3B6d/gdL6+OAEX566vCf9MWdl49XwGvXWVgyktuu1onzue
SZsF7IYkVU+1GogFGR+wAXYMQ2eQ/otm4afQtS7m6y6t0HXAuIeVKDg+Bw6CQzsYog4RvwusaIPo
n2+oNb9cwjoJ9aNjSqtYOj/BC/alUpQKTS5YvHfQoFjFLbztyFefRYVA6TrXA4ydcLSeNlKliP5n
a7f9a1n3mPGATOb4XV52VbiY75PBjbXQCTibevExJ+cN/guGS9vR1UJkXqrUeDJL02P0rnWT6OIr
46jnehrcSruaThBdAfhZN4UXza8FmC66C+45Imd0TTbMw+/PfvTvkNmukc8EKlaMI7SSaemiDFJZ
//TIAx6pujAgDBhrLpKJPn7jhEsUTEYZKLxch/Zea88qnb09PBCqUDg2jTnaWs+PG0VdLnL77jCR
tVyKoCYTLFpgGjOzNYNabgTOhSEyT+6JfRXXJR7gQqYUYzradAZHq+vlc0zjEDyE2F/WGogMtcFh
ok3o7xu4wjMhd3h25Awo4X21Dqr174TtQGAxmajh82xGJ+6gh9SmoJLnWfHGzwAAXPCSaSo+8QFp
iQZp2SAg3DbUuQDCvuhiHnPlrPLPkyxe4T7tpCceWHDLOdfN9OziNEt3jMaXEv75lk2kfrmcMLN3
mMpXGenF/FCX2T8TmbpUkbV7Mx4sokkgUgrPY+Tn48BT29eSJcG2BOajxJyYWYxhqVl/R+Y9vksT
HuUbhDSObWW48T8cszNhud15J9gwmMQyUH/xAe2R6wE6d2pmXqU2+2Eidh8ySs15cwCx0as91WqA
/zuwTl9+CmpwueZHUPlqbJ6rWaaXNcY7alFplrQl3cN1ufrtXC9bC260V5gMZMj3+ojB6tTUIIze
uueFgvseGydnZR7wS27cBayUTgT+nK9zP06fiHW0uMl6mXVL167Qm/DYU6N0gD9Ez96qIrknBd+6
K173Bhs2iYkwgnj7onRO/YKFejyWCHc2cgHr60PBL6cQelTA5aerlqrCVUtZwr3aMA1q7fwRR/Aj
LVNwPydYRNrNwXmXUxGO++6NWWhjk1lZKKFeCYVtJj52h8Mc5f2aW/l+t7o8ZsRllVlZlXB/ZH3D
w7ICp3M5iDTC9Adn1SKbHOYPqQ2R9WCxdBIseZryVkmfiXk+cF3r8Y5EDBaljaSWT/driI+5Kl59
ul1kvCbYfenIEGOFxP86AwBPSYD50nfIfq7ZzZvjOj42mZvlAEJuFsA64uNdJeQ/t62GaqOVSN5F
TDQMbTgL1i5jvl43AveNtlzQQlrHWsbByYJiHuUz4Tyj2GiHE2+DxHCtR0vf8xplAHA3CeEF8qd4
4DJql7a/PFRuT7D7Kz2n34rHYN18VZXl9gP9nVs4NpFvN6lnZCRNCtHVVGZFQHU3n/1si050g7GY
d7/Y5f/g8saymNhfkyqIBZO3Lka+FSpP/05/GZ9do4nR5tm6OAgpDaC61fifN0COIxWj5OcE+02f
zvSSwSoBBsxXzotSIRKukU1A7M5w6DfqIdkrkEg0TXNvkDPAq3A6EJ0tpIpFgXIV5yJqSewwgFXQ
fd9wieDUlmZxYOfD3/wSwUn7ZoW2E+HuHvXveP0F4dsTXQQELeMvaxEizrI5Fb2XWmKIdSFN7mvp
njO/JOQZoxszou8h5CZf+EWh7MmckXBt4GMPnZa3rv/tx1nUJ2xVq+V6CA4/G3d4NmkS1QcVyiCf
w70dTwm4DtonEEl1x1UlvWPEHOD1IaL8Ys84DRA+eKq86qDp07q3KLYv7f+rWr9vHQCLGBi9f7WD
faecUjBYFZmJrawriSJdWWHxE5RzkDyFEzyeUW5P39fQETHY1GWjnXeApLgxRkHhQWGaWmR/1FUE
xdt26B0N+fCH8frm979fgTbAicahhKc+wwwzLGqOMo1KnaNQqfni/P6TmDVxluydsUEcohKfwZIu
OCtNCMtG9aO7hsLc044Asj5LARtLRHUWKsPcboUc6b4IE47utE8E1mBzLNL3MhQeS+CN8DyUE9Hk
bglTFqrhpngmqbEg596edVvWi+lZCMa4ruHcuDgv+uGz2OLk2U/e/nzZQkzryTAEUVnrBy9kLN3J
fmmzatOwvEjjO+Eb1W8bAFBGsGlLjnMOYiSRUN92cg3pfjA3AchuzfI0KKg0lJ7fv1ImV5AxC8tz
g2RngS9FUdHTQo2oecBo+BAfdHmcZ8sYYpKNqpdPu/QGd/6eD534XAKsmKEkSu7h0/tb5E0iWPiJ
UsiD9avSRAaDwzVCoaWairNB1Ev86aNK/19tW3XHn43usmsKWn3p7dnR/aWw6c0s8MTmxMmHDPZu
WGkho8xUzWNIVEOZ5/7PPfub4q9/inGYej23jTfRJ4MFygv5pHhWAaVoMuZ6n6W9OLyqF0KGRg2w
VtyYLhxgaEgA4OqNAYsVov62Lb3yoe+Lw7JfePOEGijfdb0j/Ni0QYwsW3Owhvxwkwy0TpgXeFA6
76pczSRgoBj1BItvjETbfrFUCYyk13jDF2i5cgFShHchPGfRs0IecaTMgBIVUwlfkT2FOMV8oBsn
MqGuyhPUGcMKxlE91cqP9+oqGs7qzcZXbRabMNPKCV2iBD0OYPTDYgcPoVN9KXTpFUrmp37kPQWn
QA3X/ZhvJpJ8VBH3qHuSrzkGsPXNxoS01Mk9uKhAvLXpFb/fBsLKqZYcrueryZsjxVR8ZWi582Mo
w5wMYq0u2bz5nZWh/C4TG1B8Wb00i6R0eOgCawpeaLQH1ocFvCOGVK12Z8DeO4O2poGx0P8bPeq3
FiW4i5dJZJv5HKDsGxPEG0EwcB6tYbWxSoSjN6UAuPH3wUeP2JqbmHJVXJos0f8z6XWainTFO+Qt
I8RpNods5gMJWw5kaxWV5bRZie7wbAFl6QkBeE9qrLR+lldEB4G/lbM2vY2XMV2QU2Lpi1GqCvgE
s+w8/guqNtUOICATTXvfZXV3FzxuDw2abgXd5g8FHzZxNuDDAbzLALEFG2uLEzTSEA0jMekpWYMk
IW8yBOSQqGUu2xl3q27HM2r8b4oOd6tsnqv2hhpksztEZBYOamQqtjGX0Sv6vf5uRKD86C1TjyH8
jMaHvHNIqJFy+bUze7kFl3scvHd+TbE4jD6MZyzwiPCOVwhF0v+Y7GA8l7zQPiuRosLxFvyu3vSO
gv41IEGe26bRIkJsYhhVUVzOrPjJP28JE9mtnr8ex5ciHNAHE1imIVMRNCNpnP64TSwv5LWDMXRO
CP+DEHBdbldRtGy95tj0xr44biG5iWNnxSI81eDSLLq+FslYfTStqKbRzzkzJARojIJ92+eAEp8M
g0Dmwi92Wbq08X0owEEMw524pfBUBrdJWhYZOdCftF+5qUnaKB3K3iwliGvv9lMm7ftVGbisl3iz
ssWN2j+uVdx2Iy5Dz1mbYISuMfL6Z0KVvz/rt6r6C05ItwRyuGzmum26Ljp2B6/xr5SbFMGG28Bj
0MWrHrBnUJohEjA36yGGy95l0arlxudXpLYB/lmjNcauP6QHY787hJ3dX62ymMChOOZXtzuMDFTn
daA4iFnMkCiPDGgZ8EAoYGxkpg3lTbRIkIt65yJi9QPT0d8ZefxApUFapYA3r54iWvHXCxIROSs3
Vj7OwSvut/hemCKpn/mvmdpnP5ThD35qtm3tJGOoaZBFgKVAxsI8kSbMymOVbHHnanIurnK/jOgE
rRIubt/XeQkjxuGr1efdUVLIvFgOXVH6pruP6w+2G5dMVXKcCakWmZlg72cj8j+9uglQyyvp5qP5
taFeG41hsV24TrgjdKj/5H9a+uEmhciF/xTK/2LlFRBlBn2YZl6BWC7bbfbf39fgeqjcqkFdM3+G
mIxVyXBzEDia5Y7tdPcIglgy2nLhW33JsvSlDmL0yyHXSHTXxlUcfZ0zgfAC3EkgV4OMQ1JhZOL4
NVvQXrfDvx02ageOKPQ5PbruYH1zguHzvWReG7rduBz50Yrz+S82WzZJEyyrkp3G7l0U2ER4Ckak
QVqqM42XHb4JCtxBwfd8G3JIyE5vFKZOzbq0pvrblh7ZqOG0WSfnrU13o9uZfOHNcao3lIYh9hbY
KtstnYyL4wLi3Y9280fvnICquzIU93SsOvTy96YlnqOzH6EbD3xczW0EUxMEngiCYzqAElhxrwCx
SzyLrIbWhmKiHDjv9xiwKJq6HyZou+flcPnuFrdC/992xoEska0B2xhY423+srR0TrnK93SRXALg
4iMpx5SElcUTQCPvL0bkyzb00JkO8+EJgeT0nw+XZx2fCowPWkwcizg+GrDndJBL2aUv0nNeLcmS
gutBffmYuZWpxhiQcyGL7fON5Wt9sX04qXUY4hSqGzKGpkfJtMQlbHyZtBTE+U4V9ws+Zs5Ayr09
GA126ie46krGTZReHnyn/hpjKqmlJOMPPkXZsDYCeH0Q5V0fwcXpnkXapi4KVI7mlGAHu5p5cBW9
24HBh4ZVq8JU2p8i8TVofiZ0sXP3jYoTqfjELWmHj6bdHjf2Sur4tVBV38tRyhUfQvcgu3oR74Gt
jO69bP86qeNG4c5ZzqgoIzX3hubJL1wKMpxul5yY/6CxFROtRwVaI4Ps7V8W0RD/pC99fjxda/Hx
cZlXmlLx6aJuSF/R+7UqPLr/Cobt+pxjeNWvOaebq3Ymfpdq0kc0r9RXl6AJ8whfa16ffe2N/vZ7
I4rKu76ZuHDHX1RhAi2gh083fHgZdR5ZKWbLMzozbgxkuqRrZm3bcewA8ugu2t0+/DPTEy3E8Bza
cyVB3yLQ+/fhk3z8APofFGVTKhNdfVPCIqUq1fyOl1a9DuOccg8p7qcMuwrMkJeXr4FmmsGLnAUO
zmkxdlCjn/UjSANU8/KdIXGbrbVr1dubnpKn9gkwvraqsRi1yxriJnyWO/eAoTBvPt0uYKrsioBd
oTlLQkU8yTdF+xmndvSWVJCb75SRrKSrT3XkTNKXIQAeQeKe0RtMdlq0REpz5QCQNDcxAk2n5ls3
mD7ugbsMgzb6NWWb7uiPFOCdncyihS6N8KYXAUC14+BnvL6oVBA2zPUvtveMobSHGy7gkIZguboY
ZD0k6B/R1+LjaMFqMPHDDnO+/Bg2NXPbi/xbLoTwyeBRUVw42/zX3mlKBB67xtfh6DhEcnqtoVwv
hAp1UPyw0oTHzIoMZ0ArrpYoKNmvjFumKAusScL1zFzEk9lADsPn9bZfDBV6rK0idE9X6uHzCiL6
SGGMCYXTAnZJpt0hytpf/PpjrxTQFGKUuvx/UpKio8klpVgmcrpdIS5x4D9u5hlfeGufuvCRqYpg
bRmkSAgecGYP8YqDEU0rQ+6MzlmfsyIwRS9BOCGtigcfV+4ZR6IsyF4V7kVxV+ejvRMaWnBKBsd4
XWqxRXjiZ/ky/NFvRBNyX/VrorORBLfb/IiwPGW6QL7VxxTO+zLUj0sdu2mCJcUqh3/d2kuWms7R
Zhgk4hnxoX3G0RCZROD7ezE4FzvgV3tnTqL6ZHi0M93rECFOyeTcIA8mQZ84Y4STl6foYei+AIVy
e7XctojDkXLu+jSdQregs9pUtAHSe9UzrQQ9k6CO1zxJhrIjApvVlpzT9dlJSOHeyZtCDIlMTJlV
gVhzjcxYp4Ys8C9Q6S9iARNNWDfXpd9+KuNPOebRQMt0HmdApVJCgICTWO16MLN6Wb/MEpe+GzAG
+7x3ZdIH1BrLa/rmKvkSqyuRVgtgN0G2LSy8GS7WHl8g9blkRYhMAdqgsK72tXQ9fQNF8if48fal
ZxCtfb7qO4jcrPO0XIgVTVpHgvdMrbqLZ1JKE8zM5mxMYMm/XZ8UYrbYWjOdCahfi/l47TBlYUrT
3e39Tiz2V2UpI9oq/uH7sLIh73ffuhZWdPRSPIGXhKSdL6lLe1mXyZPwTg0RiDyuq/cdJeEtZv+i
sGsyj13iBTQ5y7pCMdRKBqlH3xFRxlQ2PhqFuDQgkN+Zi6lLX05yF1POfDQJHkHyxVl7Fto/cBqc
MGlGlB6GSKmmNt/rdRQmfssHme2tilwnDGkPon6ljlzdV1XA1mgELfLVChEbj1DzS4xCZeN8mPoa
j6zBiWEhOmSgIM0+siXdrNHx4VBDLL6MIsxRb8hq+AOjf0nQ2AoXTzVB+hNGXiCscJLD8BCZ2dc8
S59BMbdvmEhxeKS0oGYe1AKzBUPmqcmV3rahvt/pT6OuZwVP41XccRqwJGkViQsRkfiUjywJF8WT
DIEO+nNWFQ+GJYujN7ULc8RP/G2Fuo1GcRUjL3zyMVDZNYLFFndHllR7rK9FpcrN1QWiwC0NwO0Z
BQAjz2l1oUtE3lpNWJ6L8NSNR2Pk8wrwdbMOTGytsXsOenzcmVIe0MjAusD5u5ETrZULhrDABcUN
QEfdpHYY0g9CC/URIz218vSXR2YQUyQSrZwzRcCxM6C5Qq8r8TtVmkp3EIkvZg3Ovsb7ymeziYJK
2QfQVksxdjpP99930/CMPJ0sonTHiqSHnTgAigx7/hXkQzmRg47s2OAmKsT/UwMvUy0BSNcts1tq
ESYXG3Hdyl5OftwF7QO2Zw2h2E7P7JbZAA4sC7us3EooqBLjUXaY/IX3n5CkMuQEKQuEUoDU0yLy
PL8EI9Sf9GeuMWs1mXymG1dY0ysYaHnrqfc5qXziAVwm9gc/Eu5nmXsv3U/hV6ghye8cwRlgKSMi
kKAroReRagMAQ1l36F2Jlyfkb6Eww32XsH8ms2s4Ln69K5Y/7L02aIy0hjtfJpFWi1Z1hQsc47EO
zwZgCnW/XoTywchGUOEbE6Gt89VW26/31KmHqHjYTHlbv6Pq7qQ+RmzysoGVushb9co28rU8MF5K
b2DvlcS5mUcAGWa/0OJ2Tqw5ebKu4fwR0RSgq97A8dNBbDxJp3/KPdK4JWuF1S0pxPfxxIugAr9Z
/Ryz0XaQYqj4Ul8nHOSDTzgqJOMMrioHstahbOMDlWE5n/GQC8e9XHSfkodSXkPgzIReyM+EIZgv
T0ITUw7hF6dQzR2EDAuG3/cXtoRgu7QlGtKtmCHvH/7rSpHEPblDnZJDJVYxmKwoWLNmS1Dhax1T
Uy70UqYwfbrHqC+8XnhoEWRh7nxq/8pJ92Vkv0C8oLzXcSqWy0INEZOvteFs6tGCX/k5CFYeKPrE
qRBjtVBZMbqm8lyoocJsLQV5okvfyXaT9+xpXUbH7JUCWCgsIj/gTz6P6ryettBswv6XmgbupGF8
sSgLFtbBAk550VHXIr+S4+VW1OGWHwnqGy+ZiDUL4AWiVj2HM3VGaXL4J6MG9lXkcsut5Utxh57k
C83I+qmTZqvYafkPM8djlMWuT4zV9JKFrr7xpu/VAappNbi4gWdzjqTvDrUHN3Yni3V48b2fUUpj
6g+D9iljg5kETGDqiYCVNjunuE8ZsU75HO0wgna2B63Gc5eFf4Tr4Bx9VKmsNEXoBIHP0AkDKbgm
zHzS1Rc7CGC50gVbqjJIN1L1mu/M0pVToOIjlmjDFmbx+f5lv6rO7xilG8ZKnvLNypLOJ978ZMvY
9zdunH0WT92AqX1XQM71C/w/cQevq35boa3OXOmxJ5wSo0sv8bNtR0uZTokSTLlJxSAhH+AWFwdh
hJZO8IJAQhnn8XtVLM39O9OJs0hHFDDB9v3ssS6RCUBdfEC379tkyogWxfeF/kXEknqC82FYbayN
i4puxdk0HuXIQQlvuSuR1o42W6Y0P48Ys7kZMAPwv6JuTnc0HHsDF32doMBTNTmxViYJILj6rZdf
+nYjDsQQs/fGClM/mBxYoXlA7U4sK141mtkq9O/sv9Wlb6H/QPk0akxXBTiOwFGru277+GlWDh41
LOtJ0sndA2VvmQibdhf5/yZhr7go2fHdLKKtsnkV6vZlab7IIXF4+dZ54HnfJL3ea1fWK1lK0z09
U+H+oRZJkBUWnMd3MRRrZ2XPdNs2AY7z/703HewgISIEuMF1YBGwGJU32YP0eoqsPC9g+0zi7E2g
aBckUBtAGxIj03fa8/QvlAbvsxFhss+P6RrzQ6G0aGjzg6Wlk/QlWNCL03bEl/QyPCiJCFviaGPY
/fO/RTCaevU+FMw/LTg8Feucf7uIroeWnCE8Bsjc9/hj1mmK53vPXRZ+eg/LupfFneIFP4dewtww
PY9sZuZF2msHwbnujf5jDqF2Qe4ufnFsDpMYg8/k2W5kjsGC6N6spGxUBTdiTV7R9epaFrwxmb8/
ri8YbIQ//8Q/GpxwEWd74iKOIkjQo4ztSjg8Bdw9Fil3lR3t9t0D0NzUG/nE/eOnoZGe2P/x2WUq
h9IEQvtGOhaCxXePY0I3T1JLIcFUv9FB1IxFDbgBgaxgfCbdVqQ0Fvo6AMyVDAhUKWPtLF4MbOwy
h/NLIYEHjMUXJVYqhGoHNAvvcDAbPjfBc1xLj2Ur45WK0GoAONZsDBcpfX2bqexgEAqvHWqCw0AJ
ZRfNYxvHIZ5ft5ablOJYLonBlcWmfGf0XDeYVndd5ofHlZe38GGVR7WAekMrllcbbKkAUuTl205y
V55kopJyjuXbbALmCM+Ch7VXBAIQrlwcWjZYsoeKbbE3TCs5OzHHSJIfWdQ/7HpTZbdTUy+HTSMv
vFEjKJkzZnNtATiLePDjLMpzdnbcGRhalWsaXFvBW5PiRyB0kohhJn6hzD/ko4c6LsbmkbQUcew4
5yN1faZeDautzLhzbh3kR6Eq00bAzpVic4KLjhf3eAf61A3YfLLJVa88CWvTWGUewQXzff+VYvqn
QjRmL+LjCaoX/ixbZUkPIdlhEON4xO/lDBAxylqeVyxoyTHVsu7OJdqDZyZja7dvEzsODqhAdoJQ
vbUkMqf8ZoPDfOhpO6mPGiyGc9679Ss/MFWHYn97vKW7k5EGmWmTGH8wsuUHDJxS28bTCzDCu82f
1FyPH18ctB1ndMrMxd/2KtoHDdvh5KBcnQAKXCMW2WXl29KhMJ7saeqpVLP+sQNY5WgAde5EtqqT
QrlSIMSmV8x5hHj7MQM4aey0bPNb8ZhRwatzdrgktjM+xP/rvrV9psHAw+mhaPnng+qnDZ6vR0XT
RT/yim0MyGAhzKgCRr6D5RUm1G9A2alC0gOtZTKN5hW19k1fo6A8tCZ7miqKq0XprfR6W+lqXkbU
PB1EC8g5Ls6FLREQtkit5v5hH8AJpaLRu7h3LRFn68hS1EWFA4I1k5O26lqyFom3oHmgHZbzQRBg
tRgqJC/l+xa2cqL2eKnyPRFK2WYwgaPRYsVSoY7t+GQLFik2U5OzUnBcHXUcqwf/md0JSilGClvY
nHHbgF/LWNbBv05mGsJXDG2GT/innK0oC7ZPaCmXoB+QEmJUtqQUt0PvbnSKMi4/DqAg9PtZp1H7
qW3zvm9F1zi3+JkvPA3Adj68bCGL1fWWxOML6F4ePI3DdM0vr2KvwqFO9NlrEJ5nIbqf5ZyxFPsp
lMl2hkEDkhicdL95phael1wp6mVYgZmYfuSpTJISetUKH9Txq8U633CQihfMM1WZvFH9IJNEKI8M
ahql7VR+mJZPQz6iL4wHT7kxspkHbL8x+2zhMNu0xpMn9W3Od+ZKAy1RXXZinVUygrnk2cDp+sGZ
+D+rtpqaj8kxnnMmqrhqXsMCUwvKNDqA9J37ZEZIGfpxlUth3psEee/uDozUdm8rGiw9i4o89avz
1RnWt9wi9M9OORipBHe415v1t9+xHF176B/iQY0gse2L1ZqO2MYQMtxZVm/qdYSdIsUv1XuL3noO
O1yljnuX835yUmudsoqdIhMpaDGeSdEQ1JeXEILGjmrdu8cLWC1va9t09Jo7hCIqUuhe6oHbkHQN
2ibCnCUdUPEhOnEJRhv0bLeZ01BTUFdlXlzLaoAtpQdUSps8ib5E1c/HGP73YChMo1fp0YzRJw/U
+Pv5fVhIJuklF+jgjwYxlOPUuYtQxr9zvf43HEx5z6Le7/XPOWjYYQWIl7k6X8EI/uBICTgJ4IA/
+dBikvlSchI0fHUYgwTBT1j4X0lk85/mkwC6tD4Pq7B/Hx+BJjXX8p3NijUQSdEJXZNWPeIaLHo9
MgximQC6qQ2sNEkqqH4jzR9Smycz8FFR4QoCBvJfO58ZvXIq1DX2JkxiNeSVhChvC/vBYJDycgjb
4iHyqwT1oD42rh5FxG98e2jo40tqBmCaGsSzcKnHk1WaVy3aTbH4Y34g4EgUQ4SCmcSk7gws8kRE
j9/Kdi7KzZpolfpwiy/+sVeKK4N6CizT+dvBwLMg9apHtTVgQ4pKfLEFkHRtVx5QJ5/Q/Pd2/EfZ
KKLcitTxdr71D3Q2904lL85SNQVNxNGwsfmvYUXtVMn/eUvhqDj3COX+td76cKD86uZQTU+Ek+es
z8koBMl/QuSKcXg6N+/haiJRpW6JGJZXXccpv1ozJuwY+XYYCtpl7Xbm9FcpJbX2uJc4XKEU+gbq
VvGTrLrrLbZlAkmxQ5IQrF5EZ/XvlH3qOdqrh9tiX/mDkmFjmYxPBhG5uZlUO3fZGCUb/+pfRKbm
KF9QgygcGlorvbILfhbiNRjJMDhlVMC4v+JVfU3tuxHoFQVn0G7F6Y0cPPJfHhjGb7AGT/HHbMOZ
gaoNwT0I7DKbUun6c7Jry12LpixRIkrjczO8P5RH37O9kRn9J4dgxMQx01tcz7FQuygzfchL2FcH
g6RuGabcEdgO/tGIKr6+c2Bo2gNhouXDcfabqAGF1I3rTUBjBBhXMG8CfnrJVqeIyujKTBPI5gk3
tt0H0Y1grS/U3RaGJRhLXFe70JhBCkZ99JueAyIzlNIQ3YI3xODUpvNcaKDgImHNSLimc3eP0aDc
2IORqaFWHC6lB5ilZDIFZx9I1Q3ycK6KOzPk/wtIxue8uwo1YGCZSzzufMueDEXofJVHzyAIOUVq
rt5sRFGGRCBCh5Y6CoofwTSS771beQdsH3VOIyZVKjpXV6zquOfVpO+EOB3XLoEvUGivw8nL4rjv
VKmjiRCGPZ7Lxs/QMI7xhnh2iOc43+m96DmLUuV9jOBurWq4s8Mb+aPw9vLQJgQR2bt954LaNv39
TkB3OsyEPB/wsaE9VWvzF7IUAGKvaGIQI67g/+/pQF2EpSlakzIeYfT4Wc1gCbZge2FCzgpMMn0N
gzYd/7i9XLVNgItyfSh9veRH85jfatLYolKd90N1wG22oToDOK2xPV3fXV1EPQa3MwyEzrTzASZP
OyzFC68aBc/RfWE8NOUYB6f9e7jqv8cZJRVuW7S2B2fc47xT+BvjYro3FBaWm5PBgjO3h1yL+oRt
FYzEsiYbRi4Mmraphz/aKlha4rVC9kuhR8XVULyOAYxXJPLBIHrhz6Z0LltOdKTOeNO1uy3RNjE4
5LT2+tVZlCpcfrCZwG0AX80U5xP7RtyImGLzMEm5vcZ1uyqsOpzZRBPo5btxchRqnIeyDvO2WTkb
GOTlPBnWEdYA2RYD1ZhLCQmg0v8taD/Pc58YtJ10Lyt1aqTWeUjyRhQKg3gzi32FkGwceULygzmw
3SzzHm8tLaIGSkkBX6j4wuxOAd22WGiciP/rF/FFmL6GVC8M7zdsaKV1kwKeEjTXQsGD6XNe9ZqE
QBag26cPZXCnHPObrwOql5DOW7SDtAmR+oEeD+TGNT4RzUhYubgk/McmVVBJjksKYCkKuL48W0qE
4+6XOx/6rCgMhybmG9zLW4X2M2YqsVLy4pcoR5kGQRjoGKSxUDz7RaB+vpM6Jj9bhpmlLKR79DDB
IX1xwMKw7Q7ty6NFBj4I60nUoB4VFx3JhDtkdKpVqhZFwCCqsYshxZtnfA9qzpgBFE1/Y0fJjzoA
zyCZLBrg7sgGFSynMDP2uPPQa4lQ2rXCcq7N1ZFrjQ8NmXjLD6LrAZpawn5ri5VxAIjjno4XBxWl
Q6NyRA5Fr+oeRwVWZrGJS2qH3CfIfilvPqXMLYkxFn+32QKxjJt92WnONj28HIqk0b9ER8IYxcih
WDaLM1sWAscUoEVskTaItoxJ27E5kFbua6Ji9V8k6zSlUPj1OCHfvpoWjPfOjW8Lhik2CFgFRpux
Y9bjiSA0iet0Qti2zUtBgJXTQdLEBpZoPY1X0SWBpVQOI4KILhxYx1hiedIS3ir5rI4EIPRpyYd+
ySq4Y4TfDiYW8jbVyFzibe7kemoPRoPY+KGvu1d5i+BOvqGS+jINkVrRDQf/njDvPDNLFV40tK3C
rO70I3RcW9l/2/2vrHFuiGZo3GnFhY6RSXk0aBGoma7vsQEgo1rLvVjqzCFHpP2flkM27Xuu0mgc
KEenGs9sAjXlDtxTguC04m/8S1in8u63xOvcSB0mepXmYeHskCDlhEWxqiEVrfZrO2E7e7R5LZfG
KwrPOzw9yWfXQt3OCd8ljh7Dszm10NAOSrf55ffADrOT4miyDjD8680EGxN4MO2vqHHiS6nj6Wqu
eKbOvdBzoI9v+8DdHf4KfoCTE98gnDqyjls8r+JoZwZxZv9TwdPtInCFO+PfC7jIk1ifyQC/Y5hH
OPIWJ/l55moDdbRtWT4wevWJXEIHhRpvWZ4g0E0+J0ys023QCebdHuA/ioXKNgkV59T6Ng2F5zsh
Mampsohmmf9XqctMivGIi1oJ5gaZKRuuAoz8jhLHNUvorivX3g2usvLQncwldWQm4gg69wdaLk6N
mOK5fA9qIeERhKGLyyt2lNrdfWIHMy2v4PkNolVjOw/7tMZU4RYbAPA6JfM2EjQaq6Mq5yj6OABH
4g59WvUzM+Fpkna/KabX+UnRxsA3CgG9tCYhQkzxJUmwgXcnd9WTZSvzLVXqtE7NVKptyXx1vQVx
P8fAm7K2XNQLptl2lk2MfjMbh24AuiwvXJgY5nz/FMllH5qmvFnoqZm269bDAAPZ235/wUQmHcCT
HNtcaMKlAyJRj8/FLL/GzuAbUWG4E2tY7CVBp3/HDrdHbOwxv6DWPbNdgX2ajbWtt3FHIgyv30dc
kxo2vM07uhAt76xJ9pggodeGgZ5KtRL6jHyypHcPj+KH8efoCAWhZEiIpcqRa+RQ6t3CAiCf94qq
0B+7Cx/6YBgsKDU+WD6/6TuEsZovvD3rhQ9UEDso6K3DgGSOFOCqjAivlVsV48kSbzEjiO6DhS9i
+q/G7GxJYjkVDekUEMnJZjuuU1g4Cx8S75zJ1A9sOLS5Q48Tzy/ytXk1ELciVE4YUVw+gvvbQTqv
tz/BG/Ra/BMlf6I8hm7pWqryjYvadF5KvCELPhEosyxe2ZiZOF+489ENZ6qJKudxteMvwGsXw68b
w/Qct7LxcU/j4DYtidwQVsFcjPX06yBntt4NQa2nnPnytD3HD/PeUoLKvx9gY/EwK7tWzXGn+6vt
TcZuDvYR4vLhkHjUwi5O+5uPreQFrMrUR7w13DGE2c5og7Sr0LJuM4PrVj2Hq86+kxd6Paby41jR
utW+PnWuXmL4pMK1Nmc5DCL8FudZX/1uBAYf4Nmd9MY8RCXc3gjPjQhPEzAMMDJvzn7i7QJW9trM
gsbklf0A09JKaYwWySS7cHxwZQdVX9xSTCr2EgJS0HUoajomnvGU+agZWU6BXlNegRfYFFvcPRH8
gzzjPdimzG9NE8tS+tASJ3x8jalhw1K40gYHDLa10nmmwhDSn81sdOpBGvkJ9DGt6ckBLw7c9q5w
Mw4BUyKSi2XeNZlG9Q5q+7ZpqEZwMMu3XuOVWaM09WPRqXezXrdJx/hENP7gsgD3MNZTf3n8PZuf
q1y9dEWykffDqRQTxuEeRhp2lzfOZ5itiqOycCsStXaqYjSZ9Q1VsrZDrs8kID3lFIS7eaL8or5M
kmAN6T1Xw0qzyMm/kjCmHkNv7WjHhPHbCa0wgVUB0mqcAETDVMdTuLAKS3+qkA1+9iQGDCpLEb5+
QGqxI3MeNNFG9K/Uz2D7BvD3V9kYTjW/PHd5LOtHzr3SYFPh3gLEmN/UzRCoIRRpmOWxiSKtjqZV
1Tl3eDCIvDVZpL8iVHdfTk6mgAve//AL01jJ9PahwTHDaUNfTZIbRDz2GyKUeOQRk0F1THDTxv9y
hK+xRox8fzxRvnagkP6h+zGuLBjyWMcEdiXw0fprIDIAXfkB3RD7lsGY665/vt7xhYBdFUh18s5p
e9bj8Hb6Kp8sNv26bRhFYCMzDeEFhTLVRU8Z/3EEh9DB+BW/pkvLpDMeB0B1bb62P7U1aMciGKn0
C7QRhJXcyHGozwwLRSlPZcrUQGPYOPrD1yge/IgxfGJSFQ68J1aOeKvj5FowJV28PGA+2nI2tD93
t1ZpVYEKzzMuMcwIiNrhzdiL4YXYt1OTYrGOahzffcike/w6qwYtpccF1TM+udLsvILDsRWtIxYm
CeehTAkHUvB91zZinByYhIy0kzDKyyBRXlQxFA3jsCvejYHHhqJXSexR+w7qtSi7xK3hka1ojMlo
gz0XIww+pq7XC2nM64WYXPf2YHD2JrMuUJaH73THKP+OGTvPc4zdDTiRGFwR4INFeJTRmCEn/CZR
KX08G7Xc0aPGvwR+Na222LAXXUuYvwH63CZbKPctH3snv5YRdq2sUZnClM6t5U/zXO71bjbLgdTf
vWe4l98gIhtRtHd7fdPv7JGdnqNpku7Av62xicjYrQSfiHPjlJrxgphi4iWthn/Ek179AScSwdUd
bvIBAgEkNLH3q1uQLyMGT90FspLfPSiGblHdBexol/U1iy7Odi0rklsq0JHypTt07P+PsmHhBjfZ
m546Fdj1uvV/MnZvUzMhl/eFkCKGLLrVzEpbosW6qs7k0TNEoK9XujjWfdQ/RCjrr/8LSliu5goI
d8HGNLqF8lS4rm5l1vnWjaYzu4hzKLlbUyRPnwjz4Al2jYYMCKlBn6Cyy3sANBTezCs0Y6vl+vW3
x6WrulIL1m5+oWGdkE8Slsrfb16KiNvI/CkXclvz5IbBUkMV/IWviZJlppoohJARoM31F+oJzkzC
DZxrsjXQ8X1dISTeF9yR7F+cjegVvbcGXs9MoIeicjvK925d4ijWjJ+y5u05nByrc/Om/HprWjSX
sydv+02CXZsbtKnhFFc3kuoHAKi8fU3qCtd5jDgClH+MAzsYetslmBx5bchCb7r5ITGGXGnw7WNu
wj/bUQRA731sULHTaZrdf+0a1iz+79QvJabje6gUmQUXUM0CEFRW2AhbgWw2pmOFmhFHkHn8+HHd
NYRHQZ1Fl/NlaXz/9Ftz166i/fzM28I5NgFiGU3Zl5Jm60UmhSOb1AUnISuRxeg1aDiTSDJsVftY
n8pZMXwjrArMx6EnxNwXLTPmWjBbrQ/9DKi2VgTpRpLGpcgiAxrOUHRicarhEI66YYXmyEaeFtOK
WfQ6FcFczM40ngJhDbXMKjQtRhgHT35MO5CPmugs1sLoOZjfSPc1XpahqRaij/O1V7pUxre9Mpf0
OinNRzHVA4Pg8Kxy8TK6Ud4JHuuCGlRWPIJVkb1f4pulLlrKeyGhSEgd821KlWn7wVFZsZuMgNDI
NkALxlLtMfPic/dEUpwf+ZNkL8JuNx28eFtAe5d2Lv6UsMJvpI9qKvt47DBfs467wE/40d+eGqvo
uoGJPcU/Q+7aR6tt3w/MKSBSZQ/QigNn0BC1QCxYeZXN0dKHZPXUJybMY1TLb2U7sdzOFpzNcssV
GJ1NMTfF4JFzZC6KmoZQ1QjBFv0/G9Wi086mAi7jezwsl1YNPq4nzdSkklKY2kcQRfmlAnzWnXBe
MTL1GCJqvSwv54VUbx2npEnOAqtj/U/Z/ucHBv4FUpcEPw3+/0P2g9nTB60++WgW7CA0BGaSGjvg
9zDPETj28WNf34y1+DqQoNrUcPvQt9I1gPjSRZhZehBHIOmCr5AuHIV/kYdW0V/JRtzMYg+0V/Up
kW49FbXM9YF2TSEkJQ7Z6kLyDs3s5A/j0aKiniMijBoqdzAl1bZ6eBXl2x7ERXEn05qkVTcYGWRX
SB1a+PdNA+YYlK95jAnVFZk6Zg7ZEqC9BZVyW7wyWnFKNNLnwmiuIhhTkOKRu1geH3NOIAiG6Zzd
lN2eVe0mpo4sGgLuAr2bENe3f70fVu2umtni9a/3WNqz2GjJVal4/rskQdqvQTNdRyxAgaWE7Qdi
VfCJU7feMTrLkQLZ4MiwZtJd2E4yYDfvT7PTZq6sOfoEy9B05Gvk76RfYIMFDymtlMvsRZcYhEOn
WkcKvWMkj1SaIxVT1sI9F8Yfl413EbXN8Kekw+eiTg/aKCGUiC6DasN5guFr27f7vJYKka8PaLpc
H+4vRl2a3qiIrii+7TbKMJDHpaTlNmixO+Q0geyJMo40if8xWgdDMZ6yVbHTVEXvRO7zpGZ8k3Us
lQz3tMLEUkdttlk8HO31FKGIf2QzW6lQaiwxqHLsvpXCmf7O2yumpmbFScMaCpVMsnKN0Rk+FcLo
jbf7ZHAlutS9kOz4AaIF1Vew6Qt/LjHbVXOLsTAmsdUsAgekNjbFEZHiHTFf5vPd9xlEVLiOXl7+
e2gndpDNW3kfgDiTC7hfvX09JUBVJkEYcYz/rZbQmrQwEAF8hfsUGREQvBrusaMa7EQvJao9qU5Q
PmUu/uBe52Xt0Fk06uIgwpWAHhYaey8xRlaTOgmYZGBlnNREU6Lf7nd9nveODG59Xq31rdCg5wBM
zWOHTrfFnZStjulnUSPyVljazRYSpDrZ4PDiCrnEvp6Uv31iGCWw29laAZ6ipRWp2bY9wghwWNqL
Z6qdja1YRiM6UOqktTiIAJXPET7VAEBqIoU26ZkFJYE/8Qr+BuO8gxgtFbYbdT4vzMhUewfSgDuq
QOHWkKTOXd2p+/Qc6XjPYcNdvuKmO66W+aEuw7G6/W8CGFQINSG54I5bCJq+NynWO5Cd+CsAcYPr
RJ/KuAATl/MaOMYbattym00et6ry/zTP9zaxTP/gTbioa91V7F9VbJqKPAjJxLXT7AnuuyZTyxHd
miwhPZ8EqOpfkJf6IIeOhAtkL2/NPrfwq5gW+MGWsTUSF9GrzZH7QDBusjtfyJb2ZDpK9Ivyli+Y
apIlkQzqzwg1rlqluHKycdqUST2BS+o2cdDeak8sJu1AIk8t+3Np2aVObrSXVU67S2q7JeQJV6U1
u2QARuEyufgLFY9Jl6Yy986/zJAVnW48Fuz7eiykoi6RoA3zzpp84IIRWTo+w8I1HcN9EN6Kkm6Z
DGcXGYImusSBc8uqpJ0E9/XWjo14wcMzXfYHJnVDAxHPQ3x9j3CU/7vMTRsaZyeH4nh4dbcMj45Z
rXPO7N/xYHPlOvq/QhykdvHC8dh54QJ68vlGcryO2yrH5Bvh9gOdOzZyvcSX7Csjr4GETy5oJb0P
ZHMlwuLDNTyKikNnMPVtcbCI6h+b0H1SxjA1/pRXJlK6PQ3tVvwhxP8qxOinqmqlTXAE8TmMH3M/
dFiPslgZ0JjTMCdg8x5Py0gTwmfSIXUXP8dISoXeuoMZnvFzBY+c9ynYK6l2ht4BxFe7bxTyC3pm
Q3Qns0RorhkmJ5NbtNVdLUPhc7Arpt0sWKKKiniou623SefwRqdiHTX7a1CwSI3BlQYJXaSO2S6N
gz8cOt56iuUWkPhM2ZrZ3kufBhTqXJS5tl0Utr0EgOArETFkatuEWY/1i9POrq1O+sEj5U7MrozY
zTl4CmJvmJUsuelhbw3/lcykrb4TRsGRPhGiGrt4PzQx8yve09ctRDwe7NMMrm6FWvYFttw/Hany
s7yuobPE9vuLnZokI1zkKOckc3hbLygAsjfYH/Mv2gzgEVQKvcyfMQQMx0bWFIRFT8eeU4YM5DV/
kIylEWpKhs1ctxdLtjITQqZHMOee8m5pVyBcOT20SQkQg91kiyLAvpkiliIjYWnYLuuMhauEVRrz
a2y2AFRLtn6g7+S7eFSE8MbZ4C5ORQ9L/UUu77eFHVnfDQdFWbPjlz8w1apNJ/33VtrCIT+z3l+m
67nZpn6oTRMx5Tv/6YWgmND/lXD2OUeTdEKVlhHVfgGKukCX3ZZ/IrIe4PLAsssENa3Kvtz/IzCR
Luo30wq54lChx9Irsht7z9RxLIOC0IXdtp+GrbFnvs4NGzI4YLq5B39NrQL7M6wmTTLHPwIKLOq7
/K6WAxSL2kGQnFo62ZzQqAJ02yJacMZ/kGM/KYVDwhGRYmFHEnif8KiMlyxvCdce15pnqGoPhN65
KUkDCWzZB+mtqjbXjAkD8nWi9jSNZ7lyuiuHdi9kPnRjC2ZM8gFHQTP4IS6OEqTMfJjKCjZDQQo8
cmveykGF3BX2U6IXcgFhtwIoyITNUT9utLQkr6I/DSiB4xPQBEmA2WPoMSWRDynmsBeh9ghvouCS
rYUVggE/+8MOmEhl8W4eiE13HZJ5R3wRngnWHLaURtY8EYU80TyM93LF4jvMJ9FMj/7lMs8MTFf5
RfzSAMBJTwYt37FVn0gY/kdstbCoft/jvRDnerRxDLq3SCCz0Pypx7g6T2T4TMqzPr9mFjOh7VMY
I64dBcNy0+ZmozrfMYZZ3y3DjoG6chJ2ZnzfnlSTfI+AjXN+BekUgj/MRJjYnJtc8DfjNfS5HAX9
KwUKDKRqghYbs6BCURfX4YJUeFjH4wnPZvu1Yp10lmtHWPAkh86HUiuv4quszaLCPmmzX/3pzJve
M3CdjMvPEA3prA9axb05anyGc+2M3LPgX5jkuSAXa3rvHu46lxFAFJhTAuVgx3LWmpNrQYYQRO4g
QAEcaezeZqX9gmFY8ZVvavqi7LfjDeWH2OeyA4N6AEKeb4VDvHjKz/ut7acU2ZkHcFaKJ81u64ur
PF6ZAVafWPOLBxV5uCGT+xTjRFnX/7yFSc6PIwfvZJwyVyy5Qi8hrqYcN2wADjZzSU5owB1tKwYQ
0aRxiNKEYIAHVP/rHYvaGKDbQiSsFuEa322YuLTdfkYZ0579NR9VxFnhMvBD2lkDOhGEPam2zmae
vsa7DSLvv6n7BoDXOAKoxHu2NVZyu9wsb2xVEX2FWiNaaCnkBEp5hHVy+WcPdKGrSkcb9GEhF82h
NJgvdtuQpZsuR2SPpuBkEOwXI3yk0fCilEG6Oxfb3juQB6fl1sEn0gGQ5zvv1v9jAGCnzu9mRDFJ
PdXwk4YsVuZVoU+gM61QU1wsy5RpPcN6toI7+1cqI3GOdcXcY0axF/t0CA8O5gaoUGjLZlUQPnd8
Qgzm6MBRZXuN4U3g1adTlRIiUzQU9hgQMi0cMIhVviloeArIAkUeCvyqssNHhTZD+JqFLOPQGAGB
zBFtMoVSKDiwqQqBm24LMm91oE43TvuKrKKIsr1UtAu35MVNeDsumBZESAnwZoCaGLnaS1pEiYR4
kVIWPoDQARY7xCuCUDbbly6jTopbxAz8aU5rkMqPCTTOhMF32Xn0/bucvqxNNueTOMUVR64MIMIC
D6Dz0urdrrvGFyiNzG5N0gnAZqqhZII5Nd+Skyof0dhr4Uxj5/j2ijaA/aI4FdoF1yAAUSfZxlEn
5zIPFGWgo+Te5HIVTMVtOYqxeyd6Ke+bLiTiDlUIFf5axE6isPj2B1l/4Z5x5CnuVBQLsZMsNMGP
sPTnVE1w7mtS8gHcB3YqyfdZUQJ+7plzj4BzVyC0wFGrYrfmpkOTnzE524CvIWUwzX6jPY5429m0
it6ySo6hnkdrNuhtGhzeH6DorHBg+c1joWofHuH8ihUbfwxJTkRO0sKTb2+7JPwheJB/iLawKv0K
A8ssBSVLn2noy3kNLHfKbcynqEqQW6xmVD8BdUkH4a+qoR3UJXn0AGOR5BnO4ozdPTynOZPsvXvn
PDSC879SiSCRUXajeuffOn2852SDpS94f2KdG/Op+UnP39mE1dWQvGfl87bFCQPp3rWt4AfaDCsA
yh7/pxzE4Zfa7i/k5K/Rddl5vHd1/lWoIkqO4mTS5Y6eAOgN04Ga1XHD6Y5SZsvatOp4ju4a/+Uu
bX9mVaB4v5DUOENaMmT1wOmWYr0/dCbfLsUotd0bB+y8izGHayFhmhIxPWtdVMok1ff6KzADSxal
uUvOMkt0vrEJq5vjt7RY8vcDxou0KxnFXewKdihrD8hJdhGkqaNzv5Rh4y9yegTk/78BjxuH8tEy
mXQfVTOo0+9InRyv11EtkGC42l2zJR0Ll6/yGGPl4d/Zvxh96XVEpQTsFKWEPpz1tfqpnjhpqf8t
sqgbHdP8F+iXzkzOo+nkI9WsVxRiDTdpj12b3sW7dBWwsD339TdJj66YBIG/akKDI0nxXFR5CxEo
ILa7twkZ08oBXCynNm1rhj0SAvSfCXBJZ5IDom7kUwCADXCeo/De8nuyQERGzdGyPIrCAEwbi/2L
GivvYKFQKiZzywj0xI2N0XRHE2F62fY5rpg3WjULZL54OKSm3LjTXenjPxsoQodp/ARQ7wka5weE
eKP4pmTjRYuazTTzbtaYbNn3AoOicWvPdgrwYp02QOqv4my48FO6fXIF1eKTN2gt9pTzflJfCfAZ
cLcPGotifBW/ANlkk84AvKHEy0dZx9UTo3nvVNnnFHPGJwtcPQMnAPhpNSMilUUTfou/53gKn5nV
HhEGSwqeJ5Eo1T/fK3Mi4aTbHRCV4vmW7juazWsCMcgL1HQcPV4jY95W7GmgaxDvTr1575LQnFpb
owTTkCkbadPIMybJG+qSQMY6s0pTc4sip9DXqQ5I/N9yahhUYkf42YXgEW/lMETO5Mn/sZqeCKC7
F/F+gZuEEUUhTUlxAEp3XaRb2nN8vrDn3EzPdB0JspMdOpkePiW6HRbhyjmZJ4jLm5gLF4FbOpp9
jFBYVLZ/4hPfiDJcUi1Vxfs0IXZ/aLQJ4cba6VY50Cg147+BAGcUwUyZ3Ky7U6tbAU7N9g/+da14
eOelPIE23yXvYl3PpzRClNzq4emfHMDirXboV323J5f9XCJlX5Ag/jBkJYCiXc9tj0wut80i+GmK
CkaegEmf5IkfjmI809dJp94EzdMoJJjF0DMB888EaHHHBpo9N1h3HbevkgyVAdkl7XzH2wNMlXHc
Y8ks1tBYTY0yHqntZXeqWI49J27zVUvXMJeh8phRO2HMMbdhhJ4jcxITroEFhHsEUVeyVoeao1pj
qJxOT3JjSomqpSgDaVMzMCxKEAF2BcUdFZrmPbilCV4Zq3cFYMqpZHr1MOw6tqmWGCHgwkzTeRQZ
WuNdnM5kvheFh5Fpbq2vauA6axbMcwjU4S/kst5pCra9ES9zZjUwQH+teZ5n6EcBG7vN7kKAKKAs
8Ev/ZEdbG8bFwyqPYGkMSlWlKqgXk8wFxrE2Bk38sGEB/VufVFEVEXL1EcE8Km6jXvcUSBKnyX1t
0WO+9g/MszfkC0HEMm3fgVcb4VBRTFmEjLe3+MtXGiJtmemX6rARIKcl2WQZnfMoxJ1+/5EVjiJC
48VjRvI8gTmpT2EVTpiSRON/D7ATScVrurHbb0k0tlRRbserGM3FWscitDcKJuOn7ziC9tX4uhAd
E4OLFw/IC3lF2bO75yeK7o5TlE+n9QJex/g8Pv2NkKhprWebYN3jW/we/T5QgXfBf7y4scJRltH/
zG8K9aO+4iM1iaBLXTFde/c1d7q8ud/CVMlNURXfG9r4YiU7+kIlioPuNiwxovAxijxSvmQ+GD/6
XUwueXc/r7cuvjs2CwKpeDyH5WoJ2cwUHnvkZd3hm/ugHr8Aw4sigB+bE7xX6ZSBSx7m0kTk2Z0i
eAFwWzsDPbD+mXih3U1leCBomb3EtnZcs3Z7GHjKrgK2m2XSjvMNqtJwhvF0lKs8AXO72qJxp5FD
Gzv6JYO1q7k4rRg3F/+7qUKhT2p5PNZ1U3fUmBBxhbziT978NzrxdUfmOgBo8ZFEcyiMRR1Jl2+J
Wg3iVSRX3RnW8zmFbm5Ex7UOgZplj5YNZHa6kLZPd+yZ3BF/kt0XFftL5dT1jQMBT+dCYyJpF/TE
pX8Bm4r/+XBIn6xW75k5MUXqvqsCCDP8feZq3kY85YzaxN8oHLAMLSXE26VLNBLiAEnzXi/vllQL
Po9QRg46ZOjDFWHz6wU8gvgWCpiLEEULpT71GMORP/jtvJd5ZEuSoAGmykf73Fw78/U6M754tNCi
6ILDq8b9HXmFsruCyrGWErrPv2Z18xhwZ/7jStesSO7vjsdRwoMMJZdaTv3s5TiqGWXX4uUCiipR
1yFm049Yv+BoaIf6qA13v1g86oHKEwJBvam31hxC+S+i7ItpK5qFDRf7SF3GULYDrwa4MVptm7WU
eUM6O56Xw2Y8fgWjyq50I2wljP6mgdKr+k9YSs6UON3zeqA/9ymBEO65axaWbQ4r4okvygLdbvwc
qglaUYlluLBK1ckBfphz1SzRxJY1Alja+zHM1RIy/1Y7GgMUUfHIsZUzKn0t5UdpBmn66zD+L4M1
g0a8pDvDBMt/VmW+Mbn3d9XcK9GcY9H4+1pEeBSb1XVebFrOeb4lZ05tRUw5YtjIDCNhzxpc+O7A
GOEaeaxM/xqZWtyPycNQClzUDs4e9UhJxlDa/sdtza7EMU3rkfhCL3i5sizumqqtyrbpMbodh3oG
F3lIbzWUx4JYUUByGxKSWzxariI++nP2ID7tMnCQS1Qu/tI9OO9cXADDRpOqL6YV9pejeJy8gCyx
YAkqTZJ+oykXOl9IgzfzQh5QkBHsjb0Sa9PzlvFlPxel+V1+6BuR+O4bWunL0X4QtLDAo2lWDDOD
HLMdhT3Bcjr5gn5yM0lrnyTZeMMOe1NYIBDNSPcLbhveplmG52Tk+3/7iZot502D+EBTi25I0yJK
Jid52qJyDfZ/6GHh8Fa8uzk0NohYdrCDhjX220HHQZleX/Egd1nDLNBCUk5Ofjr8g0MxbGbjSeew
EuO2g5rvYpAoC13heNGkxjcRsUGxNsf57IR0JPTetIUgEkUDzyCxM8Tpu1Nrw3r/lsgkZ/UcPY2Y
1uSK/ErA9w26/Q286VZrL2z9ysUphcOnpgUkwFTBHS0frAeYZaWfYlzn+nnWCQGnN69PLanciTWt
Eqh7cTKrAeRha3rS0ca1UnqIymdpZO5rwF6qUQCZzVqZBMJke3r1b6E+u6cEobTtCozGtLq4952R
lehbtVkRt+KLVWA3o9/F3Fv4bNGrFgMZu0voWcAd0e79EtxwuSurR/u9y082k0QqPnF3pbZ+UKIl
TManUU+wn1PFQbSb1kRzCpDno3rM58T6BGktjsCwdOQhFlxDdujC6WRI+36aQoRaSM760aZUE1Ju
lPWElKTr8qQuhp+pGdHBtgvcsr+nI1m6R6SnblMEGuiXwnQ1mibcT/JKzpjyYE3Q9/Yb9Egb/gl8
tyrJvXoahfnyiJsddijM6THhhQP8ljl68/nlNLoktdMbKAOtzZjxRW7SKntjM+crmbvSZyeOdEeh
vanvxwXR5GKsiZu3nXv5n1Qhi8WDHbSyBjWmFNOdeCDux5WaNR9oIustG34Rd67/lnZAEgMaPUEa
GXF86aawnE4JARjPJtqjsuIArlaXoUPguP0BHzAiMW04PSunjjmewQ7cAgZP1/tLN0zpe3USTfTa
yFTsEaNvd62vblv1B90ui3M/PfvFVM9Pw+gv0lMotllGab9TkfNvq2BFhq/kz1KtN9yEW3D+oxEb
ddFSBIZMZEhhcHHjUYYQdI6E2FgLpS0yCiTY99aPLHNXBg4B2+pB4uqEad9I7cIpbMMwtZBTiFir
9MKxXMahsRzciBr5EAc7oivevtqpolyD2LHEAUYO38BlN6JuYwTFCEj7/eKZzmCJw/ZHEnYn2b7u
cRu+rZJi/x/ozDX5rKqh9TK1R6nDHQ/ykzEmHwzqPfxnqECHbeTwGBd11KG3ubIZq8Qc5aKrJLvN
iEOJajYdtGaPQG4/LgKNXzFDoWfjDeaFcxCshf9cpbaPTXKzK3TDsD9FC0TgKVnLRuSWqutmQUJr
vMYpRC4g3Ll/OIRNHjwTrpU9YZB5wwDRmwuxv1jpjcWLVO3D1YIzdN8OdPoLLHT8UbNg09vxnhwS
YNeqY0qoVCbbdQUAuRnlPQjCYxxUvydHRQ4z2eGoo1WMajtefY4MCdSQ1RH8nlcZYiuLLJ8x35R+
T6wT8MEPAmeXKxtwfOXZfOcBpidJNg9bv+mIoy5nhXNfZoX0iuFXYEoZGG8O/1Zd3RdFKKK9+PaV
ruQjq2bG50y/BKP6COyneAW5BfJSbeEcSTW+fDakXqKpbXgEqp6/jhOccTL3bXLjQs/0On1ZMlWk
i1qf5Xj5jKqNaDYFMd1mPTuEq9+QloUOIOAe1EtacrFF3g9lvpv5bWpKwyhb+vl6xyyTBSrg8GQa
/u351P0PN8XgsfdBqiZBGSqcQOfMqZjQkJD0QYUiplU/VzS05HE0fbt6QUeKe+vovHXG66AWOeG9
yH5BKhq6qLiu9WDVJpWHEUUVwm0Vrj95nnJj9QEBP5ZEPxYrZtQHKrCtOpCtMlnD/fVsCa+wT/BJ
8JS7jjh3JAUtJx5rHPfCp9OkvdWXFTsDPYTxifnZY2H6RoU+FHCPrFd5SXs7zbnj69dXnNHnM5mR
GKX1Z/yNnTFdzqPCvHUCbtHcymJyyUrPBcQd4+T9REXLhvLNjlLF94f5K4rG78NMEbCUBk6iy3mi
AOcNxNxQi9yU6hrKfpG2QkB+VTLpAXB+9R6ta7osqNBzVF5Zl6L9PshCbVP1q7r2FvAZUqN/bjI6
V96xHrZITGe+1nZbrc6MRND5KFQ5GGdDf+3HD5+rOGLWbwEinZLT7xusfd4BG/YYN2cxMa5NeQqv
8bJABD7KpPMUoaGb/9Vg1OmvJH2nT3OVj1va2ZDaStRBRuHdumOjefwT7bnHOaG4kb9xOICVg5Ae
vx0wpXJpjLjmsN9UqdgQsa9teszXAePsAQnMjHF3er7ibxJ9NKlRUUL29bwJyaTJUbXC1HSalOFf
UDnx5H3qDELEQD3n9VRx5rOdVnTaSKiHleMBf9l+j0nSiHipjcqTinzpT/b8Ee8OjbhmtrGlkYBw
u6S0wKXwLhkTbY2mB5DQaPQ4H3FFqNGt4u1rW5PyL7sgCfuaCX/JFMUKJBnDlVMGQwIlJvRpW8NL
0n+3Tw4CPT5KecZiVcClOcNJYYGrNpA8UrUJNNpWg3D+pI0P2ZivPmzGvvso8r9GoXrsASglcBCn
f0WHicqCoHar4OjdbftbB/UR+JqgBTRkGZeAgiPcT7Z6wQukujlDLvTnKyx8hRXgxJIMt+dXT5k4
YS0MF7Qp8U2EIvlmJt5EFFka+ACRGCf+f4iZ9HXLxlevBFwOcvW8J2vYAoOi2oWsOaId6EdlqeR1
Eowhy+SwJOlB4RZGnuxvXu/tFQLjN+RzsPFy3Np2WQtqm5TSLq8A4GlU7kbC+aDVE+Z3n+kOl2OU
xAX4WGz9/jWtJe+cKXaUmEtbPkOvgKMgan8XA9nwIllSKPaHOH8rUgO2Okllcx0HMXKt8BC98v6y
nSzo3GX7RQ40Fuab0kQmpK9ebmE260wO1C1D4SljYzWP+rUmFPxCv+AsuHrqgO/RZqXuN1eg7Q1k
5ZHLbfCdTUagWg6lzN4AxPcueFwZv5GTZPNE2Jc6pOLGWaK7BGmTaaU2/RM+UZPgm3Kyd+Kb4aSd
kZLsklovsW++e14q6BZOGn/3mK/jW7iEXNDSwIm8kpJJ5ld3wySLgaapWi/fMpGOZaqROsEPTnes
N8FkzdberdwdW+sO/MW79vBGkCGLRM9yYBZ44H8WgqvAjBON0tpSO6jMR/GyMT74B3XBL8jcBlkt
qa7SaQnzUfoUukPb5HlhPeBG8xLNP50j7na1+5hHh+bLZ7ZsgBcrNcwHb9YKQYmq7rae2oAphzjD
qDdbsmf4lDJ45vDxELW7gE6O4LkpdduH1aTRQX1eWkBOKxkcjEx50zMBVI7TpRXBqJpzlssT5gI6
nTUUGvKJLtU06ApyAf+jIExW24I/jtEtdzt+h0F+U4yPNLANUwkH/chUJ8qFLR7k/cTjaJvjEWiN
PlT2VUF/FQJtc+cybArGYur+bLp8TP+vSu0jnW1TChzptfI6rCyJYOyoqUYtPUgewWBoVM9TRXC6
A1AoYmjSyn9V0Jx7OBRHXDEGbrKwEbY8C+szVCAI3lVcd4WtiTnoThx9PoBv1nAX1uQN7rogLQwS
rhTqv8UOZKO6IZWfwcCcreuJzuUDxZPWe6ODGPWTh+N7urnDchV8mXYJkLYH4jhdCtoC7HT4FPtZ
JlWz/v2eB0MyXz7j1LG5AYP6+4QA4wDg4iciXZ0zAioq/UD5WHHELj9PHC65CV7pq4d8vLDd20xJ
ma1y2obXf04vaa3MniiynnZ19Qv9UcTRgDMe1oeNCuwLs1ELHl4cX0cDoGCrwiRD2sTbFs6sL2E5
R57j/ZB3pvnS3HLaP6SyExbYKpJv1eSrCfjvCZ1vSQfxcL7qIi8J8XWkyX8oCkwT0lkx9JM3B3n7
2pXR94mOWVW6DDlzX1kwDx3FzhvvFLe6hWZ05xA0xcOnpcE0ZguTI7hqUjDPOxrpGx63nmgt+5pe
sa00d2bdbHu8x14GNA0k4wjOPCsibwScS7supFyPjTh+6T3eaQMok+bnL5v7cGQC2T86S287cSC8
AWvpui+m+xQhYibzb6xJGivY9IihoKaiX1q76n2++O6nqxg2NfGv0EhUsxlODNiuIpwyAF4cQvPQ
czPD8Mb3HYwk8kMDVYpQRmhcZ8TRmfFaY05FpYicvskyEDqc4acCu+TDB85ec801wUOm/I9DFoey
NN6c8VEnkgInLgsMs5+YOTpHLbZq12G45ADKerDhTv95P7FPyzUYLjuWN9HExxpWlurHZW6xLa8W
UXLk2bLBSMUnijraDJVVA54hDEs8k1AM8kGTl8CEi6b4pDZakMfdCLyM4COSsjhTLBVKN7JhZA4D
NPEt7JbW5HDb0ExegBHYLqHTX0oRwSXami9eiX1vbMMoJGNc6Y6+pHUq2DyvW9cVRBel3Cy8KB4O
vqhbG8LbrHi2HoTJ/kNijAlx575s1mGqMvGfed2/gIt2NP8z/3jAL3J2gnhqQgzSGDMQ1yIuDI59
ZQlEF8lK2Bf1yAi0SlhQ/SmftJKwl6Kg63sNkeHXdqm+RGMgnaKlOv8VLFIyBh7DO3VZXBhd2kfX
Gj/LlHY+KjSSQJArXa/iJ5/KdlyZWWYvg/ctY5I1JqlTF/yBA4p1AnYxQfZQRz+v+z7Lz2b+pUCb
dY6HCprH30JPi/MSFhJIKIlWDuU4dE+C4dV5CwuO+jHDipYPcHECBCk6SO/fGrFLiQy1ZB5l7R4R
f9Go+3jb5/WqiwCqYv8oAI7eh0P0cgj41JKaOCvolCrbKZmt6ybNHyT8dCzIk4FaLPFqN0g6vNut
b18Wdw00EXsm0kD81Y5YZDpuSBOhZJ/3KWg4DejcPq/fJBfOLyTLKHd01vEIxhWTHcVivvwRJN0d
vTvZsefiPuMLvYSAZ/qMV5yAUOoqaL/TIvXswru3KSji/8/pgrI2bwdeTMTE5Ffk0BDFEEaNb7gi
HuxscFajS2Es0BhEll9RP2XZW1XKTHBgIUxnBOFxc+EoArA/w3nQ0c539z0yDlg2DWAMQQ9314Pk
IbyX72Etr10m6Ai3suMZG0qsX11n7YZhUtdaZaTO/Po0LSEF6y162mCITicyoXEpqr3aq0HYGSWm
GX/j3qOHGHc1misM/zpD7WfJzHlY98IpLC1QnlaaTkCpwzF3WPSFA/n7n7QefCjFxRfNWG/ejwvp
UGwsiuRqoFTaeyKcjzQPLEqHUyNoWw7+T4ZBhp7dSLTgG3py+IlAjmIQadublS5O4rFfomdk8g2Y
KPpPeDxU0rVIcL1gcT0EFtju5OuiR/hfkPjOgNZyVZWfis4//jfQCsGgOsBuOfNLbuFhdBpGSfnP
sImAUhWyTVgKpCTWxUx9AcEJqFZCmS1B/fHyw9ngvJPhV8vcNRqqBOih82REuODg64nayV+hVw6u
p6NvgtcCOQpPpF9rdwth/nu+rJ1mlaAlYvJZLcgcOSwqrZjRFE2ePzwLnxDK8f+EhVBDk6dSJlVK
RdIq4XuGiGk0/j74sd1b1q4HR4U3UEXTVLQeR3wPG7DwS05wWCVlOYQI5YUSRRsIfW9Jc05rFPBm
vqemWvwKLltAZM+8Amwl6tg0RZ+WuHIlrQqaMunswsFPDu7R0NjsORCiEQ1vU3iSLqH1Yi0moDUa
LxyfRyotohLFkBA9iV4tJYg/KYfAHsH68t3WE1CFDqBbT+i29z4zINcPsiBXfLvs2byyrPfT70AO
+rcD5BVoQmhx/BAPFTTM8Vcf/5/3lST0rmD632Jq51da8gxU65B4a2zTvBAoTH/dCFW4f1kEjSMH
Mgft5aD+7KahOmz725VXfMxOfshaDd4QxTUsfSK0QtpH4S0hpOjqDkoiufXFnk2nGoN/Bh90ne/t
gRopjHEpnmtjEi14EFuE7aZ+7R2I0lfc2anq7e4UVbFBxx4Ssz+KdtWyL4iZSITJN92eRVZm+Kss
zT43R5+7VJt3WlbIaWJs3m/JYfciqB/BY3YPorkPtQc6ZbvI31ZUYa1xRnmp0QHzLx/uljslt1KH
ab4+U9xajXOEiqJd8LdFoD4BAtVipjmDgeKQsvDvUh+1h6zmXLhfoNXnuK7Kuv4D/kdf8fZ9+t1Z
65P0sMEiV6SF+cisB3TdBwCow+HH7I2OiMg7pM2iQysm2Vf1IOXKVf2i60mVUeuP37lb7QkZMiq8
H8Bv+gRtCmvGRDxEiM1vALBjtBFwH+0G3Flh9B6TkIdB1+z2eGBq/92SstfEKqJz4WutiEsae79d
I9ao9xuV/Wy5lvwp2vr1La90Jh7CMwOq5+N38gCUeCgx3uxHfYia1yNSX6xlqG9qiIt1hL7M+AEq
k4CTPvE2lFW6P+ZBmZkJPV3CxUzjdx95N27AgPqt8srEkDjmu7BORfFS4LJGYqpAOkrvWiXKjvOg
ca43NXzuZLONIsBLG2DHC4jr81rr1PnHZmRd4AefDC7WFXIInWB+H0iri1OuK2UzkbKMxcPUKcYi
YL9oarJRxHFe1t3lgJSD5Qpib7YokK5RyHYtIVcq8+b2JtmSn2olrZht6npyXHGbY0oDcpNr69kb
y6MAK90IpeP79hVtnSJHwUPd8hamhNHImDVSIMzn2J2k7WtCnUFf/WJJOHDzOWJJRLh1HL643qEC
05JfDm8WxKN8kD+xZpofSx+dpBJRH2iCNZ1PslLahjvEe33EsaXm16MGmIR3N6p5x+SxVECjZ2jE
4quaYPtI05T+NHaMOxxwkvjoQaHr5L1kf47M6p/3YRCv+FDOHoUxOCbqJwMVlw0ETUuwprFTZEr1
nqPUJV6Js+361ZUXdlOJndtaelS987bKKa0y3UVL2jQUrpnSjBi/I3MjW4ERiqe3+MqyUGQDKTrI
UjR2oQRJuaEsbnaSJYDIMMitzAXYR8s81QH8qYpFGoPGG9nAJrEuB27tcUxVNCKLNpVC1OpIwXZp
hze8pWc4b9kbN3KWtN6cqoIKxFhtpCAhjwWO5l1nN7YPwL69cW04YuHKSGyjPrzoyuk7iWRlCsyl
0ZDL00IZT3hnZXY0CnDBIZuQ93I4iiFCCEGDIxLD1T+iBfhC2MaBSlZ9PE3TPE98L6qs3xWbcv56
BeNmQMlwhAePVV1J6ZMTUMH/dZwX4BER7MxunwtIlEiZrm513ZMjnZnJcf0fmFtxAxN5sLdNt/X0
3OPxFzk+lv6R4ikSgP8Lrze9trqzRE7SPjqzsW/VONpQBdnHItNys8Ut7p4DjBSm2DDLefX7xUr2
YMsvmrJfQX6r+p4AIkc5Ch7NpgCBD8CftE0t37SIWRuKccL9SW5JmAiKJmL9mqRIb5gc5KKVWKTg
2rmWvNPHsoK4wyU9xAZNUf1o5ePT6Yc1kXCV/HMiapm1MM+eAnCDsI+cwdDFG4S/5goTuIiEfqvM
8LXYU71N6HpDfk86OvnwmwqR6zVRvTqslIwHDRLLJsVWKk06BeMhXStFtsedToewOcjU7Wacn+zG
j7d/+LAgahr+1Duw62077WNkyeb4jsea3B+JxF4vz4XCJNX0NHiHN3MwziLHYAPaRTn0jBnLaM3E
r3cFt90ddwGZHzb4aNyBln/3r+gpJqR6rzldOjnTUGP52fbvxrCimi4A6gq4drgqCHQE5sDivlUp
NO7q6TKmRwTotpsUsJl6peMtlrAnOS0UsuOlxttJY+XnVEDWcg8aaBajStKyNFuUSoMfkIteWe4t
AqKTT8ia9if3faRBGSuuoqHPCqSWTQQZ2vxqWKNUipnWV0leBdFRPa1YciMdvbyfSlxCLCyO6aK8
/JbULe5KXQhR7StgIDnK0Vs8BPfiTD+hOWTnVNNQDPbD2ApjB2lXiKKqXQFWGLPxsHoHShgqH8CE
IhympysV/D84uubn636UsDN6OWeFDNigOIVZMybpUfC7a8TcBgnzo9Qtgp6SuQxtoQqeLZQ3+jB6
pgXGh+wn1g+K1exyjYr3EWbKq9Ablzj/gvd19PwBf06o9O1NtL0OGBB7X4gOJdFawOGMf7IVbe5d
iSpFiPCSFuXmc0zHfnH69C1P1tM1nY5zk6G9prhYE+0CK30MUvv4X4B/YH0g7esmYlIWl+tFuVAv
7c597dgRFum21gOlKipPhSS2HJI5EV4gNYXo3CFuJ5igzem1p9P+wMd+lWxmxPcP4dwLsKQXog46
Xcpey6oHwep0cDqODPljAWMzClk5OcFuzyJx8rkc729T8VV2t+7RytXIYON6VWmR+JntL1eyWqun
xg1eQRjb/Sp7nyQjnJRNyweMtjR5CRPU+r8IQ2FJNsuxIXg/huAosdqJB6L49P/5pqMU7rV1245P
ugDvkQV7VfdmprblIj/mEiIyaoWChI/lCzdrQ7unpxAgw33kTtSoHyXYxGK35lfdNPJtf+tW92w+
JS7Q33/oikSsHkpXhFnc2laoYN1Boh5fr1IkKgzeCdW7JFcZZTthG/f4MIGZRpcqofOlupNIg4kN
GtED9d/sgU6kuSc86gnsJyBJ6AAWYjpaoTp43IZpClDFSoXT8IoDzpWGGXxtPJaYys1+K4U11oO8
W+gLWC3fzNyc8jxAe4ZlRRoBjcoApoPh66HIWy3Zm0cSaKepTFwNJqEyEkuCXKLXraS6KFn2kDL+
00jzhMAJrFHE7np/aoZFPi6TXdZVVKlJFI/p7g3ny1lnuBCIEMdiAMdSuh22/+NUDytxjQRraCRq
5l0jRvqzd+//Po7Ydcrd10vRlE1UUNrgTWGzBoIU9y+3ATFYho7rhLJGdY5VB/gtL1BzqZLF1VjM
fSoXDLmpLkEGMmgqpe3DsdV1xsnX7637den94pcuYDgUJU/Vd11hy3hoUiFnIvh5FK5hmAyufUMw
Xmyn6NsbCfzVzHCDy57hqUektFyL6hxSB/npZoe0Cf+L1wXi2as/+0vl+RiQDKZTnv429siQuDxQ
2ahyxY8zkS4Zzhsawkc/C3+DfmNCj2/CZwqsuNBMQc5sWPbWcQiBq9sce2s8fVhfIKj/xzGENzpO
+JLpbtxiQm9+O0mxgD6CQuwgCd7lFjQ6lwO/T5l7w3xQvfa2mRVU08CDYcvG7Y4696oOkgQuEZmG
ah2uWsYp7qg4W0vmGtRNpqDpCMlGjW+mzCnypkr0NEvJhN4hKb3NGyL/zU+maLf8dk+3jLLIQBY9
5si0Zy802utF1td/yTVO4bVKoQFgONkeVsFL7woAOg5XzpQPBK4plxBF1aK+uW/CZsXsPbgIVoIi
DjdXhvcl7Vu0rEX+abq6rqfuJnHqNMewQR6MuPJxcVuuT7Ym5IZpOmBKUkP2ORPVPcizNvdBxM2W
iUflxMApAkNguXElTK+i1f2V+vz9xg2/erKC1P7GAvPFDBF+TDQ9ueEinsqObI8G3Cq4APwr5aZF
/iCL24cwxSZebO2s2qWOPQV/Xn0bmPzTsQ5/P9Ms6kQbRINyLpEK0k0BW6yuDbCdejxLhCXrrlAJ
raqj78HeWynDU0v1lzu/PMMMh7Mj9syLnx2oT/Cggr72ralQ4odKpEWIuVMPjHbWaHaNsYDWO9si
jcsydjvvHqkZt6pfjASX2JNupnSp95NYqATokuxcTgPx7XH41f8wJPLc6O9wdhgyunVEC3rEZ4AY
j8fwa5wywg+dUAHqLu1n+zuz8FqulrTrVd7cKAjjhkeJeKolX6XT5R/+pFssRobXpEC/YZEH8Ac3
QKZEqgR+wknM5SPaVJ+ImYWIAl3P9OwwuFPPEwBSNqv+H7LYEjZJZlqBkZ4CWJvAedTLo6Owcg6D
EgPadXIrmE0RXtRrbzXiJKFYa+GohlrSWoN2dsvzgn233NF91xI2osULB4Ei/eALTg7+9K+gHURp
tXnb1zAj7NwaHwhuWT4RYmAHvwY43UJjw5MIAbeYjZf8Tqyd59FHnZZqvNrYtmfQO/Tfw4qeS+NU
Fg70WVVLwYKZPy6YU75+yjAA2gGNHBiWw9ZH6X5mSnrPamsidjyHYaPz/Yd0ZDUC5HPM+gfi75dv
KJ+tnPpZRtPm1m9nUtLstElE7KPinlVosygeIfFDB5eGNiPxDJ13xHQXMXhexWpYVIj10RSCE5EU
Temv6khyjZnRR2XMqoI7TedfaTXWIO2g65tbRzlaCz4z1pP5cYKxTx52mvDSPo8G+akcblx/xLqu
zt8Ft3wzWmOFMGdQdXAKQT9rcyb2v6JA1roETihDWTdHAMNkYPdkZGKHzs52wqK+1bzpUtddwLyM
opjApcQpmPVgVAmU8pC9yHsSbQ6b5YWIDC/2g9TU+hbU8vuYsrnedzdqCXc+3ZsN/Hp1AwjlKPpt
k0V/5uU4D3KRT3z9hersFOF6Zqo54CBm7obzobz3NzgjB8d0HAGiCpPe5/PRpDGuy9u2h58APydg
wWwJEzTsPE51MNZJKzn29hUAYOErmATYGf828dNppQcyjvg4k0Afx8PSW9YmrKjdcKd+KAw6JQTb
uiHzjpSgd0kZZVueS4xSOWcBLM3wjj/GtRtc2UcGV3R2x78X+oW7XuOtmdrn1Z2+xNjKiX1vbWg+
khaW5GTfduHm4/dBjqoyWfflOpn4iPeL/j0PA8d531tUHeUgG+Iuykc5Loxm6xa1yzSNl/ckODfG
aOovQjcNEU6xFyOtsWS9f4Xab+nR8e39JWCzO172eAd4h9433yI2/8hO5w0Fzy9jWtGdDFZPoxNx
EQndvNIGnDQkGebAsPt9nAB+EUb4a/ZzfHxRCLUf3U1YG3wwDCaU1C9yKSCOqZDieIJXDMeWfgQL
fn9JzmLd62hUdXdnFsb4TsRfx7JVJtrYSZTV1FZUydf16BLPRvdQ6b36QE2CIRMI3lQeEQE7VqLC
AgV6480E1s53aGxLuz9QXpO7VbjzUu14E+ZBDIUoBl6HilEoMyol046dwwLEQfamhxLd6KeSihSq
TQlDlVcIAWYI4r1CnrH44JDsI7c0CysqIF7ANS5yCxESSS3hzmPVFTIjTHQa1v8gsK2Jv5h9Iukg
jNJiVL4aIzQENgQ4quDNtcUaaXaKp3uVDxNRNeEOeoI4W2w/AsaDuLSSDfP/smJ1ZN/f0lVAlHFP
UKVy0Ul2BKxrAc7bEoB0hmxFms/MX9YyJdSx9XP+rSI17dL+0gMZWZIhauyg4v9f/L9sMOVI6RqH
VTojFY8OdLIb2Xg3YSVcTPL+ZjCkC2uoZEjw3Iuk/meq3aSK2lLdsbDk61C4ECs08VYWsT/j39Mo
ysGdWzdnNpXjyP/7G0FXhHt/ZLoP02pxaZmngLUdMuvUBvL5JZGxme8lTjgXZ3FmvE5g8lHC9gMt
Lqa66mIFLypE44fizJl+qX8o77AkWN/GMgW/INsc5uk+gikoIvuGoBw4wOmj6+OVtohOup4qJOP0
nsOO7ByHYDcwYDm4gfikiMSrB6lgsFLXjNn+oFpyNPlE7zjusgQdMcsk8uuIQhxWMstm703ROkoP
SsFFIxMxPDkUztMMf2FuNuBFL0C7zCNEHJ2qL50KJVsDKHfwT1Pt5wyiWMcMD3RMkLXHvFL4Jiwu
xFcBJEhqPOkqDkZ5k+7FjjGpPmFlV5L+ur/G/lecUlejw1tTUX5AdslMct9Iax7tDk+zthnsH0SD
KOUWsvJ+lvj+lLJuS3sVZ5jejQQMOqbCWlEiVPfS1QxPsnbR8ljKT5qnLj89vh0tTQK3CpQjK9NS
T/4XGnbXfpNZIfc3KIjzXZy25+o7K1pKXEcLs2XFeFWyIo/0bI6nR3BDkpc0hk9NkKr8n9rUUR7s
0ILmreGZnbl50QpNP547MiGk26EFsmAnpB3IjSibk3Nm5Ze21HyKfErT101inz4MjY+vuM2CAa30
e8F0hBtwf+34vUrWwI849kVTnAcR3sqtyBI53xnXmmt+hNA6YHk8NyY6ai+FOhCAxgAecNH7xDgS
FNDOJM5OYX4xmktvQaYaznDDKOC1C8ZVEJSdkj/o57ZloEP9HDhu9yUKKt/7G0srpKPtDgydIh4C
fNNYWuR+tAm30HPKTvOC9WfumwrxI2+Ucf0Z7wDf/zaZZcDXicFUmyrxcNpchcI4s3oYGpOL/iGl
FuesPSC1q9lxdlT8CQwYlu/RF6oCKcj5fHvMl3eqBOh28HR8TU3taKBf0d8noIZXOGiQ563Nrwib
hxlzeG3bF+UYFofIuNo1/kPt4rNQlq7OJkjv3TOVkxSKtC1or/7qGHMS/rg5V+RySCmISfxhPOfb
R+jA0wptU0fBlGqv/c+cNYgTNArHJ2QvZoqnvsUaztQumldXyPAOPTb+YIKjjaucID3x6FEa94Ym
x2KXC+4AmqadB/XDFJSwUzz+FhTAKHgZD4YrMXD7DtbKfxs2gaKt6l/t63WI0ExnwzdOwE7hqjCm
+17FyLesQyk6PGEPxIHl1GVL0WYf4AXrqbasd4ATHcC9SqFeunLohxzGIXV7GcB4MNplzfRT1lQt
1zcv/LqoGzb3F04ea4ljYllRrkL7YlDDBWuTuu+hdJhnW/JaUvVU3hqL9LQ9qTG4vs2ThlIabPoP
SJHjYk07/MRCRtzqQ+448hav6xkkuTHbYYJS+wudxkKHW9canhZcSztG1Ftf8xoJOJ0Msc3CQVQT
VDCGAltnkEssMYkXrcMdqOn+Gu2xpsNNhuyCIeg8rpTznjcfSzRaH7fibVPkp2EXipraAgafTS5c
8a2w/wRds3PAqEtCMlTDIxNQfnIm4FVblmUSHP/HXCds/BiUCSNQL0kuo786z1ROB39D0q4T3M73
h1TJGhkvFgzhwRuruGB9REm/oU26ShpWwQAH2eSzdInCqj40BDn5lM2doJi623slQ2OF3JlhMEoR
6xVrn+g7x7oy22XO35i7dBfdzFO3WgYnONhK3AM7oVLzTAJ7N7D7oKlYExrD8X+uPHGYwAkf+jtF
qI+SV8shYDwIc0FDN4WELVLAk5kOwfoMPJWaYE5FfRZWrXEbSuBN6w/mVeKQEaWkR4hYKaW15nZ6
1RBR8VO+EoAaO3yA+UGN+OTdnIpO8lIl2PYr2qAz469wDlvSguaZmASu0feNKnQdjRmE1Y2gXEvC
ZkEHQk+jp5PGmRjjc23J7w/OixcG+pE7xjFqdz6a/xxByMp+85Hm1ErGFUo4U66TkvDoO2c/bb7G
j2ChhI4YDbFrxElUJOa55TV5SbI6RgGQsQ+Pw5E+MPs42/4Eqzbg3i/lDjUsn7a4lBqie0TfhjIZ
VgL9gCnMAfVztTKrLXEEXnLW2vGg3LlHfvZn2FUAH2BoK8n9W9htp914fAoBzawv8bhcUEURASC3
AwEQ1kXcTCgMcYIrJN7KRvhS6rT0TMC0V/dA85FYz9UMdaSMV9g+a6NnhgbHVtkCYbc4Hg0IQezd
ajc33mIUBme6VrCUZ79WtCT8D9HSUjZ81okPko7D0Z9VzfVvEkLLnNE1vRwtrH1oCXhndTlvsTv8
BpesxTO5s7qcPxOlvrf0ss0s004alcCwL/dpN86w+JEugkNMjyvg1b9aT44C9FBM6U/U8S5MkYIt
mXarVPK5cgM4ukZLy+NWQFMxzNjSv1NUDn4AcaZSJp3UzZAmoR34l0RCy04xhjANuxtgfqNkbaZC
RkUPDi7t/wYR/cLIU5YvGMy21dUxyCFFifNArha8p6r5XtZbzkCI25vBnhUndREE1mDoXLL8g2Bs
xtaDqJdOROWx5E6ke6Gcq+Av4WJUQ27/2g6EDv/l8v0FQ45doHnqoFVk+oKgQ/WaqyvY8TuWZMfy
qd+9nsiTljzGdDdOt8HpWlVF8hztgkiKuocUjyOXW3pZRW76MuK/FaaZZYtkT19HQYrSxnSof2mJ
TTjUDVxxJQryawfO7PIW7dL+12GlBB9xIHGUEIuBnDWOaTy+rU1y68RSQxOG+ah/X3S+YCMZLIoc
53htrxKCJn5sxY25V4RoXIjdE8CeuqeXvNBll5OnE/302Xttz94h6Zsa41kq5T5Aif2voty/8Kj8
zdv5Cajr85Nd4mZGH+3piW/uwI7c8/8+uMrx0uGphdnKyasHBUaKIJgY1sANy29v7oH3Ao1IjmLd
ce50cZFJspSS9rI99wtsEC7lIDZvF2sOVRs8ywzt63x17P+66iWPBoEHAViqaLYF7mOdn9Qb6lR4
mWn497CIrj0P4/U3jn3nOT9eK/VwbGy2oulmJ6cBnSdK1KQcaqHW8ikpZw/f9hGuVUyrXRoSRV2x
aGmpObqJTsTLQ3SLzJbMp2fbaBKlFWU7YvnHZ2YqWwBtQJf7kQFRESCmi4Fr4q5z+k4U2YKPlFsW
XgfnyqoLnCNMWj59kvau15rqdGxisiJUWJxnfht8sVGgGYxyFz1pagsmzeZ8AcLf7usG4Y3kLfYy
ta2H3hX9HwRCSNyqgbXIQaZ4PQdoQ/gRW3YEgLkSsJQxe/rSsFIVFtrLmDn7/Dop+NB916/tHFGq
R10bjKnG32FEg+/mhY9i/mfJknnDRE4Vak5OwZplxGjG2FIDPY1jNUzwy8H8vgbYofjAMjsEUZF/
uFB4irxAmbuhEBFNKE13RaXe5xLPdRwcfqMnvSvgr9NWZxnAOEZNxPXX5Zpjsc4eOSNYDd+gZAwm
Bor0E4wDj4DC5DiOMlWhQh1nzmGdHNRgr8WYuhpJVNWDxMoZA6YL5rKNk9I8zmTQ3HM6+cjV7+bQ
i3AR6CmIXWRvp52IBoOduHfPltIeJvd+5fCaOEMqmCcBMVUFSgWopFLNrYTu11f+7XwTFOeulpp/
0aklY0LpXYuEHa1fqElYIHMAWSvYkUiIxVm01b9HmIu6x8NT9o+yCFMOg/QhrRyhdOevl283eFOG
tmVcYLEq4m61DwZAiTYTFItGUP85htm/26znNolV1VwEqoJvQxRY5kqkTBcKHzWzDveASPMzf5tP
OlIgTs/fDoCczU9GT503ydND/HbRlW4lsgyOgVPHgooTD8wp3xJ82f77bjfmvMTjYWZdFLE+rhPG
tn2+g+eer4UZZPUSvHhdzSejQHlfJvaRil5gJzNSWlkmFe636HCyKgusHj00EmeaPgZFik+DFe7x
0wydV/631xWTqZdhzpU0Lxr5x99KvVD4P7pttUIfws99z/Q3f2C6kAjhONaPDEMh9P1dj601FME3
dq5bzqUhj3I9sAoSnyiRtCYq92lLf2hBUFIiIy2045oGbXJ7QPiLDeuUoMUyIjIVZzsbtq8TjTnL
IYXZkZFLxKPeosQuRbRnrZdq1+6eCc8nkpzDhk5lqtCSZmBnxl9uMrfs0Ki9HbqRSRP/gnTITSNk
FmDcC+ddSrYrjLM3XGMdv4guJ/I5kApWTol+Lczts7WK+Wlie1qTi5rMmCaUD0035LxGIteEytki
M49oSlIWF8JUi6MAw84gh6EZyVk6Q+pCojf2JsczJs2z04aSVNjhNyoggl16xPbCYm7/pmLY5PrN
CSUkrOvCNVlj9IJBudehh7/K0JBZ/xdVDYjpSM5ccmEArTsagSxD+d1hPqGkuvkLU55HmjbTdDlx
Ne42N0meZEvbfB11o9Su/IJOAF2Q5wAtYaOZzRGJRkhKs4QaSivKp808qAlyASkJRyTYLKsZVRl+
MThswZBGSyPGF1wdByfnino7kwvZNpXP7mb6NPdCn+IFtZebm/GLiDE1UY6Af47OPxSf7gUN/CAM
5Xld2tQs8y2Ccip2sPPSo68xfaZ1PDb9U/P4fJEXsdm9IbvFEQG2++FL6MvRDlZHIYCbf8c4dECb
ATVu1D+7y1D+I+KPOPrFvzEislczNRfahAvIioq96wtr/tKwlCc8mLSA63t50ReoBmrWiZgvJOgV
C5SOXv9165dmiARIdh+HuRvNYNNVL1NnkU21n022z4ncUWpoIDZlNCetSrdhzCHp320Stp3m1/+3
pwx4Fnq3U1+4RGEfyJuIKOoQZtE0W9SufP/inFmfVXniPfznOjqkpiglEF6CJzcJdRkEk25ADSMt
O/SWT0CxKgy5yPyCC76UW7qgaGEPa8C3hHeQRpSsDiX49bs/OjEeY6WEGavZ3+7w4Tq2rrSdvm7C
MkHBdIMWrzUomZgvZjY1GFGfkSXyJlIs3Pu1QlGDYIaSUcVqpWBdbiB11wJHExROoYVdwHgmv4rY
TPgCNhojBIvYF8Y45rpc0qm1qIpTPuSdJ9D7/i0yRCrwO2roishFmeoEzcdHOQYHRKhrII8PLRtb
6m10MkTeeY+pacJfWliErqcIAzY5KACeyzyLcbMbBLcBjyuZPm4Zb4eXNzXSBR/Bs1Q1gPCXVKkI
2I3UeTTbQSpOFT/KgfSOHukpHg+CobKlD0DxVjuMkWajIE+e8pIwTQsgZJq6pMnktFQLx2es6MAS
anQIGc78kd9sw5vfxudkYMFPOYhAqaBS66CFjaslPtzz7j8ky3T02FtEpBKBsHcYeT7FxqNyidxj
mcEjGEgkTTrwD/kQOAvd8h8Igs7c8gxKEcwPoZ21YMrjzzlo9bmdE4x2eU98+QDwP8CWH/zuxHpL
8tn7DYY0YIJp0cbmuAuIQiJBJXSdnIBeJCx/Tg8A5pGU/Os688BDDOFGn6y1C+5wYEdHm18Z+vBL
oV1enUw1rem5gHRaEjExZ+xpgYlZV+K1Y9esv+44LScb1QhDGfpp6i0ivTcg99usA1VKdxLQr6tE
fvcKKM5z+Tz5HaMxwUlbNhVKPUhCg29v0m6bMRL0h0Vfzje4eWRfSVcYg0bndDpOe2hrIhyQA6P7
IVWhP4L0T86hvpb8PyxD00RUzmA8RDkmZlucz4Hb6THY5c53I/cv/lXW6cXWnb80nXlDIKAtHBwM
UBZbIC/OpAD28BZqz78uhf94WbdgO+B0qC4olDrwHBmxrzoClu988aAsIZ9Jjnl9S6RFuTMn/TGu
4A7az6C8T2BVUw6Cz7BtiEJ8LDR5N3jlEbnUpzoBtgrNW6JJKDGIOpFWmAp49Umb05GvsnjCVmIP
JmOGfYRs0ykIVQaPjRV9EwXoTeALbBpdKKZxWR6x/nTT2n6uFftv9LfH7aLkCsfNfyaWJWFbREYn
jYp/vTmkeDYo1ZD42w4p903mTouSgxpYPzuil1absWnq/iRlExDgnOQe3rbEfjwFEtdCzpudleRk
MShqb0X5UKxgpqHmYKig7Q/HjIxNHWpiXkiCQXGsWKvThuLIJqaTC7J9nnyneIbJeVQwe9/At7oJ
/iUnJ0U+AlNa6NNBygaVc0b07mjLvM+JzNKYh/kVZd5/nOXiJgt0DpLLWWdIcG6DNmGWkBg+t8UP
2aqEg16kFhYw6h2tDf+Mtw9V1ltqzTcozcLG6noxHyqLIiXBUfx56yhZlrqAxkf27PWeLsfN2Fdo
YoTa1NNdOtiUc3ThVDfUojJ1cGJpzstXvLte80akaBSM/kTvA70njdnKvirrDgbhYRSeOiaGbo8J
ci8E3y21vnp1EcVya0AqjwKBK1+yzMb3qXg3GOCJSLz5IlKijqDQB/H/k3KjhyjCW2NOKeBWkN1C
egVk7eKlj+VqOAp//ymIm7unXXmbLOIb4XUwk2Tp/34uiLiHZSl/LwsqxwX4evCC/a47Sj2VZ+8X
JWjj+pKDAEYO3IIj4VP7DwvrJrvOgi45hfoCnOJGLNdnY/NeTEU6ZwM6OyeYvmAqsRk9ZDei2bun
ZJvqd93bgmi6qJtZcJPOxDmdCI1vxZFKly6A1tpDo3Psj2AZ/XBsP5TRMO5WkpJUEqnK9MVJZZ7i
o/3zeCDSzdMR5jeDuGnuvYqcwXSHIaMLWgDRzkUpu8D0dkgA/Xa/f4NZQG6ljAl8o577LJI8ScXR
h1UhhTtCwGmqgw1YW4UOqe7NQTskr5rzXXBuo9Q/jtq5m/w1R/gKUGqk7R5o/DNCtmrVGcSPF9cj
NS8xMGFx+fvJTNEmRfxoaC5I3DIPHqodwbdE6/735oJdesBxteM6LG+PzEARuR3l6J+/qdBZQCKG
6NI65+K0LwDfx9FTMmekuiEJI1x4W8IgHOo/fHrc/5ibNsCKE4GKWSC71fQHbrjJTxC1cfyGQEFH
0JgSEWDwt9taQ3ICSZwul6OcCxDSJf4fC03ACfaRF4XwsZfznHWH02cEsuEDO8RNNHiupC0OM5Gd
BpNGgZp1rAe3wUFR98ojshREZtak7mBTj8ph3myESmH8eVmRv0Mdefb76B2gKh2Pfl0wDOnq8RdN
wTPecmO7Xt73rlKI6MDOjqnobfYSDPPqrP9zLBrSgtiVncbjkmVrd0ZtcoIWoYOYoXd1NvxCXZeN
eV9ZcBMpJs960kXtbVXJ/NtJ7aklOEAlb0HNEy1+qKFzAo6pl48A1e87CHAarw+Ee7W0e2ZMw9SL
I4FSbsh/kajaDXr2SgnOmiAny9tbkcFhmHYKdo74fCGNEMCbXr6cIPNk5NMGg75bdwhw8vd9PTCK
Rc4HTdr1LGiyjJ44CPM3RV2NnSj0yUdLG84afpetKYlU9NEcO9K7sbBApgcbELQuxYeeb2JsDJty
fUJhgP4RUTcjqi+L6itlKM6eZGOeqzGLY8bfrP+wTPWhUEO27eOFpqWc4ParIzgpIcXfz3mky0ju
fBSNXhxDmY0l/WIubfuVwdFIBcreIUIZeaIQFdB3HcJvheNfqj0TQHuFHF6IrqngAYHzDbRPLyyl
KRQITpr9DswZzUzkpTqih+TbDsEcMvXfQ/NtT+k9TJNIcWMb5Oz5Er1FR8rTmkwV1OF5tFca250W
OgEjIaLPFZuJa2CUHD57nKkiTGb3E0zEpwZzTS9O9mIErvsWJmO8DAzPW18roVP2f50ySrUC+TXw
c6WLz0bXGwKf3buQZKH5UXrUJzjXznxWZBpjJEI8/2nd8n1FfhxccsPDkNu/5M9fjtYU8EBLQqZL
dkRhwSVi9ZsLNVWWho6aMYIC8wNzcLALXKy960dxLNC9HDsfdG/NN9MEpapRI90Uki+2fKTHifU0
ikax+TBvDwIYoNb/Di0mt4Zk09ytqruVYlmFljJNhustfNxULjERWb/gUVM4gzXWdtn1M7aLlU4R
c5/Mk//0jCIiZ03pAIcD9lieyvpdIyAXvfk8Typ3kv5fJhCHutRSFehxLb1LW50KDF7iEAxiY8WC
z3awEImSiIe0Hc81GS2iWfGN3WlNz8CplyjrtLQxw+dQ+PKpw+4xgWBOhYKRJIj1LShS7QS6KC0b
ess9JagRA2et2++qQi+cEnDs7xRY0EZ9G30xF0Gyx0pNSesVNv3yrvQYEwzyJJxeKTZ8y61aosy3
mTB99yYL0ntfjQ0WiOMlFbeNxU8CHKII8iRIXCz6n5ntk7zJ3BpgKP2xdQkwAKE0a07LXYgYUU+8
uZSs5nUJ8voBnaDaFSGc0zBYVZMtXRJHGkSi+UhrmZ7Y2SQNBqTV+6lCGHbMmwnRFpPES7Hslzc6
jm2O19xEZJuOHoBvYv/hxH+JOoAFJ/PrVXQ3lA3T7MB5vwlPzk8DZii2OE1E1UKwfvyZL8XtOzsi
wU2ZclQsdy7YjGT7KvlWODG+yLCkjzzywKVwgjcrj3Ag7DtYmFOQF4pjamDaHFwt7PD70wU4UMTX
2CF/FVF7T3Qid+hT3lgX19GHgEMZPYfjWDQ2stsxIFfql61xl2tCsuOBuqBaTkw0u20sq5fHWeai
E+BfhvOZFVI4AzPRyY09NUQlauo0Frz1Xv7gKasXtugt21lhMQI0xzIUrujdxpU9VnkhnpF6Szej
6zxColbhvzQZNcch2zCphlARtBrVKpvLcU3N215nKIufNolSQ3lu45rGhcFw7QFrRMRF7gILDSir
n/fkwmjFbNFMTsMxCwlcgUqinW1xRbQtesCtCmvW7CEyXPqtNm6r1kLSet5vXR+sBrMw94oi3d6n
FNFXdY/lsk0v86Zyta8e0I94lnAMwB9qtVtPIs7D5u1toPMV+9UCPgyskLvhBSmjcpOdXl4536OJ
Pkpr4FlZ4hQh2rVZ/qUuBpn4/i5PIr0moqVykqMY8Dd1WJ770YieJOLFaWR3rdA/6A7RWK3zFbNa
S011K88qXgKXMEHiBal5OLurLjL81HBwjguSbr3MXVmj1I78rIFOZZTKuUw4bsKetFdq5PwXyAaj
rJo30wV8TT1SXUIMXsVWtcNd4MMSUQcOOEV35xt+FSR9k9TV1ibdQuoBKJ6kOxnYoNxYhGElj8uR
wvx51OsnInaBnaaCAxgOpK6Z06C8K4fS92Q6K+rT8caoXQCX0+7ZObzr/lyUfk4HAw3Wkvcp3Lvl
sXoPm9p6w3PTheu/MuKhkYk/Db9g/vx0OkVYwYjJsbDUyvHnTmEBKhg8zZUcEMoZAI3QovR6SGHA
Nb38R3Uqg+Jf57gHznNKVa7ldh1s7/xnh9K8aNp0ceE5sfftwDB2iZsHUnz0dFbfpHnNwAZm6ySF
1D1GzdDUUgmMwZF+/xUsYoc9p3Eoh40GHAEvi34FVJRHCA0igcWfIVVqXCFZIGeHQ+gJTi/4ZN4i
lRrIJDhG4qN5ogdBWdYlYv4XYdpSQHxWjyc8ohN8YhS+pbM/2s5pLv5MbhJ8zrj4Enxx91+3gdVz
hyVUfX5pyQKHjhCktvOSrfFkGVk38swC0YkUgeu6I+8IFr0OMzpDFXCZVVrCrzTBxE3EBuPrzs+t
x7z47re19D4vwhM0ShJvNt+A9g1E+uLoUNdRbj2YbJ3KyqYEL3TykYMcsFFkcKc2PkvIao6ALP0q
0oqh/tudIG2rdRnmtPFZ35+jtwPMEU8Vv0J/X7qH2TeTvnxwjWqF06ysqQGXNeYo4aNIZDcG3QxB
JE/H8tdFOOUsj0CGNLHoOFbp6IzQg64tB3LOM1f0VVle+QYf8wDpf4MOgUVvITmKBhQgQMP2e32X
o+X9RND6InZGPkuuWw7vlreHtgp4WOnKaGhGotcrgvx+AuFs8SxOTWfiBcr/2XwA0XJUvxkJtFyk
DpE+kPu41805ybL/T20Y38ULFvdAZ/d/560Li0zOzouOOn310jzvdGEoN1HM5BLVPlnZ2yr8yXZW
FIak3Ll3C7PZzfG3MOO2LbcBTKh7hl3+fbgaRz3s7thDW1Hedr/APSC/nUWMS3VXcPUtIgbcL8q3
oXPrPo0ec0ATt0jkwFg9WpUJ2ewDl6XFDQ5dGAwZM7XR1I7JDdptkxlj1DaGwKlRlxF2LJY9QYio
Y2y6Ey6P6TnwT9oQ6YVv8JbbsjAWwMzNVvpTE9J2Vi82fPjtlsDQSg5l31WfQq949JrpRJ8E5y3o
F033x/LUNSSfPgr4cdTOmlVPRJlNDdTmwtvGjAk1YT2lyWs1hWRJ3jUYuzPdgwDtx2qBS9n4AUA7
FONec3XVBzplKqxt2A+FyB8ai2gduzHhJcpn/TpQVzAbwe7j4ja8Ya1P0tKGfrNlnB8LvLui1d/Q
x8fofwztTD166nYvxL3y42QXGTGHp7lmLGRDcyP3bov8y04sQSolLse2otFif4W2yZnnOgzgpAh9
fovuO9hDTFB342siGYQ3c+ZicLTZ68t0YEKXC3iDcsBEYN97PpmlhIUMXRiRf2b8mTJPYQzr0JwY
LGGdK4MmjRUqYwhaXwXhdoEahn4AQ2hoIELXo7q7ZKw/lntMQvKNIVE9+F5d1oMHNSe0mdP3TolC
KpSyxhRIr5XY60LlCP+s+4bSinWqShg99WYniyH3azN4jryrZzX5jB++i/RviQM8Uck7D/qZkKxq
9fJj0L+yh1FOUxdQqEDubbSsdFaS0d7oZqL0HiXDROJnodlet8n0JbXrhK/WVfKvq+JWCEaXKU/W
+oPRn0def0Iqu0Vzj72oS0BJ2KCRjFaZR4Ue9Qh3HvM8zmQRzVaiPBXcCMw4swBIz0MoXe8jn/85
9Df5dWAFrZ/v7GjC8WHq7NYGMayuWynmTM3rKjqNof9JcogAMO/lsx5wiS/v6YLoyoIfS3R3tONd
/RMm6BWPQwH2p1Tqc6Jl5YoENUmRJqFOxTa4EEFAQgqFaRAXJY0AOA0KAp+6F83FtxiGfjyARiH3
TrME361X5X8SduuE7Pit9+FC2BZy7FGCE6ZIbSIWxfvyF2fZGrX5eM76StTKnDfsKlHxwPFGr+Id
rUcD9PtN3RT54fICpOEI4D+BSRsN5o0pRjTmvkOy0rObo5hgp/H/NQJJOmCcLgxfC4LwPhrlWo+M
aMvAxKICXtgT9tglWe5CaOaYJETtAECeMKXSpm4BCnjtWlgfMsdByx/8PMTYhcfuPv28DDkCZaEN
eX/OkgMz/tZsBFbyuzRHOI6LpSe+XIlURy4SMNveTqvjl+ZDIwp6XqTl8uXnAaN+5d4+S0pMxyAG
VdVo74ddqTtKoUAmxtor6l/2m77eoBjYB/XtfOMVYnmJmzCr/zTYt1CUNayDfsBA+MGyY872dnU2
12WhOaBZAvgyMlBWYIRD0rO/KwDnAolr4zqgRR0hJNEGtqIjHbOb8oOoxFBPnoOBn9ibuWYqO2RN
ieCWOfmnIV46CfI12KCzyRTQnzJlKSovC08UpKUyRMdETmyZYQHAkrhELORC4tYpkCGR5z/C3bim
wrvbtIvKBuBeeH9Cbpsv/3/devcFXmwekzzpsLAzPs9rUPVYXCYZzTRxipMT96PKea/SKVpwONY0
BIFOKAgK2xxfptQsNLS0x0SPQkDsxr/yc0Dw+fVFzIiXELjCMQLVZksiQt5qBvYQ2k/s5R/RImY5
cWGCPzp6kh4FElPMKUBXtglImzabuCWEiZ9SjJuU5cxT7Oqzud0pWYWnxs9aYfGlK/uHs4xE4dDa
KQMC+Ra1lF/n1WROoxXGmIO943kNNz9ZcjVObOWgs0xecxvbIGE4C0NTZmpjjL+ikxVzCDAaWu58
wtG7A05m3MPq+xza6Lc2GB8FpwUjZb2KEr1//hQCY4oVXXAtFGMZpy+xVOv7PhDIWZrAIbYGTqZL
evfeqC5QdKe9B1UNjp7JkYf6ySy+WCetA3NY93eS34+ukLmH85yMq08r22fe03p0NH1cLfSbPdSM
Ln3prn356rrS1rifVuE6xOVHbtm+xI8sqEwqdQxw3w82lzXJUNXhwUFfhfNC99q4jH/AcjZQ/xZz
3h+I6Cd6OXJRj1fB178S1IWPYFstZeMipM5IIh1bHUC0t7yV4CDaDDKuVrENgkhtcI4BzYG29Oda
/sp50YMeXP4trQjXSkKFFRq71WOOSMDODd5UH4+qj41f2QMuPvedYJ998B7RPphtq6PjkE+I+eAO
maYoIqTLVQFE2HwPdTmvZbevtkwi0CssYJNZRFt7NupnTlfKvw6x8JmTYl5mZFFzfKJJuL5MLb1i
RUplmmp6E94KH/Uto5NpXUnt7R3+cOj1iosKUB1ZmaBM5woUkkYD9dSQC9HRV0ya667KYNKxOyUP
PmP6fuvEE+jSTdXKNRGiWi4Kd7mlnr01P4ZiLbbVFGE07gN72A3kWdVxPZjCW6adDM9WYmDdTE68
p9rIlp5w5JpZoXaK4mGk/IQAMJRfSlkMIz4FhLJEQtCorAS6uYkNKj3sErjN46IXy+CzlT1HWm1q
oY7GZC/OReAK/T3O+BQn8TNwhgUdrEjDjB5MtUeAS2rbnZc3rC45zQWa6ZHTWQlpr1h61pBrUS/i
0xXxrsEok9BtadoK9weGL01HQAvaGlPVLhT+YrhDNgHP9+b+Z0XbE2xK+4NiDvPozlrKBi4rYnGu
MhgYGXgqxCEy7S6G4XksAokrDkSgIqcJUPyrXNGb53uhV1DRSdTlQbK/ZN0UJRAsKQ9rvc7ETsnp
MKMiOUMQtqeNfLLc/RKuNX6WM0yZ86iBXVVksvRl+zuRCX8ki3RHVicGdtfBLRWCP5IEys1l3Jr+
zmWioX4724jDNYdSiR7YwXy28FgKaePGf2xr2pRApZ2nzgwLTN4B07mjckhAVLLpa3wpct67kniI
DsVHFyJP90XPSVbSh6JPEB4W0uwKTpoCY5M8LBYKsX3C7uvnHYPKXp7VRFyqKKJ1LbdFCLanBnIh
rZ1yBGuyLpNbwAiuXhe36Ow3SEqEohslu5CyJ1xOFcg2hhd/DYBBSF31OuyG+OD8bToKSrldBgFl
H0bGA102rRkSnYnSCbbsloTOmFkeDTplZs1Doi2F1m971zZA+saPfYRU9jLfh0IA5QMfL/lY7NOM
FX2dKSW+HQzccCBaduODhpnXIG9bg8zFbSZL8xX4kO0+sbmWFg6RtC/HE0nLZnRTZX+tksHHdnYk
CjptoAsDE/xwtI8tk8S797VDmp5s4bU77gIVEIqDdSFBrrmWU3TuHU5K2MYeTnt3UYXbkvmvEzrK
mFEvoXIfVfnLLwjBfYKsycZTEDqgQam/eoOjgOiYQ66tw1vWVgfAuFbl/AklxNsF79K847Uu1Bi1
SLvKIMB6UeaMZF8g4LIqLePgHk8pQ2YT1z/M3Jkql2wjWVD/uoKXP6Y9eN8WZxqPmDovwos0FMzu
Dsav684s6iHuCbS2+79a1ufdMjFQo70LNk01cbBYqjbXHjhmvv8sHND2Z1WaOL7Q3jHAINkH0vPh
YUHJCq5IYq9wbIYGOBmpaZEX0Hqab4WQ+6ICIyh5PVxFY3gxXJ/VDW+kHW+J3HO4qMAxAoq+00Ad
Xjj2wsi8BJrob3pRUdW+ywhQepisiQF+PfQiKilgS9Mm1KVexU0xGQk4PnfSUSlihBrNV6W+HCYc
bKp5I2fv2NXT/sEuZfMAimcdYT5zyYAxW4pe4fXhQVGDtCKQiK+4yIqV7zVLOkLzTAlrTnkdHLlA
5quJpCh3HSokxJAaZU3cndmrkDNI+hjALrHIYw1XkUaIUGwROiOlP1uOnLEwSZL8G3ZV10adqmsO
F94yviMsVT1Z0u1Awe0rrmAZ7YWEnVFVyDTA4Xvz0TgnUB1oDWtCFeSzqUmLTWl/rOE7XODKYyQH
4FGh+t7yU9MAGOOI4xbhM1q+TMsN+p9KwAkRCntKsGnHrLxqkJlMHYTOhSOiD5R6XMm15tDhd7gw
4vWnnFOfNOebMuPc00pmDgIdEjoikMoHU7JcaHxEhWfvPdvNm04g65PkfZY2v/AwEh8LqCreN6fo
ElyUFtd82FRNNhXm75779F9f744e3QSfYqyqz42gp8PMmnNFbBRVVx7UimnSymNg2blxuIRpJjWn
Vt71ZRVh4BkCsTWSzFBO+MY73vxRRIQewPYsU6ZH0z/ga7DB5j8pofpfz1QFoWwIsxfgALNqFvH8
HKEP2Fk6yKmsZFpuEIaaaSba400O/f67pfxUA2o4KE/Ee2x0PsUpcwGgvo9gQYXnaVzmrWyy2e/3
HtuteSYrVD/H0HjzyhxDzv2/rICssnkr+gZokUAMY8itDnTmZrAjhefvBMp2vezUQzTDo84URhiA
dTR9+KARdRilmnO+vIyYXrn8/2E6wAdNr0H8DTaFSajbAqZyG362fifFtkwxoc9/eO+mvtOfzjTx
CtvlWxHUwX3XXJZCvtlqzABjtPZ3bpmbFpHDzxN+JLa7OIryIspIRf7sjfc+24FuP205ifxyl/xj
ySapDsHl7fAlA5OQKro8ap4INLk+maOptHdiSU+39KlMWB/Cq+ZHZpU3VNPtocM/PTUcSE+Jur8m
fDVf99gGIPzKapW5ZHUhKXXYfe0PxZa1MXxQqNAa5vj2Gdp6cth0o56ZdTwpcithLqkOVqUEeCl4
AGG+dq3LPSzu4fmiI4MTADj+RCyjDJqM/oXzhnxo//NUZw6QKXFFCF5+uGWCnOAag9iJrr93gYUk
6I811SpfDdWY1sGCjf6VpHYC8vdxDeWDew3whT1x8Lpaa4YJVu7D410QpEU+G2W2GRsMwcDXAgXZ
h1vRaW+YG7Bxm55QDAiGGxBqnYRruSOarZcd5rXXTaTgd98YNi7Rcb2fqphh2zjGS4zD2pDTHXPc
Ka7n2QOFMYE226LphbuTAkgrgIMZyw5Wg3O4pJGjlwm9654LlPtVXlXbWzjTmeKHsUhu/ZReefWu
/UAXFoFh9Q2ciZN7YwSDVNtzGF935MjUAxkyNz1YHIPKpQBnAKD9H2oJ/eIXnS8bc+aZEhr56maZ
EzFGR99KhlSoEob1gwE9XaIgLRzCE40uzBNHASpDmvBH12lgl75pFagAiRZe3L9J35gvGaf6QazM
qxaso/zS0gxv9e1SLgdxjBaIOraL9yzbSEluRjzWbL95LULZKzhY9tzB5Hbaz9IC8ldmri69gPMp
la4SUfkqYSiM48hAbhFDyOdozq574XpEnjk4TInlV0Kc+Of8r81QmO5cs2AZo+MAE5/e0cXYKpU1
tVQwx+lZHfHUbzH99Z3Ph9KmDcs4xw8JTnM47TFqo9gcS0VoOBnavxoZB8rSjOthNxTRv2s6yqz9
Q68RNqIcy257LvjWut0B1GFncxew1gfaPqvUQHISwoJ2uP23AXY4kAPoYwI/Ia6ps4HugMwur8rW
SAXtjJcTB0kC9B77m4K49RQZ13+dSTG69A5GXu1OQv7nC0pZxcwJX9GXofiimOpUxxnzGZlc9GIG
JQqyIAPzMmgVErfTdDSSw7QWyxG7p7tlW5tn5j3xkG1oa3+O2c++cwV+qCr0eP+wWmpw78RJl8kK
vjIfMhwMuE5yUrnMzjayX58jhywrSEXdBzpAkpCX/o1fQAUxtKYmvtzRz6fmKDWiKK5WIMe5n5pK
iv+HLU8vdswGUP1KmTbOmaBREPrNgvPFHAjab8Lh9Ihh0su1xc7G/GbwYHNCEgbLCB3Nl+/V5Suj
zVac+Aa/CIk8ogGBoBrKXcYwhsL38c3yahXH4fj2OxcVj5ctXmw4xYoLtXA2ITP9xaeCN79RemXz
7KlUAoFjOn1OGv6QRoPaIC5ntS8b3u6m3nUJBj+vRFfWuzczc2xjpCTFdsVzKLoZRub3wSlSHfc8
U1Az/qspMAON08e6CUeUUEH21aqHvgRime3JzaAJ2LdQo5bJ6suxqxYFVS98uMRNImVP3aSg4mej
zjw4gjFNHLzhR/re8I+GOdkE8pQKFtnZB11L/jmCWgFQWpTYednW/CMMnoJGqXe/h7K2IUPJYysM
vO6pG6A7n3NX5tKR5Tvxn9/ybm/xB5RSJ1KtrXWlUc2c3B2bQN/x05VedBUSdbsAYuqrEQOgU5lD
Db3ZSf8EogYgo4unGIB/LShgwcQr8QU3Ja6+r+HEg8ugUoEovhbEiE2hJ2ynHradspzUJgYfZy9E
XcDPlmk04EsXhCab62IyKUFv7yIgHmOJV0JwAcmtCfHOMZaA5b8alTs1LN0yA4lPKztyhP8mUYHO
2ohg0EJIPWAf6zvTyzBh2yw6iq3z+BzJEnKj1aHGLwrXAPtiGPodzqOedDl7eYJQ06b85YgDGlw5
WYB67qk3LBS8IVK8mEsKxOF6+RRDgo5ZJRgKbIiYk9QOzTkuSwdI3agMe1/cOp+93pIFyqUvU0wh
hqmJ8xk5jJqOLhFsN8OXIEi6Kw/NJwRw3HYY7wRv5g8sCUEQqWoU0lS3X8gRlJAOjxqHf6e9Ho4R
KF4RFmwCh4Nc9nnjPXHPISx7vywbc2yOEs8y1kQ3OF/AQ3jOTdlq+UFX89AcQL1U6BTbdEQdSPb3
uEhkKJwq11Fp/jlJ7D6yua9B0c2VKNRXEyHS8d/UboxzWOsQPBEAFEiOdSy4/YUB6Kl0woZLrfxN
KdMwaLJTIkjXsxn5MMvYJrpBxafYnMLEaoB4XB2VcdfNLcXQK9Ow7xWXNCVyP1fn+geiLkr3QocB
xVqLsGJjSfBPgo5nT9BRxUYDqoSAOPeDCfrXPgGZ18iG+lRWnYPieKhJDsePxbOnjNYELrQvukka
W8K3kOy6l00WsWq4UvuYGcTSo9Wco5KnZhW9SqHxJ2tehh46qRBVKLIhN9CxhuvYkZlhwSpnZtPK
/0+IIZFaYw4nVZg4b/j+srxTqCVQTbytcpWkYk83MOcOzVdGckxuwcYx3vke0eYKHpeLJioVXl+f
yTU/Xn9+tAVpKAEvzOk2YBDQnpaqH56WCKh3xG6G8QKpXbNj67O2DVmYekUtcsusumiD9neaiuPD
D5wMWy3TNCsThXCZPVHS6djcnqdfV+wuAVZHx9ly36n/rRcjregSi6xtx/VrN2fY4xpKcxlAIeG+
YsgkSSl7ftf7Hs84HnzAa/ZlU/KsitqWk8jyHPPbonLigz/T7PojKhV7sp2B3BbyWc4ATn0oQ6jm
/JDf7Y/Kdm3jKv+mMbAY7sIdcHVAYb4cwK8nfvaGfYiC8fSIEfi6YgOcrC1m0eyQO6wvcVjoaoNP
duIaeVLT6WE3fR5E3eUUIEerMsVWSmG/hhcRTEeU9lW6hnLVQ0sEby/e/4yT8aG3JMryQRNiyo+b
6Wa/0FLjZnqwNYlKIhBX1NP59Pz1ObYJM5LRuCYPfQEP3Gv/zhvWMPCh1zD0vSAn34Lkitt3wwER
XY7A6kBZUVKu2K8hEosK4eNH5relzGBJIWW8YtS3UBhP5wuVa4RD6YTJyqKY0gDyXsQNyXVIgOPq
r91L9OMJg1a8u+08becshJSmoaclT5n/CDSmt5qTy+lhvhmCxsB+VxrpKfyI0iliJcDkYCrDPv30
8+AXu9FxKBuFQ7XRwJmaoA8GCCrR6P52/6YPvdQ2y4ioLuKQAxqrDap6Uh7bPBj3g3sG3Jt7YNTJ
t8Mk6vA97G+iCEn7sx2UQzXGyJc5ydY0DbDXgH2+QEmCPDOxCHcVm4Bo3WSUoeBvmIXoytFAJutU
tQP05srCe9gAtNgC9LHTXXxBa62I4q8SHpwAFp2Va6NJWyVv3LrjAfWpPNTlxMCAUeBDYQNLa7na
gYlyyETmjbFdl8QBaX280sloLZF0QQzr6uJUTF+lBynfXQguUYL+2uU2EnVMl9pn3fCE4QwkI8XK
Cprjg5+nXdhHod3F4OmecBScVvs8n8h7bwd1yYtBsei5lAhtnn6p4kuKLEQ0e3dDPNtAkFP7AP4V
tOZub/RjR25gzr8bVxXhm/sUMXByQgaiA2WT6GrbcLxyhEyelvVMOCgTcxlDMCFKzhjqOh2EhiBJ
FNQkX5/2MUtqMuXugQ4SCeaV7As4otXYRakSXegMa5wrVePJV07N+v0d1K4eWRCmSOiKYSXhgtC3
LbHvX8OIyJQNQ1MCfMXdBqL+w14/BDt5M4VUD9BVM0keEP9/oifQwcgP9eYeS64R2iko2AZRSOgq
xQQviGVHVZHecODgmPRLHhMJiF+I/9FcQVtNivQhGB/D4f4/hLGJinCrXKnzAph2PBDt32H8t81U
kLaIyrsIDqQIY+mF+O9SHdvSYlkfP8WFnUKy6ak/B8MUUyWY3pQc0vXOi3rdTNGke5qDowrtyokQ
tihjmlGRDN1mUo592CEk+gKYX6GR+qElcCio+CeqBHJYqRPrTXe8M3Ar0IT0h6f6FjnanoT/d307
9n6bIZAiOzu2vLeVKCDbqqWYiN7QtH46dnnKxRYIs21jPTWVmRhuG/N5wWjG/UVQ6r2CNH5pJCWK
Vt79j65adWpVTalZkg0qL4HkhsHOEmthfLdDhHsED7dmb/83Sr2+d1mdsWVMF48B0DJGBt3bJ8dE
kIVXRPlva7PZAq+6KGbEOFO//HVu279OdIESM7KQ18jjJNiF61RiciYbo7RWMg5wrJGNe8DrGVgd
sg/OPYbMaBPLWZFH78cIM+tUinZyWiGYHGcxyUP2YVFXXg7/Jex5VDPjaoA55OaxPyjBEgMWZP0C
/ngbeEpl+t1ZFIwaiptHbS3aRGFBsRCqh53mJ/aHNvmhGZcy2h3DdRgLl5eGeTHFz0nK1gjvjzRN
nGJDHTHU6LZVm3maey4vIl5dAP4xtUQbwmJoPgL8CtnSwi4KfmTGYeZeVS08rqqsWsF8sfgXCQz0
zuA7DZJNCiBA4giEcR9PZoPyVBWpgt+q9RyKo8q2jCSe5HOx/4HBJ+rikNfuPTuckhTna2tc7R2N
qU9ba2Trb9CU4CYv+QCMSW6KXUFvtyDYhobIVN8egYD3fGrDBuVoE00BlqdHBDyXpi1LjLFDZuWu
PJVN9SwoRwzBvFH2A83hLTFuUrneR6easvwhnGJMp2XkCXnR7DHY/blD/bprWwTYC8JHr5kEb7wv
mD49aSbwuYKhvHqlcelTWjelduaDJqo3oB6a7VAwqiZZwYnKz3f6Y+HyYsmhiWmYaGiI4bMRneju
z27GmwE5lIRp+wDkPXs87qAK9qDTQjxtbqRWA4kGu3ofisUnBfwFR3zbASX7S1Vnu8Qixb6p8BzG
GHm0z6UF7qGgPXavfbgXRtbZMdiot+x7uYNdcuVbKVFzvNiHSdsC4aSvI15tIz/A8iktYiub0bvf
Bb9WsLp4ImS5Y4eY3rVNBpy8Tlwr6XfO7xfYyznCxBwjG+c98almZcm239JKFwNB2X0NXqQZ7DcH
TLd7GCe4tTiGTDrBBof8UwKT0brR9wGtPTWRUHy0DcGMfcFXGrQiGZwnah3/iLyCBCjqrAIyTYk8
ydFhl9IzXqgg4jI/bXOH+uL+k4EZ5uGyxsxvFz5Yfrl9trlaobNsnVVKO+9dLCeEscsvCjcqFZOc
JleKOAb/+CP6JScI60PLibNqp39vUAbSoKg/vD/xLO3IkqtHhO2sID6GBahnBdJIr5hC8VMWCyZq
YYv0vbzVnlgjMp6MZc20sU2ri5cF1TzTcKbd6vZdLx4SW646z4pbxWVf4BvlRsj4XYC47lQIEVMu
qOfCZVkYKwDZa/mfmHMNEUWnNbdFQ1rgLReusa8E6ol5WqVg1dm6kueQ5j8gFt/rIulaeI1r9vXY
KPdQBzqQm+4mAJ9P27ES9HeqdMLqgyME9vbOXZFK5x3HNBXvHXFTNefDyzhIDk/7Uic0OAPnZBqt
UH2EIBIVs1VJty/VYx2Abjj7f1p8OAVUxHH/bLjK9sVWb+IINhJraag60UUcO0hC7wMPUEML93PR
EjsJBbjL+W3GdZJAhpaq8C+9Xb19ntwyJaqHFQ72LGhJqEZ6n0wPSQbPgt6EOSq/y1bEvK+5IaGW
IMFtXL75qbebVHbfdfb5DbmURuoL5FhA6Q2umLMFfvYaAeImbZt74CDnhFGKhIzBifTt3NjRIBzd
NcIKNw5xMbjvrCS9b1RmuhY1czTDAzDwxSo+wFvFlIIzsRmnzVEy/sqj3U+ZXlKTbwqs8iZXLTPg
WWcykgiDpxy9+qPx/uI2XBHo3y0jOu+Y44fUkyk+CqmSDptpiPiBK8pJL9oCiHQegf+PM9AmLad4
XO2wz1G9q9vkCpqFuF0RsfIZWkV07rtlxLD8r62wHZHzw1AvCULMjGpHm+RfITYePTk0HjYG8Xhj
zw8NzGMmXX33yCEa8t0kJc87gnpilJVYrre3I0juWxuHtftPhJtRic3EWhnRWWYb8E9cyzQhWhcw
H8CL+AE11svQSXSfAO4LTvFnhlaaSy8WYLDYX/Uzq4ZXfVvgT0or7x9QQ1mCS/WdZgrpBuaRH7Um
fvnyLStGFPPO9B5t6E5EHvBp2Wx80onZoDfzlXUNREdhaHqoTzUl5BXFDbNRFCyQZBBOYv6fu9NX
ZAUFW36yPu8iPOlkzLrK5E3q7CsyXi6jhxxQd8fAHlfLbPgxenhrg5V9JLXhEZ5TSCqXPKnP7sNx
41jpb4Xn1g9VfRuI1oTplcNQVv9XSEtN8FbFmccyVkty9K31PAzreH0Jaa7VbkvubP2k3FwBK0KO
1EdmS5HWLhE7BYHEnG/HSLLkKuikSlL7wT/1RrhBDAYPzPQfwTHHxzOFrq8XfkCQq3Nmo7rDBgrw
NzPc4B4q6QMRN60Wi7PsUGN9z/9an9MZBFipZzqCHszW7C+xYqr5hUo2LVhxQJKjnyNUn73a+y/7
aJ58yNV4SzHfAkvNIWbcrQ6BWVWR53HqYZfQUzrvma3LD94dMhsclZobcezQJObFPzcxGaJIP/Rd
fvKKjOCGAWYimSXd4O4kQrTGnO5tn/r2NorIa3+VHOGLfXOvlCBjByY/ClilSUBGPyrZ9eReCFSo
FP3qeZBBEmsVkBQwMUjTBgtpDCxvOgwtwSX/DnbMH1e+SG5hmIQigDXyOXVMyvyv7cwItgmcyG5p
sqvKCpfydfVtSFfOoU1i4+umyRFI3j4hVLnC57ngiEj0TT1j/AM44vyXo3p4fX967VuE822h06yn
Iu4Klyk3GLIVbpKA6XY+qr+EwxiaLpKh/E4U1VMJaN5immCdruN/DSmDmXvnTAJFfM5ak6f6CTpf
z+UqBCezA5ul/dLp5b3gyV5RNaq6q2dkNHp5ykv+UwyIsWHyTIv5oZ9qw3qvzxxkgCsnZHlIwX/e
ewZGtNASbw9wTMUEund5yyBr4DGbA6Py95dyPj6xJQzzxv+Fwd1m2trAVbQE30p7XpbumEOyEVrz
erGnFkJUiuMgOGOlTJ9OkYoLS9kjBxvqisixArt+lAafUjJRS3mq1pr+Q5a+iIrAIYtfDvNEFCSA
MoNhDScjaExsTL/i/GJ7H3UeC99P5zEJ7iuCsDJjXbSq/Hg+W8Z5VF1c6UZdj9LEJ4wBhKaJ2fyZ
3fvKxO+P7Ziglym0friNKuifWYvBB7oyayAmCMle5BgYCZaIvOK0DCZ2nn85p/UCP/P12Zlx01Sm
GO+oZqQKhvX8SEJM/eCaDJTPQ+K2queQ4QzySvSQEBFKKmwomktfuAS6h29TkdmiTzK94RVYyaNG
zUnN2VXMB8fwJCr/liGQQvj1Gyj+MbdIda6SNAjkbRTbFfdWSAnDVX9r9SiO4yRl07Q2EoaUGLzV
a/jwimw9He87LVcbJNd/RGqHt/KuXPBvtD7IOLkwOQTpRHAFYHcmywtUfxwD1AHTTMXf15spkPow
xknDafq0WrlLYQShHy47+uaEEc6eVO41bkA+0Y5Wfhx1lf7r7OBtvYIpkQSnWCO2oKRpKdtV5bJx
vnL+NRw9GyCLQ0iQZGZWL/Akm+Pg31mE1q6ihTYxHYwNI1jR4z4xNpI0cA0iszt5hgTBX7bZ5mxs
fBQJ3Gkh60nDybA9HAxUnwDy/doPTHl6YL72ZkmnTrHsvUUcj7b0yjJVHTmTmHkMWGHV2sqsfvKd
ubhEniBXzawZg843C9W3m0XbOqNmk/0LYVBbrGSnUd/4bgPOnDn8hoKNlHr90wYWhu+VhHr1SBhI
j8l8tGFqbd5MCKK04BhFShEHIS6Zf6o6jBbkpeJqogIvYX/ZSoykyO/YoempVd44TbNYHUjXNYRm
AyJNNDE+40X74Vc4pg3Jmr5qcFLNTZ5Rr1kAUr+tVP902ZYJwTGD8+hwFfwkyX3NGxUVooUGkqLl
n88VCdIBkPdJTwk6YnUX5R5+PxmPWQHlfoJXdkGTfQxUH6JfmHUdSWzxcF7EJ99XNYyMfqIp7VU5
sVcbrhqPsE43gpMKp25x1xy7rNoe/A7Iz60Vz+/de83frZc+YknQ7ZSaIQm5xI+W21Qk6O8YlzFS
eWFU8/h7EpdgpiYKf2C1Fg27xnL8wyivVGQuPL72uEOBFHR3yGRcMfNdCvtnafqlnZO1DW2cWhyT
4vF39gQEl0e5rPX2TfwjjgH4/uxh8THj8Ps+WZesZwMupnSzsPSwa9ID+mgeGVY0HIAesZXQT/bL
7Zv+rB0nIJzdpOtUwt1A4ZpC6HKYkAhuITg+Pxl0Q+mx6WqsaMRJrqUDQ1ZslTr1N0tHcNfA3vEu
z6aYUWrObYIgHaiYpzzO1CL/N2s7fTsu7b1tLMI0Ilzo7TDoclYcWraD7gTirtPAiQ81hnEg9lg0
Kw3ixpXs+i4GIWj7oFdmdQ++yD5LSfGdKFVYGvhUXZ4qh9wFzs3mDnJH1nqyzKnMRAEKyRiarJXk
rR0gmE9Eub6cW2+UZt86lXO/O/tLxhcEmAqadDxKWoLwyslHuIeKdGAi6px5+0c0qEDVK0pSM+Sp
60xXfePxgrS6RjwnG7fUNavcQvAimImjvZkde5YhOdgWVW1fGzK1UnGRcVNA9xM6jyZ+O74RnCsj
aiJoJqAUHyKSGwGPAkvrfL3XVOx2/zAtwbbzYjP852fAI7bnUwrahZSkaBF7gIG/BO77Xn06k7SU
Lbt5l3o6FtHjq1PJRAS46IiX31yZa4FyhwJ9rkB3pZOG1VVwVRenqyS7jpKhaT5OKhmmoHOFe60P
rW3Hh5UaYpOsRs9ayurxMqDGSAxVfZulbzr62T/uEFFFAA9uUX4cAXjiAnEbBkiiAALm9ZVq8HXZ
5cz6AkXwLTRCQNMnKiSQ5+VIXIONGxJ8WBrcfXoExme811eE6hDBX0SBA/B6OwhV1qcUUC8BcwLW
LvZLpgpfMG52lS1o7IdvbcsWJ6fvaO1Mt9aYqNncNjBulE8s9XYfvUNf1j8pjhyzGNh6KMAqjQ46
BBA9q5dl0E/dYYJd/PXq4lOte+NMYTpMUkggmg7fdSG1eQzQn//pVnnl3HQ2kTQxhytqJQkwrSdp
ixf9R6QHSQ35ZvarNjwwjA/cDt7P7/8q219InMOKwrrbVjNaIxTxdURH2VD+uT3Vb8XnAnmmqzyA
nEHT/Ug4MEqSJLdkTogapBmlCSxAzzv1cg6HKbMZrls6Y+EUmtq5PaQTGJozSJeA7rkm4GUF1Geh
wqTd27fuwUn8f2z4FZNnq6nK1H9Bj72R/p0IaP0ECRopsyH2JZAozv1uzBU6jDN4BbYUqcCb59f2
zOx5xAyIlFm7ehqIrWOZK0ANY6RyHPHSyLKFo3oAGSRzz/BGrTb7k6mj5XcJOrLWntRf+QuJPBd8
wVvbl52GLbgsApAAhSMskL9vnKeDVzvSEEtsJcpd5zQ8vbmNGgDGxdIoj2WyshrsVoryZcDJXVTS
M787sxAmMuH15bsm5uOCRfBpwFUIHrZe3gPTGThEW5NuO7A0XljfmJXWHua5nNYl0s+PLqlQvSaB
Q7oJF/VFI4/byDdGNebrtRsYiwt0k5uWCupMNc2W9Vgja3mO9SskDD6vYlu+LcIQJ+LWgxToIyY0
goHYDb2NcNOnxu9r/T7HJm9WD2f86GENOZ8XJlA+OwOYz17/HgjdErcjwzd6D33OFnFM+sLv//hk
ICYqSKgJ5ZaaizB9qk3QAdjwF2pluyOwRK2LQwuF95Jb+mIroj9d9+ljxlf4upX+FydQfHIygASR
NiJaeb74ijMBPIgaFqDXomSDP0pTTu3mxOIxCN3qoxs38BfNBHGrJ5WoGbKHsLIBk3hSgxJK0Bta
BFN4eJKFSBBjoXBNjWanHagxgGvvVQ9dG9DNzHs9Oq2IkxW9KZ1RLGBjrjwdy6FibpF0azDKfCzU
1pX7kwijVeOEdyhWomPmINaSlMK57j0vczOabMLg1Nqh2h1DCNK7Y52MzmFEt9TxA/Ynx8w2dWCG
uDXbq/1U3XL8gh28ECWqrd70SRLrT+CXiGrf+7Z7kgQQytCAiuWSV6N83PAFnEQGBDasIRIKH31t
x8khdBHcdlTTWd8jNjbjiE+bzkim7MfqS0B6y3Yw+ui3rzPWG29ljHhaSN/pObeVW462CsQHZ0bP
ffxwyL638qX1O+XYF3ptdu+HB2C+AIFiul/aYnoJZr2EtcMtImPEeVCzxKU4NRu8hKMcg5/8QVE9
vsM1fpsDcIh/quodEn47HI0kYtNykOKc+Zmudeb2e9Nff4v3DqY1+KKBbFRoI2+/qUezmTgS4RHe
ZMs6PRmtYKz36EbGq/STUZPXqR+qH43GK0Z82W+jqJ/vUj5f5BJVajiX3d7nStjAlSMpjENjjQux
E80c0G2ywIFDRR9aCacd3If/kLk9JSD6Lm2s0HwBTmLsBlaYkIFvZKfDApYJc4sY9tg3h+dEKtCf
M9C46xFPxuk/FVaIS5SdZCWQpkdPV1BI7M5VAXZnCZP/0DjRKQf3B1KvEgHovdkbSVIS/Ehwe1sh
KwOI83qErIfFEE+Zg64RgOriEcULZJLXXmD2LfWa3vfqI9k3+zsL1LT1393jvWcexf0KbgNJNNBM
LSJ6qEz7V4TQStOkVJql/uPfuPzGfVWfeklK9pMIbelYx78mlQPsOCHPFzSwOTD4EQ27fdoBij8/
BlxGKe7my/uCC6mP274hBLnAoy+7ZbXPyN32FeoQhFos5Yf9s9ani8bNpNGZ8fTz8J9FbQJaGsDU
mRaqr4+8BHs/ESqc8XiwfL/9zFGx7DiK2PZhVP5sW/rCpeQj6LqRNSSGewwuhX/3INTfvUFBx3w1
o6y7F4uQHZ4wfJ4oTC8PdaJPSeLcd6pieEHf5Lhg0At4O59YlOmnaKa4kdNUoqBnpIjnG49fra3d
0AyJilzez4sSlIMBm/GbMLBCmghahufqwYaBwkFunWzMNLtzbt3iDjwkW+mRX+bBIKskKEWwZ5Ze
cSq2FZEIeQdOqjk7R+Z6f5GY1uhxTWlhqpNa3CRhG9HzceNMGe8sbJ3jNpcs+ofEFDlD9hPrRyec
zRlajDMSd9sgXlzwCG0MnZjUsrJ8Do3//IZ4Mc+4KzfaHwKmr263WrrYkx4lR2PazVXBKr+GuS32
ngJ5m6DPGBlpW3utV9XTrAYomYZnvGRNvtdk59G3AXxUVz/6L1zFaaGNnDZs8Srg4WcNXvRDBqWX
XQ+Vb0GehTFZAQ7SJs5fviQfkACCV03BIEnlQSiXe8J2R005vM9nzwri410RZ+IIGnQxF8N/ESyV
WKwMAamzDYh2FHZsNK/5+XQTCLzf73ZqW6tfPBYRX9nJHaDKgL1g20C85lETav0PhYgRd6R0dDv0
MPGZJEsA1ixJ7G/pxlMP4sx7qyo51hb+0xeOxQYCUcYxRDfKuSr16YjkxIhia/ERe2F7Bb9qpih2
N+3mLLFGxWea+VoRK3lPzM6EVRMHUxZGHMhXvq3w1OaMG+qSrN0+F3PQ3bCfIGYgZUfSf5nX4Bjx
AG3RvSD/6bDHPGRoCNzwwCPcJRPnWHRWtMpiSLaFa2pcSB8pGOktbW03DtezgSp2pEhaX6wQVq7g
KKADCF53zi2XrSmldTx3Ftav9y8ru6Oy00bRbEPgZfPyxDMwRg2jgmzSY+wvEWcXM5XyutnwqpCN
DjyXRrO9UxBSkxk8Kdbz3sMka410jeq+4QZTIrlptuyn1wo5XLcWKA77nKqY3EUtgTCrPngawLeT
oCBKwUuEn+JQInNHhJjK/1l+msIpFepPghcgWvGxV0OJOdkPi508CxUDvFTs0JCuxRGSVVcdlwk3
f7pllS/I1h59diqXFuWYa4Z60IaDpdlZavUaj6DQaoK+1/9RCcclsF9Xij/j0UOsXqmRZV+yx2UN
CR/d7XrNjgc79tD58I78BXZjqt3iiZnlIN/hzHXvAkcyqtFklUVOa1LPNhurGzR1zFVgS120j0pA
mhHBZ981sIJcgTI6jitwgULVPG3fKBnz+lrgnY2EpAGcRB20Eb/8MEuBtD/DCJfuFPGKiP7J0JJo
ApRO9LhuV68VJgAPqzZUpcSquQELn/vtVhgfdt+6YFiFh/4YUefC4dY0DFP01fVnUGMVNZqbv9Lz
gZojIP+/DIQKyRvvjDTQOHG2CMsl99MC3joJxC6vyAkpczXdg6Qd+VkGftGFEjYd0wmg9AE/3QvL
8CSPPc9vD4Bh6PvHeAg3uM1OfLoPRWK4Ye/rqTtT1w/+58C3rUj8P5cb4KP/HCZpJWgmUw/4h2VO
bHaxu/yTi0UHoipAaBwxP8XDshm3KYxjewoS5O4v3yBflFgmpDrLhVWbNTr9Ub6RQu4dRe1j4sq/
cc+bL1qOn7VG/LmvlBknSYF1vNzURBkkhW3FGgC5o5O7IiKF1jbmWVlfk4s6n5cS0nnjchS/PFkY
UEoimjUaxmUbGYbjs82Y25Bn9QZJWA2DD/sQy9bHAkhjAViVkAC1fiDYSIncx6WbskFu5IG9rMPc
XRPfbeTI2c8BSwssowNLscXKDfeA12MHGvO8w8X+33VSJrm3/KEC9SrsuxkQyybWKeXSwdrrOalE
d2KG2R77HgZi/YchjXaq1DnEY1545v7J+aAwLSyOMzuFCUiAJFnuNJQ5phF8td8kdrciK2iWpYsw
SnVGqceoXR/aJqjZWvB6df5xPM4hqqO4kEHOIANTqg94ErhD1z8Q/9Y9D9fsGviSL8DGX+wqKtBd
IRnrx7kZcRneAQTLCLjcfTnpX/xSvZYvmmBZCpBDansoFWhUJIUfnVfHtP97FMF2yUU2HNP/9XMd
7tM+lRV9qwVl8LabBkKbd8mM/vXiIBClC+rq3E0PWh1t1SzAcoNY4wBiu66VvhUy8qPZOS4omCDq
IV9Z+tHG7+VWPapdC/OUfvMwWccqcPE8GxQ8G26bj0ZyyuCPG3MCUWMgYVvQjMzj9+DAaktoQAxm
gagudbmr3pmcUmzRksp9747eMwG1rNXxThM0EIgNtPwfF1CuYwE/HsC6RfuXmrxm2iMpziGluBkD
uNou2ikhhNMM53C1mf/Q+6q2LTeaxwn/UUhIY0CM0oV5dXErrtL87o+8lFnLQGBUn2o3SKN301lM
jkrzzpu+WHNToPFmATJ/fARYn87G9/6t4sF5IJ9dgvhJWeCrS5WSh+8H4bLipLfVwNuGO/e+CgF1
mZJnhGlAHys1srDaRE//GRpbe8tt67UzY6eojZ7/txBofeQw8F55nePTR9KW4HMXrlNLg7dvV4wX
H8kypct9jxLjPzZqDcBUzseE93BAxOuVLRih/EBJ03ngGDbPz1JACe1+pCZ9RqnLa8jZCPSfb1OE
I0u7OGY7zDieNKClE450v/2f/eneXDtX6D1lcGtNK7VkmTeWK8wTyQZ26nOCILV0iyFWKC/W+g9J
ncnfbThNDnFcNz5IMuMzlxo/v88V6sCAIcvpPE0PBsfPHGPEo0serSLNJcKB8H6XagVzmcCWE1jz
2QneNvIxvPNfidO8mIrzpia1boD3rdIKs4wwoK6O7cftwCmFlt4rCGinfCeSsU4qGROn+QerSpPN
uvylgF6sxYgjL4NHQ35N9oaDa6uqKjLqLnx7eITOmC4FvkdJAkv8oqYXbBaK3ggMfSF9PEMwqYtx
KG+tsTe/d0XgblsKhREabZwBBbzsEEGH9uXmvbw7TUirdp99n1DUWz9nM8vVK69/PVMbHUvmCp+I
Gs+x0vA1MhjgerbLyYJkFsEz1C0Kdu1tNSYLUL0+z9kFm5U4SgPpxxFjqTf7K45HWXnS6dV5Cfl+
ALwQjhHEgx320h33HhCQIEGjVUBJunRxDDr1QBY+FWK54o8m4vCY6/uwPFKmxAHiYe/qOARKcgFb
UMuDB3uMyIlYuXnCOC5Jbzf5jvbuW4rblC1BWP4p9YKzpS61340RmC8dVTgm0WoIRGBAxZjZR/Yq
MLoNmofpV9C0GYrpL206JLLzaLeYf7BU4IwNMXpA2830ivJFINTUsuUUAw/QWqyvEH4lzMn6YM6F
3a++gVTg7JuntfLS02OuKZC7UoGUdfjwwaCYzoHCGr9mr1wk3QRLeFFkCU0NhQACi01SiDKdcg+P
moqIaLYSprgqASBxxQtbafP+tv9Ww4ccphsmel7E/o11WMQZCTyuixxZ/Iho8/u6ouAo7MVrgdZ/
VDmXZPSPjcZE+lb6pTNcAgZ6Ojpnx+8suJNF/XSRAtXhnMSyV2opn00rJ0e0TmTTDOblET01K3fs
GvvMXoEeeltvXI5m8PmXKXmCBNQRE5rUQdB4c/7qoj+ulyclVHk/sZWlRzLG1kbArIhRQDGDa/tD
u1b5z8h0I0zlxDJNVKI+fumx6qN+LIUJqMq34+CxsCEzKMI0O/WfS22yCWJ0UmppbFd/Bftv6Wpf
5SF5wq33DBuCpTb664Y0WEYgSR3gpfjS3oTBy+lzPtRh2Q3Rl8drxLFuA2PD0/PZgfYlpXWDyW87
yeChm+zlJ6NyUiNKlVK+qMBIH64hwBwRToVyNDAglFzMMhTAWq0Ebp+8ompLmxc9I96jxDi6Enwl
8zMHR7RCKmG4ObuWxtVy0jJpStzyF0HWO3fPSmhhrbqubhjdNUKItbMy7a02S04CfQGu5wrqAtUJ
b+saX6p4iOAyfzD+UOCCdMDmD7cqeZYGgsQTdMMmg0Z4Q+O8hcblJPfzBXMm09OA495hChgXV1jB
OF3WkqcSkjjhjQZnUDJq63YlDhyhG0nKLV+34Rtnx9Fj031mayL98tqtYCG749dVCtcjKWvkJFkz
hu5iS6p4a/Li0UiXP6yZtYnvOD50kxBzpEPNjHAjyWIU/UK0BprYw1Yujzjx1aRVSWRPrJCWWYNw
Ydzg1es68yHFWK2dPm6ot0XrGEmD4OOm4lC/A1UJbSRTZ13grww/qtYO0SmdJJwJOfpho1XMpxJS
G9AaM8jWnwhzyT5WTEaaQwlfcKZJFKWQdPxcTXgeAmTt9R3poM19C4I1Ch5a3WXW9iqVl05P3NWP
ZQMGCYEMDNe+SfyCGT2rYWPkRbg0LjYBAhiMAqq4/hcOSk7ELaSZj08Hbs0Rp5lSX3jxPl+9GGzV
g7YXXVeNpnvlSPiPTX45bbH8nwYQLAg9a2XsebAmW79/DaJwCDPfnMInwSrkQ4QDEFrtfUmpS9IU
ipwOe9Z5SDeOARlc+9tjHASxdMNOwBA0wukP1q0am7Ks0r6rE95x2Xbmnrcng+HqKrYM+dVDmANR
md//u1D7VZ8D2ID7SoDrnKWopfEsL3TtWekKisipeej6NcKg9MPdIbA2TQEDroTj4OuyfwU4pmrD
aRsSMOTnreuRu3nUX5qFXF75uMzp+gMfOLNPomnDVDL/sTHwgQ1Ak5atmNgelTKnF/lcwbM3Iiw+
lJQHGcSQKzAivmnzs6PqnYpDAX7OaI5GoQEPBh81Fch7NgNa0dDmXxB3l/8fQba6WFLgQ1BABAnG
S4hNagqr4HjUw5V8bc6aiMVIqeZtHhhxCmV+emloJ9+nrq9SyxxHYfYebG+SMqVwV9QM5oqckr2n
3C8j+S9XZH5jDSNqtyGqik3UOYA/qHkiz5yxGmhpAuL856nxz3xwsD4v4rdGKm6odorlFUvrN8qA
TkupKUhjJxi7cz+n+wMmqygSJq2KDKSiZddy73aNwmB6p1pbDUU2RgnrXQ77+PjOITaz1KcoXvOX
UiZKRFoW00YUeN/40N9Ye+VOJ4sEeUp7a1aiRkjfrErx3nuDd0YuQB+2X0Q93/dGTkbgNcrAibx1
bLYpJRX4OBHv0Jp9TXiN8LyJjfQDtErEhIZlEf824k6dUfMwQ6Eicgl1yjxDTcDo2pltQpWeyHR+
m9WtDbJflRrtdWkdzZZvIeQAhNSv8M68czYnavRLdrRBg3Uyj5ofDkfn10hCADp/tjDZ0XwYPqsJ
lw0b44LHmNMcktPn0PEsnmRoIXyJxIi7rn+hMIj67ScGvsccEcR/mVyRX/+uH8lPoDFIN2pclnpX
KlW7tycZ+9A1cIWTrGkINnv+CS80GYVU/AbLZZBin4BXUlZnXeSdbHH7vCrxt6kXhNWzhT4GLm7Q
/u89T7ca/1zG9inpXhRDVVo7CgU+FUBDzIRtc2xdlvkWZJT/ochUklNVxClO5B94kPRX+a8MpG+h
MQDDggjH6pB3+nDcljXtO1CGMAjxAjl3E1kW/iwf+i/nM4+Z1EHs/LD4Jb8xY6LyAfqdJSnvGRZS
o5kHHU8ERuwA8oI40l75qAW5UBMk1SWrqWavD5jlGTDDVH5NM8z9Q4HGHyRunNUxXQdKaJ6anK0W
BlqE5BxAtJH45W3qad3ODxRPcyRqTdsmW9jTWDFletf58QcP1r7hmeexy6jE/cpDG/fXxig3FsCv
qdSELGdI00ESIe+AvLhMCoHpDph1NkgWSNQc0IHqY7Ih0qiQXb4Vbzl7j8qtKR1zCrr4HKjRrkkO
ZP0w7X0rxYc5HwrewN+MO/c/R6kWFdQtC1plzyirfzjhBzekMdEAETcra/4dt+sHqFIVC05ZqiDi
mKrnWhcPfqgpnWS8jYBZlfZI6IKD9m2fbvMokleT3MQ5M4ma93sOezbdiJwQCIGZzrSokuB/h4bB
Mtnr3aEapzcFpO/rE2Lg0uo6TQrJ+W6iF87RwKmDdd4rEt8dxTcNlvC2Mw8e9BGLq1rT3zP5eSoK
ZAqLyM8tb0Qm7XNBKZ4RKbtjjlDTLz45BpvTow04ZGCqFReTcUiHZnZkxiYAIlyK6sSw7LsstGKi
QQ6F+6nibeupK5J8NxONGyLtNs7+M0eCQNoOu+gkylGoigI+fQU2TMXZOQEpOERxvbLi0Q8w38PV
NOKCI4UG3u5DG4x7csEbf9813cdllDHzptgELE9GYIYx3lESAksBMFhWdOi8Je/QSNckBgV+D3Q1
zKKV+ommOMlbP2kOaXkJ6mgw8PGystY5+mS76zmoLhXkA+ZlLUDugxbADbvQphtfV393R60m/JZN
zNnB6ou1yDQqVSAEz9t0MOd4VTQA0JvzhaUNk7hIaNtkjHURwWh1ulKQMw0fvA3D7QyG+EQJvc9+
PAPN5I1a3ITaMUfl1oTTltNh35OW71SQhrm7EXBUcYOV0gbIa0VfjWhxlVqClAK+VJu/WWDr33K4
6U1hul7YCFRSGXoGlyzrAyEWwQ55gE6xkjm0cC1ZpS77Uc72pzM5mGomdPhfyCaIeqOhPM+Rdw1g
vqEPq9iXlLJhAMD5DewkgYaTVaXz6Wmop6wYVFUv6X91kQ695AsfOhfq858/skGguAlTD5gFnRcz
vKYQANy+/n/MKjkS9EAq2/wAqID9iUasPZCeBUEJSfEeo144hclZjRbmEN+uuu4nA9JEh72dsbgb
fU5NoyuYWX9ho5sUmqxnpcymYDM2djj6cXCWk8pkhaIpMEm9OtQrh1nHasVVtBGRr9En1qvWUby0
khStFif3jf6yEwaclHR437UGG10n2debg72UFYlM2psKCr3PnSjeztocRJN7c9zmYPjXbS42xaAt
XrqX5Qed+G+sYdtTC/OIOZAnhQZEuxk8xQe47Q6+++zm4JyjG+V2qplpVODqdd7KN/b9SIaDiJVG
yZywOqvybBNVY7koYRhDtiTzRxk/Yx/D+dIUSJf57A6v3n1wyLU63J8Otn5sJaSXy4QGM5BgkZ/0
C0469D7MO72MkZZLEfA1YBiyfXmYTtL6frT4eYVw4dcjy+g1sw7SjJAm9L8zm07DT/i2dNHtzeQo
tKvUfxrI4HbcsGWCr4ED9h5YtM2duUYDYk8WCPOzBi/TtR3lbLesy6yy8nPNpH1aHEP/nOvh4td1
/aFo77J6sxAzGNUxUUaemOdHfD4zMq+9eWeaM0hA9iEXaq2/3VZfbs3ZZLeZmfDjszFgTAEl1+JF
SiNVOpMGvPC+HxzCwgzBoTbGas1AQT0x2j2qDTFtLK7kFjgr2w2/T6i2Cf+PZHoxxMP/7QODbXRI
O09TIhpETGzlquzcC7ZVR67NWjPMAfYhhrVkizoGAMBfHK67C52Z+FmlU9Yi3EENgAwVh/suJLvk
2uOrWFh8Q6pNCyEis2iK+Fyk3ctEyGtI7axmUX8/KLgV6caaowo/QuR/5Mwtf2GBA5tvBYEPi3Kj
Q3GQO1EPw0oYGUvRhTQF5ChJBgt4BgMcQfdfJkwxFKg7IhWT3BZz24KwEdkrrKFPV0Ei5ehaWQUc
1CoZZOCu+yf9lfSYtqD+awNysDy1ORehHCl0iook0YuwRdNOCdy+yRARY3Uv5h5f1BdDAMZu4Q7H
hcHNFN0pWPlpHpE1q5u/AXL/rsj3f5wPwjq6pbeRBko+xYa6x9tn5Ab4zp06d/MT2Cp3Bp7cPUhv
1HR9AxdKVpxTzuYUUqFLtZgOcibnYinCE467b9c0VaeJj234eSiU42Wo5LIuT63dxGPD1n0bLlse
bEW8LSYqaBLkpEbpw6n846c6fKquc5/7TgXU5vZOcRamXNK1BdzkeMS7d3elQziwFcTl8NJerIrk
3ordEkhuREyIql+4I62gsGeQCO4y6PczCt+idRaUGwolTpRy42TOkRxDXijG+DJs7wuNjBjaIaHE
nRx+EnqM+TUp6sRxsS65L9HnYZ6KC4VhV1Xfrgco78C5AM3IqPEJez2hj12II4Q+TzcjpJ1951ZT
CW4egt5j8HX88Lh9omAcueQK7dKu1p2kDNy249tYGZ3Ld+IEEE/mtQmkJyDvI7FpyIlXMk8OWjft
l8kc3INwLBBI9ezU1e59iXw9wqbBmAV/jr5ja+aajDB3dw9pe43KczQz1g+qpOX8EQ/fvS6Rou0T
JgMmeQQXkcIlcV6Te4yLSEOBoPyksp3kueDhwx0RMOljkQp+uBT2mIoWBsjElc3/fdydBpDfqhPC
tk+G5MvpCb/6izgzPrYj0ZqXKt0Xu2VMqk8wp2uj7+/IXVf2aZf6pJOQLD7yaGOHUYpNENNYLimt
4qPDXyT/egve4uCsGdu97VnGJAXJd1LIs4k7W7OGqP1/6ujlI/zI5nAsOzC1zO4ravzWyGKuTVP7
cn0m7pI6vHdw4dDqLY7CowVPsRyL3jBhb7adFT6U89PDcymrPBYtnNsyQWFwcSrEqyR6OYpbdo3j
V1o0K4OU3na9TakVUJfiHQb7SSs1K4DY31DajlMTSdluDZsFPUCI2DwgEaAMBddSHiTTCWik81NI
Io7wh0IKeeNJyoaC5FTRbiTLGc2fOGuldq5QBa3xqFlckAVkFdHEArFeFavhmUcmsTNGYM17HHIB
VHy2IjfbdXqw/xM5WA1hoMRFdpVsd662PAlo/y+VbkaaTLL/ImCeTiWQ7i1icxDugwOUWW/5PdEQ
JCbxyovpTx1knmXy6Fy72Pkm7GaJFb2drelFo6NNO8OrdEBbV6PuCP9wFWtfxJLnltmP1KgZX83x
mFpkNINcc1DDgn4Q5hB35Xd0WfXFKCXqLiNc4ZtSBxKKU7X+TD5mR9IMN6+kII3cc3D2bPiPkt6J
JHCB97jwuehIJ7wmNypD9cP6MldetAATjrCdUisdNXoqPCg66+2xugfpeNpGuYGc0jwPtWGXx7FX
aALZTSLOotSUlaFc/GcqVnygb5zCb9x3jcuXeunfbPFBIiRfSUUmHwZnHDcLyOF7moEsRsRSSYOy
WZ35XOHFHMxa3E5BL6BZGkg/8bQduFvPcl1RUDyd3ZPD6Q1ulexyq/NHGQVEnw5MPaqU77h5YdBT
piKRXt/OZr6b6Wy0pwbWicP7DljM937Ceycqe/RPCC+ydxL24pXJPscAoFmSGSD3eTf5ca8Rd+4/
cFlEw7s/aK9JPDvyeobAxE4Y4XcGd/B2N4g8wsAP2MxBsFU8ej31nZOKCFIA26zpHl5JZejjZt6P
iPbM87AekCAtM2CGJ5oN57yrHmOFnR+bLEM7YzjJNDMj06JoeC0pWBr5owY+J871WP2OV4CzRyhP
Soisg6vBN/GGKDfsM1n5H4kag9L6fL6DaX5/HDF9unw7SPfdwi6AMCzrUVw5joVZdf90g64sZ3p+
e8COxXg9fXQKjjH43rUFnFAz1Y/RnKrjugodUKuPEcjgj9ZVZoHPKwx9jc/NZ6uUWaBf44d559M0
0qC5u3lLT5PQaNJSk9I8+iGmOJDo7J9gTwo2dg0RlCStktz8tJByHB6G6A9n/hpQ++TkiUHQVGO7
kKtnuW82iZez007+xInSnhDG8olALMMCrvEzlxi/pnM551HMJLo8SwOeDBYCXQsAQWC1WC6HYg6o
qRDzWho2wuVObKHo196vd2j+Uc7uXYtacapipSdfJMDBtxvJCTfvP9i1AoMh39D62rt72q/B2ME4
G6WZ8em3hPeRxaF/mtDuIx3rQRKDZ8l55p4GAWszyUBsgXhX0wXmwTBKLB2zGKJtZ8ygkm1WHt6V
76SaKl8eAYigtYCQxUo2RsHjpwWJMiDvlL8HMhvfcb7LJhOCDaFxngcoFVwz7wsJ+b48CDOD6e3j
6Tor/7o4iAv2qRBvrsXppiulBSmk75CWCfP45gz6YQ1wIf1lMMf/GhpdN5GgXHC2gN0ePqkcs0Nz
S27EEEyLe7FynBfWVNU7yLXYlqmota5VUzgyfu/bo78U/9/ga0DVl76h8FqMYzf9DYrPBc5Ejgsq
KBldMP2wtuDnYvxtaDy2yW4dBmU/M1LsS3uZhZ7Xyxgnc0oM+NjXLF/u+/Sc/kzIlgMQNm4vVQN4
hW24TXhVNcT33yD1wHkDlXJHd3IKNKV3jXgtfWHaQmfqx3B1Q0fYYN3QlilXtkjuHy6wfrlB32Wz
fp8MY4qre3bLupc5tFnyXLtF1e5saPUexJNnrrRagWalINcGJ+PVgAICq8RlCctTbS6aErEMM7+7
TpG/sCFMRA+S04y7De/gRe4M15THoHce1Wd7batuzPF3mjV3ellBl8TdyWfB86jtTjp6Qqa2tmWR
y/CXY3BbQ4kr0bTzAxmytPdjTAw99+PVQ6/WLU0LUL8n453l6MK6vqXJ2V3lzmjpLtGIxdKt5ixc
kCkmpEft956Wx6Ptgu2GFA+xFDSrrqfGKc7RsTLU1fTmqn4iykpugpAnqmjvOMDcQRpL/vI2y7gk
RfPMImUFO7jDLQdfkpc2ayAkuTaNvn1DYcYdr282w1H0+a0s4czVqkNCdwwgZOEyI3l4/mOXoqPW
6BhCGjzdqjXDx1D2u2+I/9YcZsWrsTjAqbWNLy37g4/ZZwfY+rC4+aFALrDHsPXRdN1foATw7xWK
Y1gFsQXMRWa1rnxE7MzCqFhYTaINrf0UFGcMh+gC7o/blg3bqfUR98CSzYYveO5I+457CyyV22G/
C5be4qthHjGu8vH5Uc0LwDfsgPu0K4uUv8g+phPXqcBvsQq2ar3R3Bv1luZylZNpf50XlXKGEurm
PL6p2TBXbIELyEh2cA0UnAr6suP8UeemqImZFxWWE1vFub9ssimmEwW/8ohd+9x9Tf5qQlu7/6EP
xtzHAjXRKne9F6he0ZX0m/JUhbt7TQaeg4O5R14ulLhYl2ynn8EQjuPIEafoo9cP7ucQk6bOXo5T
qdEUkL/NBlXauk/UsHeAf8rL4Qoq8Z1sdVoGhT72NBfJC4mPZEhyiBGeGKure12Alw4Rs5405qxE
9lQdiYUxRFI3sDb4S0SlPxyonyd6NvACF/FfwWl3966foskQYRsuO0ShiOIu2Uo5phW3rOqzy75G
oGicD/slkimKfowtio0b/dWOriE1GH4FFgX4+bpXP0KcCNiX+pHJ9YBnF6GuizNM1frKtKs3fNqS
GUq/sdBNRG9oqf8C/0D8BQy42MltujPKWvUP44OnQSb4EXFuzWwnw8TTR5vk8Fd83dOkNT8ngjgh
sSUfQZ13FXx7pNC7TJCISCiVah/D7P7xIrItM+qNLCQwcbu5DiRIryhIux7DtU0nqhPhQO73m8VO
msAZ47DYahSbY8z2/OZw0FTyWJJu0y5t4M7f1zj2u2QnOWIWIfEXfJmVarSmeICNoSBWA1G/wIJw
4td9zJGA1Kk/r6urowKRih0oFuCQzyxDbJ2HcxYO83W/ImDya4OTHEb+tRZxbDnwl1ktFs/hdy2o
vJ4vMQFnQVGe7lJSV2mSAK25em8vBbUN/glypuiYee7a4FTBTg/vNi1OFl6x9yUvtjL8nEz9+wpn
1s30V0gNcUSlwOUtKD+rtwDBADbPrkAAuGyrXeuN9VOvjoFIwqmIwBfSvYOeUaNxEZ/O7H+vPTod
EkTuRZw+Uc9iogqopO9UYTpg2h+kke9la7q/M7t1CJsQoRz3eei6i0wtGAs8s9eZoJhHMDXa8Ra7
run59AzCDAHjiDMXjp40YOhAfjOvz8VhwftRhpFjd6TsZ1CqNbi6QOcY1wrmpKbvgWm/y3srYERz
8OymJuRdjrrPnc5C7ZOqqYp28NvF0+A3wIDesKjIaG7xhkV7DeVnvwytXimj0qrsJDGczdXtAtNu
6+ZniWYDDqe5xZS/0w1/CxufhdX+ncDwYa7bo1oHe/dWvBI3zd/Z2/r6/dmcsAs0VkHU5GSZW3RR
DuItG0AtkVzKKoQSXmrMGsi4pLIzk44L1c8k63yKi4RraFp+c7ADPUO3iTnY1atPnsdHYWptHxSw
drEhzJZMYdMZTYG9Ru9U0re7cAauCZTTfn9El+Wcr6qQK0Zo+ByuPrn0vnV+puRHt2bY/nR5QyHl
ycjVRR23qrKpCMhrkQeZQGJAoSMNaWdtwvF+UPvYe28mtDqFTqACaQN1JbAqICqYueEotNVGOZlM
uiqys7OXCWIs9DILnc5UKhjLx7l8nekIKWeyLmBEM3gmHdSPHX8dzh9A5IuAm2v8ZeXVOQf9/3D6
uQUlZYhbDa8m5GzEGQDzxUhGerf9/006IrtF8FzB0NZ1DurjB/ZLJdP+Q5hXkktdxwexHf0SuI0c
t/Pi5xvMw8g5lNIx/KtQw8tK8Q4JJ7kMHVd3vjCtH/cOGYIpdtPoKeZ35LBfK2PrwJv5wc8EFpkh
pOCLxnr/GAGhuwBdfz9ZF2koZfqgVSB5Z+rqkB8E8Ea1mUeJuQTW3eMBAJ2QS0Zw0FAIJYWQnIJv
XbE1ZXbgXXRJYy7eSoU2PiRvGUyhI2xuGwETnV5fGDXc0zqo5L0N8d2icv8dhJW/tEdJEruD4+DJ
yVxOYJ5uFiewnIaZ9t7FAFJioaNxdEzX1a7xSl7VlP56o0ceZ1tZM37Uy4WRAHklc36ihtzUnAde
hKZy4B8I+FDRLJYSnmgVi1NbrC8EqS/+TUeD4BEs3pbs3n4ai/TCha2JlTs6nyovUuJuCOUnNNp3
cxjRBVHyZ8migcT4UtT52WfluESmiCa05J+jmbs4ac4OZO07549LDYpx4o09dnwUs3yVcrblZnYy
/un2D6xcjcm6OKUP78c3PW9YV+0ijK8tphP8NKWQP4sxd63ctYgAW1YILIWjrmK44mzzeNG9liqU
3HFXzX+h9H3lZ+/E+E3iXPLBE2ahNbPtgYyVL7RDvQp37HUP3C95jAOqC2OhPmR9StYyxaHlxGW8
MAS9k21kdxB2VwYemq4KcnAj0tqGLrYhfdvLRw47b/F+ii5F/KugoEpoLMK4Iu9aJ7R+6ngndEZl
cZSzR6nsRPvebKSj4YzGGcIuupk45QasafYdvkCZQdbBKiVZCWSKHisOZXd3diQmX10oGu2H2kZU
uiPhPs2o8rpgfWaWfJXgf4xfm0MWb55V73ax6JMZHeHzwoaau9Yh06PyWe9w59GhEdB5hAJ9JfMx
IN+LL78g7SaGOeQWHENhOZ2yJ28e2FWcqy3Y1FAMDdZpPN23Jj8x6TOiNU2KupPukn6LGhWs7zLW
L3MvDYLtHOqrw5/HTZm4don826wYIlNnaRftMWTFGmRbWp2IDziKELV9c+/KTxab0nsjgTAtw9bl
n9BUxNBTqaOau3OmwQmlVKJ4C65tiDySzVQJ85qv3XEy7dFCAPXRY9+lBpHRRE1gkvvtzONqAj7I
jSFB4s4D4g2W0w68zJGXu6PP296Pd6PkFm0cbu2Q9abZRmLlHoxJOvGvpRqA56l/t9lDVBLFfKBL
odLCCXkXw0Bs4rMG6niapC+apyiTa2jOSdUm46mu3C66d4v8VXzdPspF8WiNv6Z26nktC7qcsm2s
HwUjye1YejGrEyWkh8j3b9E7zyJmgnGgnaJzE8u/yg/ZLo1UmldFDkkGObsoRZfvTKNX0t2j79PL
aM0btP/be5cHUFUJX8HEiGh/W1/Tl9qX8TLF98LHBeN2cKcXHjI8bLkzm9TTO2+avpa1GBKDogfl
LzrrODtha2G59NvCLUrt+THvTEAlFrxmcA9crmdh35cowUS0DbzDCsr7IKN2DyBuqFZElRNdtL9r
5QVfzq8SnfTMHqBluUMiYpjbXw2t+hAVesARbBmjnWLw2YefmGq83nHVGhe8kQWrwJh/O8EYGrKu
/RDarsyT9ZOsJthJoPZpIuYvPDp4PQwfZDiOAUWsjzrNCMOm0gH6zfQO3MfW9jhXr8tLcUdur1og
aUnv/J9tqgHxQCPC+3TxT43Sybbyg/FYRxk0rlum2a2ZCIFKLELu5ld4NSQHpRrRSl65yVMhAkPQ
hr0e2sC+C1Ccc7vC7hbpTBYv7IQzif7WUBZMw9ZPEehA9DJs30FxvbzNQm/hdBbe/Imv+drrkYVL
ovO8EUW9Ek/aL89lw5I6S3k3BC7PpVBEnNAM1ptwWmTUdWAqTjVtMk/FsJuQdu/QCc+jJnFBkV8D
uA7UqJXoaQs6l6f2EAbC3TJ04g37SZWrMxMbLwNEJfKAl9tkou8dVIcbIB3XsbQTY4kfpTS8gQ6u
PEAxeBNQuf9AxGlMCglPGcvd9R0XIkd6Hl2erxTY9g6IP2MusO8w+hIScTxxVHwbdCZKdrB4+Jat
sB4CyMEQL3DLLfHZETb44mUx5X/XaO7jO6jdWK0PNLhiFMH9C6JGiR/umopGv14v2wUFc30stadO
BqkPHC2PH85z8BPslkd6Z183y0sADF3IrWkOCnwWlOaetj4hNn2tbffQhjQd79h56+XldeSeiDdX
7yo4gUt9YbRuI2erx8Q5eJ4QJr2S+MGsd7lJMdh0/eUSTCY34+Q9T2IW2r/Jaz0Ii0zOElJp2vJ5
/26xL+Sy/J+ZTkN/WEb4LNP0u1L9JZvDyiXE3dCgXXPM1kLKNHfBAQEbrtyJEZZqhqU3V6tp8OMv
MzJXCRdDGKWx/oOqCYYaQVC/a0KSfFS7cylT2JXkRBsxIjKB5mpLRfOvHckqMJa35EGAKN15annR
vgR/XvtdJDc5t5RV98I1hxmzV1TPE4+XEPXuivhYMuGsHYar0DXB/sJr5zrNmN6duRGbW886YSDH
IpGJFAhmo066QILbQ8ITB1XoOdtbgR/3nYXx1SLsfLlzcNaikefroyuKog02zNe2oBPhM4Qp2nos
+YNlJMuVlXQkA6J/FEwzWnK2uzAY37Qukj4jQq3KoEc1Zgcpecm070I/m43e743IDWXYmO0H7waR
TuFoQcfnsw78K6KPEXk3DWrNB6iXdYAwffEipqJE3WjyMwe2PXYYG5o1jtgrT0QYXEUhln5FbsOQ
+DW7hZDDzcUT4ODXoL6grWd8Tow1tfciTQl5Uc9/gNMPP2rH/gMneJ+xU+94YMOEtbzRpGGvrL4i
ZmKccF0vS0wljwnezA3OHykD2bAhmtFySFKQfdB7dnhO8CCg9rZcPoA9bkOJ+kk+9bfTu5FU00Mo
1rKqBl6WoQia5Amk/alHoQbwWiZnkeAiu6V122IvIUPn6ky91pT1geEC6rhzDh0Upk+rtSW/pbnk
YcKvNfjUn0kMiEXho8t4/wz7Jy2s/gxuB36IrlynA1drBhuuOUgaFbyB2DdzDydUtixNQYeBgxrA
cxH6hRjrRwrF+14yA7plfe3sh6zWMy80JAhz913Yxigai9P4r8iP9UyTiTXAGkAawVCp/z9/45ag
ESXLUQRTEkYyN83h90WfOGMqPWuEnJD1p+z8IC7Ohpf+HATEGxzSP3AAwtbSyG1HKus7+21+PyYe
gszTw3oTTRczy57lja7S3wnoLAhojQJHbFc88bvPHDM1JhsedLQplmYWblgWdlZnYdJLXCBJGq7p
k7kMkCC4wTMyC1tWvg0tsI7Md0bNBVIvp+i1HoYNKDXsunXd65nXMYSD9OOqBFM7sriA8o1OdVEa
rTWRK0ParT2LBzZLXUlwPW/nhlTSkzEW638RCpN+8x9IaryL3ca5NGf4HVSKazJLFxAaXGUXcgSz
C7uhfHqA2Hbv2otU8yeuiwK8yP0JmMn/AFx75QI5l/mq8zF9uV74XB3yFwJexGy9dSfeaih1I8nQ
478PJHBqnYRdo0fokjtN7MciedCK3qOh1rIfN77xh55xhN7eaEpS08me/e3O21/ycy/Al6xeTkLg
VrZD6bHu+ztyII4YB3bBzwIYqmdHH96Kpx+Jwr1PEl30APSxEFqUHACy4wRWUuEmkCv5L9HcTLik
fra6+mptBOn9lZever7toZT/iG0Sl5qUb+mKhO3J8tIHq3EYikbespPXMyPhFgytiZEgOiBXy4iX
kfuU9pXFqlDZz6uZW2Eg3yAjtgrqDaov6dT4bIfAYs+1dNdH/nzzCGkitnfP3gCYcdB6HzxC4iQh
t7FW9iIP5EigUmsm25/iD+2aqe/EEVBMhYnuQljpRZ9IW1rFNPBKoqlVD+V3JtghNWDKw76syrem
uxv+AthRqTY5SSfTMKWxV3dbvRezVZKnAOG/tm39T2FKdYGg8Hu/xbXXcPtOrdxup80e3ueZXEWY
8uM763Wkv9O89tsZUgk9ssO85LOk2EFBSgeR7mU9H4GDNfnbYrCBB1LBhKjQoPb/bU2/HJfoXypY
t9gtzXJy/GY07eg0342Seu4leWb8tbEh6h/K5yQlotowmCY5Khvx7SauQ6nvtbKmsGFNvqfqlaYn
+NggN/mWdpR/ah1FxmWqeYNDrIEXOpuQjT0xRRg6+p1yLnYuKVJMewtZTCFD6UW+arglBHsm30JL
GNda63OTILPynmhUoalHWOg10T7aGoVLA5x/xSgGD/ws1ZTmqeKz6zj0S2BkDcwB/mBMN5pClxHm
izKO/T9wHt8gxwFnuMN7Q5FHjQEGiSbgHth7FRWc5J5HyaiWuC/lYXhtlKxTdi1HDqdQCAGcTllo
ywEGpXAnmlewhl47FqePg7mNXGP3Db2jplzYcR00S7n16Y9IIKem77eQfeTrZ5Yxf+gsURI11yB0
/pUGkdY4OEyHeWbFr+7PAc2tw6RoKYFUhgjwsFMWceC9+d8oPhvg4phawJ3Q6BYtDKXLNakGJ8Uj
TX3FxfH0xf+px/UgCbQkhfvgJvq/Bc0ELKhuOBcEkHYjTuHcYRuPCyKdenjAU0sFg/0YaE1Uf/Dg
84iuiqgpmbN0/RquwsVVLgBVyZZG3w65YmmPL3l7f+iK7m5d274YxFlwRK1daJd3y1XOuo6+b+tN
aBwDg40E2GXv+5nudyFCYpA7ghiit53PziWz8TrTQSzjh3f4MI4ullMcTDiUsL5+Mi9r6xyaV8PJ
l7lSaBoqTFygkoeu21xcD7XBXUVu9H1g3iUCqPEpa6920vGlySJMVCj+cQbpiw6Svv7yVLAH+vTb
wzBKZifZ3qRg/b4tdHebcePTRpdPrlJ8ESJrH0iy7OADLjGdL3D38ZZ5vzxGHfz7kPnnz5/KxylK
CeKvJmjrXIvxUqkRDxf5/pPYYIpIgIdVhsRkw7smtHg0lFZUbl6sdRH7Gb8YQ4CFxJ4el1Ab0dSb
S9AovUX60vKKqTeRAqYisvwcalYwiW2K4VArsoFV0ZBBKlgVbek2mDjMty8naeLvANwaf4A8asB+
6RaNBJhDzprYNGx1x65PZ66QPUixfiYhBKaOoPJNQTNXvrvmfMYDO1Rv4WbNpwrDVicdpFpHv179
/kVa9huZmDPX47p8P7p+1k7mpl9xOmBEryiATLjzA22k5qOVtwBizz/+wou37RoIDHYTwHK1FKei
xYUyF2awA0jen4D14UebKT/4eyilIwIyuIx3y71I8pHwr/BdtRRzTO7WYfVSgIkn8gXBvuPcMNTj
1BH3LY+wBVdtp5q6JMvC+QknUQMlWOmhl+azhiqZ40fc12u/RVjowgI4Rytpis5gvEZ4426MRHpK
nlj/j/+4SrCBtwvWYpz9yAQ56OO2UhgkxvmpVkObOYfVGXjE69wJz1pWvtQ4nMFwNJBPl6lGVWMq
PhOi0/N99jMgbnz/h9hwWSHxfeYpHEYJm/1yEMnIDrwVU01ya+yLPgQZLVk+SDcAEB6jwZpfr893
mMbpMQ8oSaGXuEHrmGnpL140bkVc9uOg+Dmf/NvbGtx8aLrjQOKMk4t/zEo1rdnyJuC9vYdaa1jx
RfBAHsaD/IeNCY/Mcnb68IqR1sPbFW6um1cd9AEV/1ZYxngA1res5XQhumyEw5pZtmRyHyf3tVVy
N70C6+vlq1TAjzYQnlQrntSzGdzMd0m2fI156PZm3sH0ToD7i82Qu3MHg57CjrwMudwJJlq3QlGw
e/bZDDDUKaRqIatmv0a9zuBlM/DG/rOd2l0HC3fuXS6diMfVFyjO2wqNHKuBvs9XBqJJb+ABSUIZ
WVGKK533ggLwVCSbFKa4OiLRVmyHeiU1msukSdxUH5SwRrjHtW5JmtqIEnDHu6lNzPQUOqUGhFZM
geqFecV1rwTvd3ONMWQ/Qv23KT+gwr7if7JG1vf2YQXvVmbC7ytsqJ3OzB2j/GbLh8G/U4U/7/TE
oT/+SuOgxrEE7Hk2TRji45otT1Q32xNjDBVABWxzIYmrbNp82JKvHcGUeqvA/dbU4FfQRkYh7PVh
ppL+zF/rgBIKCerywxpo0/Vhebb3WO8veEB8iboth7G7P47hMRKL/9rR77M8bNfTZfS69BPUzqa1
VFlv0YdAbbP06kMl+cVSEwFGSDNbcK1Lvb1euhzNdIm+pt7vVfWo3hhAYwO+ndSBtiG5/MTcwTf3
2bxLet0eghSr8i1VlVOrqneDAkESB9oVGrvshOTr5OWu8lYP6rj7uJqtOghpTTC7/2FLE+KKGkaK
ef2e1mEYr6eUzVLvkzU8LzTOpmjeN8IDiqL8/SnAxjdCcwwpZaidgyMuPGSIHD5qGjd5J+XYrllj
2Gbjo8+O6NtFk6N7GzaYZ+cm/OmIRR+US0W7m7QYj7Pi4RfMRAUv4NhrWV/x+C6Fk1+5i7ccvyz7
78eJUJrvJjrh646T8NCz79gtwL0E63whTeknj7xNezYn3p248aDKt9d///kGbdjTQ7yx4yaYzIHD
53J+tp4qdSjJ75MF1m0Ta++GiOA/OcBPH9sOEsTSRvG25TsM+XLf9AG/Zd7H7iT8Z9nJ1C0MohWE
iR1zJr6tMx2gw78f33qUSR0GCEbCZJmEhdmJUNIxSCX6LXl3X9aSsDbGL20p2COEd9U1cEOCtyYG
wyItP9e8oJt20GN4ZsuzLBCHeGbDbRzbafwPnzKNmjLzDHyRHQ2Zh98HdAIv/hUJ2ozdVrD/n1b6
hZii0vHD40LhqEJElhiLtXAqcwnUps3cFMuq5XpQZOLDD/vlKOEwUe7jazjpVKVJ3LkDT0I/LK5C
GQOAKBvjYB81fvj9E106XKxXRwKPULx96zM69KTnKFug/Jp+M4D0ak+5qyMVl8HUj2h0pScjDVel
OVskzO41ucB+GzSlKmy6n64d+xZJ6JxSTyv+mWyahxCvLjr8a4qtrBck6r1jV4SGF4G9zpyX5lSz
ZNzv04fIEo3u/Z3v9UhfWu+/MUgreko1px23dwhXBpMOGuAP34W0Urs0g/RTyZJ9tdp18S1807eR
A2i0dtUOkNfGkXqx0zv23JFB/9ZdHZYk47eTiUtKfnvkbHLqhBn+UwdXId1A5bZZxWFi3RV4tstM
FQlHzcp4vlLtz88jtdOEuPrEbxYNc1tOCBHLQ+nCV2/05LcMOxnVEw5dcK4mLn/qbuXXJ+TvA+2S
qyA2fG+5G5TmY/BJ2XY99Pa/6/8Q4Zc+snwUqzifVqlJR+EmigBJpm5iyk/3RRiIQnyPvZpDApz/
bTlYUvTukLlNzebFuYJs8NdxR5QeAOl16pxvlD6ch8gzLaAC5LE5k3jeIgb0Wnhgcb/wkZCpYa78
1psBlhBu1YOYG8XZEmLpxWGlPLgFCCS/bb8T2x6HvKb/MmuGq1YREDl36WWie84TOwhtY91IdLOT
ZyRd7pnCrK+daukfTEwAGqhLvhJ+bYyFOqgQgkpBYae1gG9iojvQgkugYa2smQv4g7I/O+ZPu1bw
LthUMZ4uI6xQnygG/3DxvKREk9zKhk46FKd2W2vgge0RlKPcFHgyAMhvM6/JmiDoVnEN5ooevISR
pzCWBaXBCjepVLNfSdSlG84IAh2t6tatRUyXXJHSxFO7KRX+Y0TKkTwzHXJWHf0Pzs/SJ2NRovhu
Kg9b6qgCMRCMl1ZFQ1PIgfuBUFynnxrYn3CZvAuA1zIdykEBzpUopWUVHNh500Dg2Ltt+6uZQqZs
wMTAVQGA7hFckObDT/edVgd4+fEJL9G2gkwVFf99G+F6wZuXv9M4bcC3wnYGo6YFbBzAmsko9NVI
PzEs6br1TYBgjcdF5ODr//+D4n4LhV6v9O1llLjyRzSko1iNpPPF7PyL3NNQrE/av75rSOCvX+pc
CSz3Vy19pASn8+gGJ7rcDCRl3C41gp0xzrB9gQJy9SDwtz5GrlXygWswd/teNMG+ZzDUyVEUId2N
f/0XAJbCRxSSOy4mR7oO/1x2/jm1HrzWT+gVzXT6z+tkX/zuXBRBVE2v5XRInPFsVqRaRtY40qGv
WFzGOq//YJOz2y8b2LV0kjUY2mrkf/Nzl5O/ZrtHVwDr3R/kMjVWGeIQ+/iqYO0YLD/e8m89W1TO
oE9r8snX73QKMBmvWBE86odpTqaE/CwnXd2bA2rpBid64703NI4/zwAc+BRlgAbt2xBxsgdqwgDA
pvSmis3vHeasw035d3v2bxicAQh/N1p6jKuL3d+LIxfyf0wcsjROEY9Z5A4zyA+LlsdUkX2v2mPK
RT3WQBLXLFZScUlQ+nYHQSSWJM9C2/iNKR5u/b1sQamDuWgKHjd2muXWriEeyc3Imw9X4rjDMcgn
0H3HWW6Dz1AxdUIJnUxLGPq2BTYeX1wwWXSxa+zyl3r3QAr/9BzkWz5bOpYO1dXW9iE+2VyU4ocJ
G8FiIiXYIy7j6PHDhFtXfpfgiIElz8Yzfj8Gf+JZpOgwPUxX8iDv6Y1qZ//l7Ep13lonpHR1syiz
04E603L7w6K1QAEAJVGv4URnjqSkDjrsWx2/UEFsyjTvqEs1OGz9G8GA/v/nM26TtzkOpUAUnG87
PjY2cYSCBIvAdlJN98yHYEffEZ1K38gzxQoTa7OztxlVQPUFCMiK1+wSaWcfy6pNst0ilAq7hOJW
gdBreQFN+pQ194mTahFtibI0EcNKVDw+VQFTQMAD3LvrhpgPnxkbdTuu1WSphxo7XsYYT3oLkxOL
WA2FHhWKa6ytGhH07hNk39gU5QrILOMFpIHiuEVcuWZWRelImpvSTjAjTEk07L1XRfhMnJDnRdmI
tftWxcBGqev/niSAaeWw78GhqUihEHSLpGl9xlF2YIxElxtHRdoedhOmx5jGkvi82er4oettUu5l
m+aUCwnpS12JWQ1o7Oc15pR82RHpopOgBb3vkwP5CMgTFZiIxzYxBIkULmZTPjrvDVk555EcyYJQ
2mCvMW+xmhkimEvmVZnvSLy2/FJf7HchGqDM3gBL3X4BOWh7ieYONIQdjY39bJA6V2PV/SOAWoj9
Zq154uY9cPfr13+2Q6ublTIK8R5K0ecYSF7KjBJkTDbAsEfhg3qtS2s4XRs5K0Y+pDlz6J3RLenr
OucnyI+V8zewPQNGIJGnLP8sZ7bm6ftlV6vQYX6dUPqq6zLEbgwsvbmRPbl+0qCjBBeHKN9oYQBM
CAjTMvuoyyWBIZySsX0ciFX3vqbo0Zbmbbo1/JoE3gyIV5HZaFt8RC+kkBlz9OH/FHeYJ1xH+G7U
1JUiIAcEvLgCzNeO47SFHp0OZKczSZEo4S6wcfovS/ILtudgqBX9zBjfA2SM8UM6Jypzmre68lsI
UDE+5zjKsH6SnpIsyS4FibZb/cfNNRTeK+N6a0kPqCixIrmIfSKAbUGz7Xa7dM1o91R4OO+cYDXF
dcJq58vcP+lQGYideVLk34yyJs9o8/iW9WYErWEHnD9YcJX2vIHhiyT1d01df+pF63VYfNWG8+T8
QK86mz1YGif07nxOrP8Fx/HbDrvR51e9bW4rGE4vkAkRnhVPcZQ5ITILZex4Kh3DjH/rPXyxHgzc
uIg8J4zPpqXlnXyJ2dYaeCgHBrxbpGg0zsu/vFf8jes45I8vkU1uG9uHelL8dwZlD33ACq6yrk8N
dBjBkaDVIF8z5DBjUcuPqlLRDt4fGdalIbxbB9sNQQSe5LvtyV9Y+tRdY6M8pLv5iCJu9evuYht1
f8iU0Ye8j3boCKuX0SNYunALw47vLMP+WQ3cUVzd57aoAJuYMCehhMly7QxkI8TOeLNPmZStOQIb
241g9EtAUAkL5QRZGxRjBCeCAu7qMPcvJZW7hfiE3U9jrO5fv8FEZT8gVr1A/lxYgL++k6JRBtzO
6Bs9swpmaWIvZxAUZz7/dhCOt9B7nhT2Ra0+chhoZ4x3uy1cQgiknALEh2c9lby7CGSqkHCl+6ZA
RV7+FPAP3zXQhcsWBPwd9IIqRX4KBJM1z8xDZqQmPqGuhuQaqq0zqqJDQfTXLxgyfydQWLx403Nx
Hx/rvYkvD9Ipe7FUeQLYfzsN6jV2p1bgNKJiRl8JZGk1QHJW8VOiLEndVk1+FxLjMO4+rG00+q9y
qThiFWE7bmCFNo2lyX7xpg0LQ0ZgalDRaeVyLUmv/Bxfb2vzTPYZxp8QwSroAy77jI0FI3VEk/L4
5R/GTRQT6V3KJM8h7/CQsnM4DNqGFE9FXEmb1sE5VnckqEZ76bPpkQx5YkcQHWgPYGbDpHH1YmQd
VjtK/1k0H5UtCZSaEMyolZ0V9f8PymUdRy40Uw/KV5St91k2zmWVqg+DFeA00iFIYqZi668M48y9
5CEY2Pg8S6aqArpNpTZjF2niOKJr3WvgDWDnN5JZU0ecYLW+4AHe3UVReTvNICrCfNPPJKnuq5LG
RYJO+/Pv+XeKqx75r7xJaJcCyCpUmKdfSc5Kjod9KbbH+61F9jMph9fXeDC0sUK4TKcu0w9PYB2E
4XxRuaCRBBhPgbQP4D1EtecRhz6heLuiFevdCoxLwHWjmnMhVxTHEjhm47igvJeK5w+EVeiqB2ej
L0GdcZAx+JEECKNC8NFvSjyQ0ePC25rs+PmtbEONkSs7gOmD4BXj94VYfbQaUhzLVHFM0X3CG8yX
1fuE8fYzK8L3hrf4srNE0rLZNBjpxpV0ug6csrwAjiv0LFsPLFo79Lp/vVBIiGyvXQdNnHoV+vqf
7WvPlqiXNAbZsmKZQpAQ4KKNcaTuoxEWzxY6YUEoX+V0MQ0p/BlC5dDVXfvOkTAt96SXD0vhhSpx
wK2xqmK+oN0iSk13qt6rxdT9Syyv7naXxtbJs95EoLRJYnLg1P/WNVBOjnlz0Gvx7wRF+W/0oU/j
z/K6MeH2oU5HnP1dIe3nF743LtZpMXu1ltcYSjr8n5TpCM5mXFmzlnVSxk+0y9yePt/nIhVxDIY2
duFV8MZV2F1y9iMOtc1+hRkPHFSnDc+kl9mVmZMemHArk5AmpL1NQHmbE9x6Srj42P0NXwyr1zCY
HUTHmoCsnvweLDJuKJSlSsvuwzw5jbbpZyoKqFGRLOucZJ+3S0wWUyewzLzdhlt+RS5Q0oQOhQZY
tJ6pZk788BlMK4ZvILVi3T68J54K9YCK1yE0HZJ9pM6+Ca0k1WorkvY87GNOusYC9G/1FIERIcHR
eBqdO9pIFmqxtN+aQeIiqoqLJoONh5zq/faTP9M8CPUFRyEDrRnksguX0GzM+Y0QoKAdxrtlQjTr
fIx5KOUnK91LVwO5zn/NsQ5KsvMCTqDqYemfNON6ZwFtxv1vSOWKM3KCjP3fihsZSFbUM9twDhXH
a3VQv3SFc8PPPwdFr+6CQu/x3wpGVn08N8Ma+HBBiAVyBKn+5CAKcHByrTycOZsLMCHUe6iP2Hz7
C3ZY2tEw0Yzpyr/AatHGabeCPcNkaH2eC75tKX6lF9R9Yz4f+NyV1sV92u8Eui+LmIByfrpORYbu
yTh+vPSxpzV54FMhLOw8pPIJS5prf4f5Z86FPq5Ls454RAorAWnz2/yDKB2slXZzYw6Msu5O8i/5
9BZKjGwCAUrSSk9QTGEJW4Fa3h0etCtQjUV6SF9udUwJid0jv4UYUqAteJdcaxdzQEzFLkBMVdXC
RyqegfFRajagkSV1/ptYJ+itInPI0BTgsYBCkuDxObjVGg/PLW5UF+ffuH4iJ1QztzgDBbVgt5Ml
tLBXBrIBtCMPsH5hMNelIDgVsoU3fYt8Osmrp2EnEY6+ZZ4zHer50O04aHVPoBOqwfDcNLSDTcSa
uRjy4wMq8zVuofuh8aL6SYm0AEIthJGeF25uB7Wlkz3EYQZK0/jphnAQsecHRg0MVwCIbsXHI6XZ
XQoQd2qlebYO3CiKJMk2BF8pG/pAH3cOsVFwr/hzj4WKfdePsXxlmsdOMJIxR2bYs+/hoLgvnZbO
/YAVipCu6SlB4UXLjDugLkAbfB1xTQzRJUHrY9z+T7wrrZlSbopAuTbloTsk1SExRpCIz7k9GcoS
2/o+eJk9WCa0failjwhqkbmMXT3B3MA4omMY1+YpS4NBOAoZ620YMjacxi6fBMAD9GdV11ukyNmu
QvyXQpoM13fzq4bx3EtFeD/d0k9QYKv7QAWQATha9HKTZnP2Kjjyzc8casGdr34BpW8ypquoVmS4
/GjqDmY5MsoukaaC5/2B5b0Iu5Rt9cjd7lQzsITJ5BnY/c4LRoaWgMxPxrFgaqvk1he6raNPUUfJ
t7Yz28Uhc379WmGZenEDUdmWjx6fotAXeWK9plhKtWEpkCOlJgJrHzeuDo8yJHxswlbjnjVXxmYM
hK9kqVMenZeQSVlLWHZjfjhpjPby6DIyb0iq4xsOQ4U83GgDgKTfAyLFarFtu/rMfTE0K8sc/Wnl
J/Mzf9tTSGX2/Hqg4ejs/lJhmysn9BDdvOKNwH77u7DzFdnpRevDLHnk4HejB1fhqCWHM6xZeG4j
p/ZxNHp0kvoqPh1j5HKBPEJIGhVZRxvmkWCSnRDKS3xUQm7oYhGPEzS9BS8zxcqKwJJ4wJ+5I8Rj
EKzrMNsvN18k5QWFl0wHNMc2z2UdvZ3NonoRS+0btnXhz1nLHiEyFYJbVnC4Xx1F1cPmoJgBom2T
fB5s32mSfZeuMCgfi4j1xiDEYplqxgrwLpQhA7Zg2Byb1ojbr3/qfuOhsFXlQyOM9wttut4xMolP
8osojAfpcwXQN92xZVK5n7n9iMBeDRUTdbGL2HyNv7eYD5gZzsfe4r2o72eEYzgLEdO3LKUeUThB
HrT5rb4/a8XGGaVHUHEQUcdegoNd3pHWAyrh9QTbTQuzMSfpT71KKl2HKMdNzoflmG6/SBNorbEl
F3FnXYn79wB/Mtoq6xoOc6GcV1G2XKxkdoQIuwwU418uNc93NqHOxVFcUkSgX57CNEltWdQv/+HA
tHRDI3+DIBtU/qgTeEV803jN1X5PWp7dE9JGESSGJZ+FpU22EA0xbgUBCQUQ2e/jN9aP+cGwv1FV
z5mvK1b5zgazvEXqPZLqOlyw+cS4TBcVNNmMH2O3/PO1U0Fw6LVEW0R0Ya+0PqdCgHkqXnCqw6IK
wZIfD0lYSR+7zzr/4FiLlr0JjFVeJsAMY5Zrg8Y2mfiUYKjYbPT/HSrfEwPQLeA/Hn2A+zSt5jBU
xyO4T1GPHYJjchWReyXQl8LlN8mlfJHci+lshGlz3xfEyxSkJB9TnwbU6DytbsARtDe7GKLQGhZR
5KhZjns+L3JQ5e4iSkYZ9d6N46TXLet0S+eXAIvBPsa6a4nQb9EcH1Q0lk3d0BVkGTAcpSbJOOSB
HCu8ZL4nknne7+hiG197C5cHC+lMk/7DHxdZg+RJtWKuV/x5I7VgWuT2xCIxwBEikJGe9Qcaw/5h
wazXrjPoq+msIdml4EtrWHuohKZHEbZ9f9lKesWNIvscqoJHZ0SA0z2In3D8nE7V9cLnedLZKyoY
/CrCf3r4XNTmkAVi2BkDU+6yGdfiylAnH6GkfhPkOH6I5qf+QIr1NfbZ7q+toDk6veQtBaKIe1xx
1nvGWBmRC8UkVAc8JD8OI1IjAVPfPKYS0S6mDnKre+lKA+VwkULZVo07JKtc9IA8v4+IU0i6kud9
xyZrweKTtWfbapa/W6t6HYLaWveq1+dz5Cjt28sN06EYY4HhdNKnTPhjnRzDU7P4paOjhx4mfhUo
U4K7uo5i+PiazAVvMNZUpkvkUApUKdxB5Y8qVJg9r4iQcjS+wCGlG+cgeNY2bAvFIjPMdEs0DSYT
YmM8bxp5HQ/HhSozsscWgXGtTr5qOv/LzhEmqgzM/QaS4sEEbv9tkhXvjkpkMdKupUPCQme0HjPv
yzgFs9HCthmvAmBJ6djR6hEFA2uXx/axxoS4YMOOPnG2juJUAX6hUxFSRbmQEepGh5KlPTE4bHFZ
jdB1P9+JCbO12pQ1nh9iFz5YLkI2+heoaITDhuJIYQndUcZ6laK8rurMK3dIF81AYM4B+gvx8eSu
RL45E3n7mx5zd4+d1PyGHRhtmHu6nzp+JNMokNHkFZ+YJ04AupbgbRXU3kDPeP0mGeMQU5wPPeLM
S5G+xs9Rdp732Ku/UF8K46J2lTD1sCjaXbdUoNK587N+sbfBqGEzAT6GU1WLnKKs86pIvhP++EkD
cT2s2AOa9lSv3JyRp46Of9J48cO3M3pKKYJnBP3RtivVzHrnB2FZXBNxgNLEUhzuavP2A8JxK1uI
nHmxkVB2FFX40cIpkxMdSyxc+Y34jaq1c0HeChL+XRw/sfpT8IzkyivqiObzzL5AVO2TAcwAS+5o
HyQVk7EVX91nlc6+ZXtuq38jSx+Bz/GmtqXpFmAm4mae4RKRc5TpR7BbCSrbi8+R4DLMqPSzNewg
gPBom7ytTpHdBJglnbxB8GRmDOPzQrBExUafPme9fkUwD+AM0gkNJ2yQE+8caeBNHi0gOSIIWq4O
sPqRUgRhTW/LbPWmvO4IjPjYN39tykS+0xUDqACWAscxh3f42X12BvGo29rhGM9OMdzqBL5OoF54
Y5qWgTSZ8hnXqx1GhzLLqV+SIrHcgnOjtqcgaH55rbzW0nqcqsHJ4ECRekokQyQKmzseXmzcPycT
w0MwZXdGENK/ONw/6bZ89YhyleQqDK+J3st8RSl/SpbedxLKzg4NYak9bBxe/KsYnZ7w6EAF4rJ+
8Ja5B+sc1tdL22eSyJfkStOfXtdBW/jDlUd8t25BPAD2DX2LUFLUHfjKOgz/4dy6EhMcm37I2M8G
6UF8qkLR5wqNgTJRFiN94bRI5DrL7tWoEJ3Fl8t/HquD4kpX1JH6RguU25xqKw3BBx4DNX9NtNa4
bHMeGXMt3dLkusHgM+sBIHdlkOjQdurP+nJVNTMTKqmXJOdMmXp54hl40D6gwo3to0ShGZxq3dGK
GdYpKci6mCgtNcJCuv5hmpWGAB2Pm0aWE0Gx2cjGG0aiwmEcxDYSXIOHzFtwzU6qFDPQpiDyw7IE
pTMCejy7Id2kNsm+/Bzvbc/SOd1TNE4+y6E/uxQsfbbt20tuc9FtdtUV3Yc+wsXoRqgT4rQ90qNh
92JQ1Tq2ImiqpW2spyTOgqswbpASDPKo6Jj/VOdPYMo/771ewJAtSNjOhBC21u+5PHI1HzigGJ0Z
7IOuBusNz2yXjbGb7Vnk7Z1FcsIAAsVP30G61AmuGg2U5QGfGYkOgcrVhbCWS1qcCj7z/WvNpRPi
BJJLxOVyPZU8fXEmcTaPk0MWQPJSsTP8UA0v6yEX2Ot9+HH4Wm90Yj8O9mOF9C1p9la1AygGzV2F
+MneUdvRlZtfRDJvCU9m8ktqnhlohVoYJpuaPNugVdjrw/V/zSpemSkuw4bwyFg2ctzJddAINnRR
5leU/qHbkkh3bDP+u0dfILf6kfnUGjXVoO9w2dWMPRacMS681Bq59Cubz4aHme7PdfpMgRszabD+
sItt/3PdNmuKCb+5PKnXc06TXXC9GCqJs58ejQwyJ7qol0pLP439V9Rj6Bm7VSClK+SY4lg8xcqo
IY0dJQkB03Ddn3jVGKQNli5lThzaoITzFm6agN/HLBBgkJhUDjmuucfhf/OnlXykc+T9gUtOwg9I
k4LB+6MuhAbZ6UWpA65LkjYM3yWBYQ5uZuAUj7SH40Cg7ngPYAjxBK5eI6nDMHYbREeZgLxqrdbK
bJQaDuUuWduTw3rVEe3UePk6O5YXqll8kK894pN7fIRE2W13NO1VX4sM9l+BcDypMA8t0bt6igby
zFur6LXE4/YdWJHTO58IBiXbHziB5qpnQ4ZBZ3DF5/aM6RGbmxUWP7c63V19zbRBuDxoxpASLiFU
pOKEzRX3VjXilT5ldIw8QGwaGrltSecwrrWnoZXDo/VbiQ/g4hDazWF/TuhknxoHWltkAZc50Yaa
XYuMTSMVyH4FsOtEuCGPe6EoNTcWcb15RXA4oLUaLNG1JvGN4flwfoDA/lb+ekqWBzQnAx9UkUuL
b2SZv1/M+LH4ugUxfUji1daoY9ySyAT8EAzDnsF4BFMDVumrKN3jbQijrtOREUFAyMduWOZl3IjW
rn19r9SfXk7B5SlXorErIOMF/qv/M0/oCtwiKpg7UQPh0k4evkRBuO2n+C5LzwnezMC5GzFJrbWu
zcQdH0uggq+WT1UNKhPIgnkaGg0duNAqxzjID5v0O68TT4Bwy3wfmLrDslHxvL/qK1c5hjZbOoG5
o8G/w8jEpHlXqt+KOtI1YSrmEaYdmYKxaKE1mb+HQGjgY0rR+VaUTC1SaL+Y/UL1IcB7KcLvc/qz
m2CXoVXYNLr3+TvBc5drSBQFwB2WY69WrZ66ITslGQgFXne3RcrAhooOzPZl1orkv+X7ecaVA0Xu
gBfk+aVu8iqeK7dEq/JeOPwmEB2EBtebnyfNiqoU6a5aGbe3DONAi4ZvfnuGl56l0niV3m2w/7wA
ZUq/L+RdLz3pIJsAS5Io+KrXprDWtQD480DicPnNKR6MRy7XrVotQ0aeNCkv6NCPx8sgdqIwdXfe
BkEBX+31zS7313r95cej1nhktQqV63yqoKSJ/j6M3i4Ll6H8BkPjRQD5pwozYD6wlUG0N7dt7YRT
YhmzfhkVBDYTAZ2bvy7LWEzQNNsPHR9J15UiUPmLGOY91VAaB36yRiKJYhiH6BM0Mc+e2IfDu3AE
ChFxKpYlugRDu+hOXsHOAB7/blarFu/LsePniRH3cW1WfFm3+0RQnJwDX7m9oyFZuXyBAakjzVe/
//A980zP1IxJUpZhScRFvDjAQ4CTA6RI5RUvhp928N5t/NZXswfW6L9Gk8H/PaMGjLsjo/F5oJKM
/nP/BHkFEvP8CK/Vcuewi70CM9phrlZVh0IsTpAsMuOXyQgwfo2XAOsb5ZISnQq7/BsrO1F/McLA
cuKyQ934D90TRbligZ6oUoD+fLtHg7B43WyXuqle4+6BMa+RTIP1TuQSBKfw656dbbLgJ9DMckiN
0/mXctsosIhXUrPWdHI/iXoBqyIVzXgU04F69yavVsgsq9jJdFf73ztIoBooeDTyzhstQE8AVgq/
uqHmII/R+dPK2pgjeKq4tKAL1nIefYgUh7fbIn/CHJHD2azEaeF/LQJ7CtJqPOPUXwSvjN/i0Pwe
mzPLxH396czWJmJiaLVcluxo2DhpzScNbBysGJ4rtf5Yj32nfS/b+pRcghrqV6ZdRC7FhTnwnfBY
yrFXV/C9CIUjVxxPNTx2MKg37b2q+lcnPaGPXTH0zzH1uLopA2YZ1M5drIfXftHecVZBdCjyIcLm
EWTsnJvr8SYYx+w9a4quCoHj2/vOnLssy5nYuJZaX2TsGKVaIzW8rtHibHOMfSUzJ0xwD7w90XTI
gwQk2VvUI7UcG3er2BKcvtbYV79M89uYliTZmhkaMK4xyRZqc4pMCEakmHpfXrnjgS2otigdV0EK
tNgfjI6gFhgLfJxylhOdhBtp5ejOe/pUm7lIjtBxEthN83JJk2F0ylcqSJ3talwvAbAEtHtsTBBz
u08KWJseqYABCBEUIRmgVqj/iJDXhH+O+8d+FOM0YPvRzdZ7AVYVOHj3zyHNG+h7YoDOv+aZkf78
g5RA19fp8LA7kz8C5yQxDzP/XzzxdWw1p4u1q5vZxwuPE2/Z49Lq6d4vnO87ah/FjjSo/gRwz8/X
+8ovB+4gtrOv/KFqETkwtTxCRmt16oGcLmf6XGenvc15KqEpXcUtbCYPbH/gqq8OJy1e2yrO/L+8
fkQrhXylnZSaYEJwKpAi9eoJwF5sx7o0z+yMjIVkiyBJqi+vWAAVJcpo1MniVUc7dwcyGZfzL28t
C3XGFtTHL+ysK7Dv5N9p9qZs3EfBYeWYXeTAHDxMnwnSRIA7M1uaN/or6aEB9L/nwNm0sABLQ07L
/NlzqBUZRtf9bye3puQ1JGzxwKfkvUxoW3fhVwoFJp8aFJk65CTGzqXCS/dBDz3qHT7A44BjnzQz
Eydmheegm2RE5Q0ndBYNx9ZKeMSL3J2sQQV52w/WcW1xXqyTSFyMRynHKw+hQqbiPHV+jVKNT9yf
2wP9DJF+TFk2ONmj+MsaZy+fUmaJ30Ux6xQ+DGhK0X2a7vPHzJph2p2eTtLqDCbbsiydmKolLNAp
hobk5GmFRjH7CfBXREH1mHbBIXfUgnlHSVklPTBrETPJXCf9kFXHxSTjQSw0c4tQ9s74oz8+2bT1
fSjRX4GJBmS98z4wHaTYQHCyGbmUfkm67fgxIfEaecaKmOzWiJA1lj+ExcmAemMyZM7xnckp3pYt
wtdzw/6v2TFT/eyvRzwOG5nWVQl9M2SBSMHe/PRhs6gza07KBKKRlQ4sn3M12zF7fo9h5AQbdn80
5ErMZuKhJqihALRxkC6VEQ9UI5sn5eAc7x2ebsdgf3rG0iMZ1g0nhS5haoMGKwArVEl/pQIdr+NP
+ESGZOfF5bvJdPI5FMLPIUnEcHCyLc01OqFEw8yfVoTC4RKjdofEjDMLD/lawp3SIqLmSUtzrwvj
/vJEx03V2zo2bOrqHtAFONQsHkiUVwBYXlr9w2enDW579pLaOiBMOjd0PoEj2ajCPnOm4b8H8G4e
njk7DyIXMcJnfl4Po0vn2p4KkxvbWb9wF8YN7PZtMeJxTOBEOLXvHuZRuut7prdAcbWK/DT46m2f
E+dUSVNCOilvoA90c1UxXEaaX9UCGzYV1Bh/EVqGiy9CAiI1qMpf2DqxSZmqOHuVG/ElaqYYrNTc
NLjOEJH7WePRSDwPPOcjvyz4mYZqRLoGlbCZFJKYvA0f20s7TYON+QaxrTt/moPrCu1hClDbKZWK
XYt8ibRo/3rMjOO6plTTlv3d4XbP7XRUXzHzDc1xILhXvNXoraVxB/iRrLxfcmSQ9BNV/94kiQUr
6+QloFJEYoW4loEzh9UnqKnH4cqVmTqXDt86qEDUmhxiLvu0xSaLXrSzW7j8eUsiPdx6wodFn+Gj
s2S/fJFZEGQzoxYyeoebO7xEng8s9lRj+OafXlTUNx6v0Z2stIUY8HLeek/rzCKo6S+5ijcWcin6
twoSrmlwVYTCUZmo3c2NvqS9Q2b+16nurIMDWOZQLDnZe828oN5BH6sqlLFxHMAB72o2UBBEQU92
9+QCszyEb/xBwRmf5SDQApHqZp8N6JS07cqq99E5LWqZ8yypkWSC5pL7j+T+PTz+UlmlAOLByx18
BQlkaqLl57muLu95PXGkeFUtYZuMAkf6gVJ5ogRCLjydMPWJ3AqH31LiUmrvxu43BRhbidV6A3pp
L6SbfIJeoOSjYnit8X0d2mMe/LYkFClinT3EWajU37jp8lAEzk7Fx+Jn4tZqzqEFqKCECTgHs71h
LpR0HgUgEc4cCQNK44ZwS7u8tVb9yVrBCGdJ43CsO8fY9xIGl9raznu5mhOcZlTI6h+m5cluZFxX
2otV0Sqzw+wHZEOjAFpwlMYNwoDosyi9t6MnBahjfc/Nf8FddAO5B1WXx0J8bQ9J4tnvgf4ZaPkS
r3ARtAQDfrUvnpyOKvEjknwdQtp9Qe3WaEKw4joxudWdSDyOYA9UkPTKmgd7t8UafzuSwAVFfYNw
2a/7mLjcXQ+lBLR0MXNxCBTmGPCVoC3bEqaG8kcvFsPC97hS5L7sI57tx2kB2E03dpWnCpkAGQGN
wG7q5T399XiMl3GK2aj+Vpv29YOi/c0vxhOvPAbSTZtdI4laNy6gQTlI/KGzDXa4dzTP+K5rbOHX
99yIl3TIjRH7ANnFHhz0mrBRiKxD1iwVM12W4cne1a3QpBwDwx4Wu62wa5CzcuDYBsU2ZWLw5b3H
NrFg29vD0dcGYFHTDzAlL/KVkWf6YyPhEDAdymvLhkythaqWZBf2G+rzrFAloplCb33yOJoQbex0
yO0tORrUF21xDGTV52gAL3VWeJP9GrckZH87rLc3cjqTt0HWYjLLYZPvIMsigMZWiCTEfJVtmptU
vvkwC84FquHlGiXmWHFblrCb3NcFdC5pT2F4aciKATigSw7cDrAQYe7FeCAQXvMADpBteH+jZTPI
fWc9s1di26+XzD3ShgxjkDV0T7JNONN4/IRCvVdO605+3wDTyoGlgv5f7loIPqc7WqwSXpcrWGx/
ERbVWThcyXri5sJUK27DfcJC/nrXv0O7RkgrP3GeuFfq7UOOQ2oysns/6qf8Ru3IzhP7S/BIRVZu
ZmwftkuSfjL2wQ1kxxeFhhL5g0YmA5rmeFw9FNgo+AAvYpAqPDscj+J5+FMg1X2Chf4EDPTyYq1V
z23EhIvXxqElg6dAhtw7dAwOctIQyM1e2qdkY0gzlQ3/nsg88HmRNQJ08bey6SHn0ocgzCQY58+a
zqV2i3PCJxvRSW1+haNaDhA0qTxFXDPY/A13PthFfPPYk4+ef7QGJla0R0t0NMWLxH5laQATjnMA
bF7YW1ewVvdYQxjAAUqspA0ZgA4zw3WSXpHR+VQqz3aLTKeFOPcJWloeFyM1UV/2JcYp4R1CqmF+
lh2TxV379C18tLf2+ht8gDX/YLw7b0uB2DmX+liSyJD++OEVLOi+XuL/k6CT1xZH3Oy60mjI+7uM
0ioHQEF4bCH8KoC9MRJZboap8ObF3Golot7QAdAubIVz9fZ3dsvGwUB/1X8bkRBdHvy5yb129z1z
TRxq0SkPlgcyeKh5I1zUMgFN9+ep2cv+4+lHWGYymP9JdFaxJsUQn7ytNEMp9//iR2M6R8rkQAYp
wQ6LGm+N8DWh08BgXgQQo39GAvnrVgerM+6H3Lv7oxS5bNcjFA9iiehK92DD+EMbjsVKQnxv5IRf
h+vA21/mnvTm1Xhhh6ER4oXGvFwq+RjcVR9pIXJNr6cFMI3L0zzOsplWGqhOvOBbPcKs5DavMzXx
X+MJ7PU3np9V/FpICwOZ2dnyUsv0lGYHUkMD9oFSr1K/QUORkSW6DbKg7L8p/tm+C2LkYFMykVck
xnBIrfvXN7Q2pRBDPtHDCz006dLhAVGgwV+E6HOLyWHgHfTy5dYgAqNd7lN8auA4wDVTytzFCEgf
/MwcWn/b7xQrWy+uoMIplbEKrtxAIgpBqXMaWRertR1c1LGrNlw3XDs6DI/cndt0ovDMb9svig3I
RQvXcjwKHZwhmbiEGzNN9bsoiblBcQCiindKc6MGNCAcHa2JZvpTihrrO5Q8ZE2xIMrN3ktMeFS8
+0IF95l+NHtBynUmKqSTEhNoRS4heqGk37U8YRE2FKQiEuwd6qyVzm+wM73rch2faeNAw/VP6RA+
y5ntxFHqBL+1vnbe5tJawtn41LMuj27pfji0oqcswhUgg0Vb5+7F30X6H79N8A2Y9kNk1CyRWZ5G
AbzjS0UCIz+TluoogUimbHasZRC3mQtO4aWvY7PVovTNzTzOFt5mwMIlAq5H+bh8CaonjYI1SEWf
dWygS+tqj9eQeDT9GqXthNDCpCSb2r2KUFb8p2X+Qqm2JpEBceOxM6de+GoK7L8CZ+fzMdv260wN
WtHhmWxdZEMi4LvxqTJn02l0a8DmsRdJJExC/tQWntB9+2g113TVEZxGK/juBfymdwuTqP0BkYmt
OF8vz99tZh4+7egUhlwBNAOi0YcoQ0ZynsaEOA1V+Hx4zGftMuEF2YoYopHQp55XhPeMfmgmHRh3
6G3CS/e7OS6m7F5pGI6NX2r3qb67kcHu8jXAG+z6PO0+4SvZ5s2TR962O5Dd/ZuPJljNVgL4ixCH
MmQQmwyDZzyRBhT6Ro5eXJRSE1n3k3y3mDwptLVUzeDJix1JZ43uNi8GhZS7DiI+ovxLALJqM+hU
xDOH/RoOG9uxecL3XsXk9KQ/khb4u1lsXzJqtjfhk/jAPydNFaaJCP8YTmWRMk70kBY9kf2vgfqL
9AG91TUEUtn7TB+rh8Fq202216TP0TfoY0TAAp6vevG5TSdO0AHYwuSem+jYk2NmRK8+P0s2BLH+
UET47loE1oUxKwuYcVyj3PgUZgBQEAaLa9WWXKFFY9CqR+a8vRjavjEvC/AqqGhNUNQuWAu95qJK
cHRe2QE3KtBEIp9wElYh0/IULRGK8BuIxDv/wTxHME3K2awLupvRBlXUidC/1xOueF1lh7PMNC3A
vnBu32LVqtG6jpztaUmEJn+szYO7x77IkOYwKGuwIM3Y2fFmu4qjvoKdkdVUSPdT5Ft2FMlnY3nP
0uDllJmJ3W6QkxPAa5ifjjotbNa20cV+1o0ZrEwzERpyxLSJSX+n4nIfMpu40DBMwoZAg8CizfBG
jDlx1Fzqtq8g5kSi8usDw4fw3k5cqwhEyse5NgvBHXPQYmfN3yV6mTVeNskKRNvdMAK2iFQaI8ED
oGz95a4oC2BWMsZdikUzr+wm0VfywC6dHlPWFb4ajDIyuel1C+eHrsLk+Q/Wun6MUAxE+4mDrAgt
r/m7qsUtyYSqPd7hPfIqf5hZlgv4/M1l0TvROFW/E4fHla45Hki/1WUHYiUR+R2wd8E9XVJnI1fO
sPf6YfHcFm4UsD6oR4zGiVfGnvuxl1IUr0hxN44+0xn5wmXXTydQV+/8pcK1RfN1Yrf4q3w7FLUO
ZakrRxGSJSoJlhJMmUSgpMOaUCOGRQfJigjifwjJLTrEPNv5zpCDIF2ekC6+4feJgBGpsVTRGAzR
BYwAQ0OGFYn5Yngqt+p6OldwJZCIq2KfeDKMKQRL7kkOzB/7nHxwh+DI6Az2cjX/s6NXVsCKZoTb
lX2n9OdEZv4iizzV54o3zHQnm69nlMdqGAR5ibWgU8hjPw+w8TJekp8wC2MnzLz2UNBg7KhqL+Dk
9/Z2l98AAifHN5ACs2Spt/pnBND0VzlUH/17sZCJiE/2Qi/90P6dzaNcNZ0yiUp31xFA1N3tb7V4
+Fzu1D/1xW5yO0/GfUduZqiYmIhGhSo0ujHoeMhUJe4z4IhuH2sYubiklaLNKCCkJJ5REgU04270
7mjmPNW7QDf1DPNDNBMga+iH4d76s/7rbFn56ibQKoXvPzwdzfeS3OrsHJ5U1p9N2/P08arSikp+
Crl92ps4AV8Kjaxz9F2675qwFQy0SzbpMAr4WGT7R56zKyh0XgaKPYycoiMedmAPQX81hlsk2u0O
JH48gJSxOwEHt/+jyZD43eF9vlkoQTx+E1elKTctctr1njSSawVsErHOHbjoX1LgRF2vLQBO4wLY
z5bwMYsYsfG2qfpVnMRpUX+nXe0qQTF1LkAK+iEf0VhOhZJPFbHSNbtOWUzwQIRmMtGrtctC2DX0
0ar1w7XWiJdYJRvEmBMQsZmvnB4y/OvfBM/bIZuktNqq1pacTFlL7SrUpI6S+XnqHFHL0kzOaI2p
TQ6bTphSuwyUXgz85XgOqzhtF04TlKYLcHdvn/JY65rADFTckB8nHY5+GgVswUka03y2Kbt7nLDX
rt8VwZhKE9sU3liwgjW2HTkpS7aR1QW3z2Q/glhNnn/ZFn21K8tr2sySHwb9dW+W1Z0GKmdnDfJD
WHPU3wL/41lP7+BA2VgsniSuzD4N/QqI9cnYiqKVSNEKXfTtNdJd0CwQKfrJved0jbDjDG/d6rQv
dudQx2yiNDeMxuDhVuHXi+op8Xo5+R/I+fw2CLG6s0QdpRXXIQ634FpLXwg2fNidAE1V2NIhPBPQ
mkE8p+46IFSFXDB4slM7PpJDB6NxjFI5lXbWmoMfPe9TG8Ays0C7jNMLkP4zxH/KlJiKrvbXsGGu
yHhE+9JrMS9zHdP6/H5BB4iGWIMD8ffyzTFnm38T8Z2WuZ1OIXB+9oQhVCXlgVlgveSAdQOBIF8G
1XsGr7+qlJDl3PHZSi5VXGIU0N8JcZH7hJTcGa5HGPpGNuvoUTMzX9a2TwdJMfGm4R39z6zfca5F
zlk+9NuttEbtvC4+Vm/JxMlaNSRy1WyepFg9LHzjLZutLKwhsdDEYXtXxs5dghjAQWLG6t0pJKyx
gp9QuPGOc7qdcZCqYWSUx9Eg7AmX6hxd3fBkPULf+BDR/X7zVf56SyfK6k1AWH42sjxiKSPqeQiz
m8y+LJpnIPk5lboDrW7gfD2TwJdYElx+TMLFzdyIz6vH7/DLqBh46iqzVYb/B7rg6oJDSFv/6cN3
CzxnFxmBqiG2Xp+boZx6Ce9xQ+a2zqDVpUXCBPR3QwpU0sLEPKJ+O58iIWzHV38j3JW1uCBnFA9q
UWGCBBqBS/EyL2+6wisFfGOdlb7Jf4WsYGKTJOWshW5dyerq16NzTBNSJB/lkYZpRztzunjyK59O
HfUh8C6AJZ+hJV+CuaE5iB/v1eusAlvmd5JEa6efzrRHjyJVYyokupLGbBqf9aK4noA6YTEfJOng
ppOqBtYsBW3jUyssH5he/n97zzpNZx4NHTG7PQaGydxThisW8e7CPghhizRRDg0z5cMyeoQkF9Kq
mtWHD4preTxeox6N23WdjhrK3PgR8XHBfTlhrIzHQ3Q62+kyjSKWtaJTqpoAF726rwPMkVMa09Z2
8h2+yVKSq1aSsl6hDflbdL5AUMViFMD6Ofc5sTfJTQDfR5PE/woFW/nbr6yijUxSPbA8CNx6Mo2n
5tRHIXmkQ7usApvVC7nblzLHOHtLC5JZOLjdx5ituQqCxhdWM2Q+WZbHQVp+kwZldB2wayP6oZAZ
5buKOLO4FdBAdbpCnQncGJQKZF/wrSMLphpL2C/OjvfI1xSMnGJ0cRuf1gwdOzf0wwExd9L8OOVf
7fkapsZXZrExAIDkndSOLbIFfxsWkCTutK/8eW3v+SZPxmHGx122u3dy95BNaylN2dbv/Flw5Zqs
WIqurgGFuHGt9VOptm8Br58kywn8+NRrFiV7wG12S4lYdtG/KsgomxpNYXd4UGBAAIK8BpNpVIG3
WWeKmnC8GmnwlLK+iXpydY+BjLLBU3zakK1ZaFDr0cImbdeqguApquczsGHzyzpFKxejfl0Bcavw
VPrE6fzaTNu3gVGTmCEObnD7vegpqyRInG25BmNDCSrBJRpZgXNO5oW8iI28nYJtRtevgdgMvYJf
L6EPQuspMwDzVwOMhvyFRJFgPX5vSjh5iF2SNhnHjYRSV+Vz85o6aN/o0GuG5wkkSpRCiyHEDkUG
V3TbMq8WtMfOJkg0wIIsuGxmImeAcFxE374Y5BxXA3ToG5Dcze1AkufxFUWYE6on8gt3plCo3ZsS
cC+0S448neT1NQ7d0yz9k/byAQqzhv3sdA1aOnRUEJZpVAucExFMYTN6bpPfocw2xzCOrq0HCqw5
duVKJO2aEDplh3Y84ur1UGab33RFPnNtvbv4cZXoYlRRda+QVL84oN5oyPKSN6FB921/k6stBacl
u/K+Z8Qa/QJAxPmOSk30KTtEx/MzOgHCkFZ+kSr5+crPqRIEgCNFXEDeMGTVgIfY3z3hEw2e1VL8
/hVo4YEH+HXUA8yXyWBkZAb+b9u9ZZK+lyqA5nweqVF+9URRsSTAlTu4ST9nsUxB15HQU/hUVkJO
VY7+PqcISxyJmU2446OxFE6GkW+HV73fxn6WsMUxdXM9UoaoH7NSu4n71XvujAF3bI+qtUgCpAp8
a5tCo2ZvG1sbcjM8Yx7QNAnxwr7uiuIzDGACfofw3ZVp6dvlcywTjLNC3J1LanSW5s1uDJnmREve
yHP1gVMFumNi/bPTf+hMK2deCc/HTgfl5IdYn+lGpdZNI7iTh928rhlu/+0bXuYjQQCJh21nlc7d
OMvw/CAuvSoxzUG5BlJZnb1LwwPRMSPf30mzeL2l+PDayQ2RhW4dpQDwIQ0BA+rg6CTtTV12rkLr
x5F4jgI7/uQK/W1arX5S9zIJyeYcT/B7KInqwTSKf8bm4lkFoF8TTjrCCy/PvDnhnkdJqVDVycI2
vtchy4iEmSxVs5xVQKi49Zujl6XRtyCLTF1fwPKkXwktNse/+ghdczWExw0I8ERQiJM0WeSR2ywq
Dcla7ipNRhi82LVwwqZMMf7ur448sznWaNUsylyPPzH1BWF1uEJGRVp3mCf5iI01HIXB5d4zQhVS
IeWI0ZJdfAS8LKppmMdPUdOCkaVl7adbjuDc8b+t8hXzvL314jogKn0INMDxjtYoAwfpjXk8MSlo
XSTdd/SBUSP5zSzstT3yOYZtbm9uxQNzrN8JHOXpVOrpy0MFEtjSpYdlhhnAERUhAqWCNEROfGW6
vvZWe5SvKHkXsbjG8V66edw8sTgfcaiVezVay+VOE2jXHzNo6sdec/Ew5a6WRc7W0YzBWotstL5n
u+RAK1t2p3ik9KTd+mjC11j5fv7oWXEg4ShBhKk1wnBrwKJq1LBFMhVGAs6xf09UT5NRhWmLfwar
8aCrVeiU/VE8uil+ciEjVxzi84Sm239zK0LSFe9Vf2HIBCd74n1NcDuFd6gsIJTeyovNIhUmyktM
2DW80wPpicUtCzuUoFjZ/Fvi35iJmAJF/vJs4QH7bbG6AgSBfJwCs9Xr8E2tGEYVgo6dA7My027t
ZAtCl+BBXwjQ+AGAl63AE4/iR8kCRhSes+eL83Q+8C451TEJrZ9lwDhg4iIXq795BsXHF9ybrorG
pB6jZVmIPx7IAkidLBKVXwer1Z4ZjCi6HWt9+FKRhFLVpW4qhLZKiRPu/IL0QHtQAd7o/9+HfiHB
9WSnaXywjpwqVRq6/XSe9lqUmDvouMQJu5OwKJeuO7wjBqvgysowdAsAxuRb7qPdjxm2S9qRQVUb
dcC9aL5IyuGpMdl5uFXg7CHx3xC2pTJXvXqPI3zZg27wkyr0CgJJn3vnE8DXVVL+kO2Q2DC+SB0i
hDV8W5/PDYAuEiKA2U51/owOt9gMVfYGIbyLZd5rIJFifOouwhSfIzBRDZH70lQidil/4RMCL/wN
dc3yUCpVngnGvoM0O/OQRxT9h4EgHITpmT4lDaTXndWDIJwroMAIRJL7Gv0xd9Bb0RPuOgjmqIsL
0TCsHZCREDD9jTtATiyJRYBC8o5D2XhqrH5Mi3ZEAyjIQK7nDes8J02tETqDZ95/10Ktpm0e44pK
YeaBJbLjf5E4wYOLTtrqpYqYA5z7qH2Wal/+D1picjRllzW4NMeA2jZ7zFQS79TwC5ZWjahjBbW1
kByA9mXz65Jv2D5NHLqXMECUWKIQw2sLyPH7quO2SMjbDUaF3xUKVm0lVISfJYdTBBxED6QAoVAP
8oUpWXUwkDzku7fbDApPVMOnXedwQN84qt15PjthB1+3oTnfBKNEhLcYs8qCW3YMebScMs8OPlzu
q+Fz4kKK63axebT6K+MC0XvOFi+4u0NMCm391Szt9nnqjL6J9L0u6xSBmjS9fbc8xzyl+DFIFPif
n0CM803XJk098xJ3iIT4zMCDltScKh1TuCSUN3wVMHMYS9h6Z9tlZB77ED3zw2eRXosr+4gMw8XQ
Jj1gEiVuIeDbKGEByQt2xBfGkyHHjA/PjBM9RkrD3Gyt3XlfKfST4Peu6GjX1dldoYReKpWAON86
U8Hdjt4PO1hCaorjDpVqTfIGtgLFteYuWCPe/d5H0hHRRIK8CVsMfPBtrP7EC5jA4cmsNubU01YZ
/bOH/F0ZoetOFhnyL5OAtEXjSOPN0y9KvfZcz8AzTLEJITz0mShH9g0zd/AEZankh1Og3jbvxThQ
NVjSQ2p2Uq/cAjhu159kZM6N+g2Gsi6QmA7X1XGDGNQvqlpL6b3nUCZpTrNHNJYJ3Sy0ImrI/reI
r/pVM/092N2lMmvpiGhZfUC4GRYIytlBxqkoZ5WjcmkbAEpa06yQuPhRXF/UOZa1nPTnHrTSZDY+
gSkHNOJW82WqIh5U9DmapNyIsnoKCOh1+hQlgdLIDXvkx9pELnQ1oS04ER3oE+tIvhevPtIQ7qdH
/rjpU/kg+FGCxvYiN6iDVbOaKwZycPbAQ2RMeetlKNTz/9Fw5DrFdadTFdyrYjsCm6R+slzUwKuB
BzK3DyS9EGcsGGMTvdPUnIIFK3a3IsfGfmglE53Kwim1mq0f5JQfuhjJYbPajZYo4h2o9n0+dfgQ
3FdEptUIlzyspVS9KBKZWcOky/9gRVpmi4A3uI3pbskK3CzJ877HSgv1dSjhRQXZDu+b2FFDkg8Y
Qcgv5wxTYDSC3/mYE8fMteHdOcEMV9KnxCpyQt84Q3usw2Dqn0aGMmtivrQVFnBiUwQ/tZEiu9gE
vfSMHxx1pujUC9jakxJT8gtziXoRXUYsFd8MJ+mH4YqbE0W1Yx1Y5TPQuJpwn7SLhtz+S/ztndj/
3jWfboWp070umEkcnTuRtM55svizsujsnQDrfEE78BSUUUEJis5ZmVuLnHs23IP/Rbd8foR39sAV
v5UAMBrQ8EuW1kmpgQf24exLmU5lYI2+qrgN18Kc9wYoSmI973seEOU8hw38whrNVZejDTZRIwpA
arp6Lq93ze16BL8yNOY2Z7amNolEDEvYIKiRTITgD+q/32pL4WvEuTvemHYL+oiWioYXVdVTPCtt
0eKnkmu5hDS0fT2GwMQgJ4/Q1CKKEtYiIzZZ2YX1gCBwBuMwxlxNUp5514xpUy60vhwT/g86tJTh
opQRBua0r6QEHN8xECPKAP33RO8/8mhgqGUtW9EUYbtOjuZ9dPUC1hrg0mEl5KYBnTTwHznuJgZd
WQgPo77d+gSETfpJ3P4Z1AFTFXZU0f72FjOagrRrKPx6+9TMAmVVO4ZeN22HUplO6SV/OscSuhni
87f8RH9l2yIQVlbGRdRGcY2WrSSfBNA5AJABBC8utEePg66xj3Lz1St9xgQ6++Pm8SBFDpQllybb
lmoeyMEtewlbeRZlFYDW4xn4PJBkvqqyh6T6ahAPj2IJbWmsi8c1wTRZ4Xod2PFLyuCrc18NLsHt
skzqZHiEns5W14XCyRwsl8vIo1w5kmsY9xZP2kfYs05RZJNjpQcoNPdtN2+RCsG/o2vk7LluTfy5
3bMs22V073nJpJHSrXRQXCLE1KFOZq9hGkAk4aGWM37CRVKeNbP75l699YZPJJsTBFTFrJ3eYJM0
2oU5gcNtfep+opi34NvLGQNtwEQdV1FKRAq5Q4+cZUdr8XajaZT8Ps/aLv/Amw4qm6z/IY+WUiSv
A91nDRDPb+9DypIacCoyBZZM9BaUXIds+n7d/4+WGTftXTX5A9Fsn2XBba4nCoYhu8xZBf+VjNd1
xo7QjOo7QEcNVX40Q0BH5y/oI1mNkZC+Iu8V2n+pNXyE7UZLNJh/barrebt60dAH3u9XaLxXsYo/
j9Tf9ATzSt4O+TgwgCHa+nL0jzYv8WfYogzAG4Izqy7SmIVaDiLkW+a6S7TY71KiAeI58fBrv1eL
bjc58QXxwxFsljPmPWazjWpKa3bxOCRUdsCK/tZkOm+lWF+TgXO11DidiuAmOK8MI8Rb28JBW2pA
ZDzvLzVB0hV5x/o6Lgltczg5GJ2KZa7ZcIC58SLlRZvBkIjHy/1CdPdPE39ynPirwsqQ8mMwVFjk
Yn8x7IuGRE+UK/qtpRqnU1wFWQhgeSClHXxCJavuL/djcEPbTC4ytGnmK8Do777xXTS0kg4QPbrU
54Ahqifk41E1Qp7K/es3cwzAlzsM48OFUGxgX4ZpMtJ2009LZ6Jac8hbzpdbVwKmfXr6abva5MyL
Rzee7WwaJuf7Ntl379JhRIexG2L4mfBF6AG1zkWu6p/fqvd7ZIJKkaiKo9GFplrlKYCNbbXvoY0W
raZyIZGgLadoQaUrTECgT38oRZXmdkzm8YMK3g8xGASdY/CH8v5lQNRv2C6EquAMpdfn03mQyGeK
VXSbKjEfdMI22ajXPe0nDIgjXgwS720V9zV5tGUAbX85Tb8HuqDfAMDdWE0e8xxuCH3EompEkxxZ
xiBAiP0Vb3shLtZzimmlRtookCPp+3oaliYbHjM7LvTrsiPNQylkJzfH75ko3kOBhdzzfUrDfnhW
tEF1/c59r0IWshQ6hh0lFkkamYF2q52Xzj3xy9Zm+rWfr8UwU00B6J5ZnBhnxwrZifpqbrcHqEwK
WcYxeLdoZNeBmBVAexuxIT96ZpEvmgAsTNRugC05RHFkG5wMQHqsf7gvLCgMoTUBi5hmWl61QNdL
aqqlbDgE3yoQjo2ZGVDg1+lIDHbuMm3652/roCGJqzgqukgCpP2kXgZzVqstPexBY2BiFAampOXE
IcLoSefk6zp42unr05OGE6Y60pz0AqLRgBWpNGubl/PzCDGkTRHMowxcdZsJIDLJutSXNW75eE1W
rrtmzUFoKnl8FJVB4KjHtINzhLImAp6xyBXzMlukPq67WzI+wha2SqcodHR/uT0USg4m70GiNxPp
CkAlX9B6+RilwA4aDEVJnhEwG++ojCLkkKotN0Zqoa3odc+A1dOI7+PZl9+dnuepWqf0MlngGR2B
V6zBePOH9yb+uOP5HDx0UHhPQZ0gOvbtwrhdKejF5EOYy7/is7cAHPAmA8mFxJjMh2uvng7TDypn
kwCc5w35+TJShKEQLGPotKzQvPQ+o9LstJRed2WapXmrX8aF+hUaSaMNfkTq5Wa/qEgcMAT+dQk8
sqarbzMDCxWgF2zrkEeiGyQyZ0FLdR8ZLoaUiFmKb1Enr0Ln+lxUoQ5AJnhqhLvxRMBRudmddpTv
EQaPblW0mw6CpgpT1UeQxSzpqol3fkGH8G0pPwdzMy1XkiL7xYWO4Zulp8uXwv83GUIC+aNiEpHd
3Iz8fCtHQtpbS2IKA29Iq5WkE5VGKOtgodV2ZIb0riDxsscsLQkgilFPQIiOA+rX/E5VtEQEDrSU
wTfMJ+kHjReK4vf444s44GjJu8pjL5JAcNS+6YQ8FFimQ1vXXOc3GVjVn5ea1EBcSRLNXZtY8Eyz
u3DBYplx8CP3dHqs+9jzzXTaeeAnAVntQwr1IrjVEh1VORHqYgImLAXfiUj2w6dbFhFW9UUL2wV6
sDblxSbJjRVsjc9gKAv+1YcpKbgJPmwxDJS6UX8BNyvltXkp8r1+ZUGQQ9p5SFycW8uGyB3pzGjk
6t1zYDwDxuv9p8b8n8FAeDxgvKAHX6B+MkxWUo4OS06PnlSAmLD6/l6XmA0yTvn8d9W3Z8N12qCY
Lo0WhbZxBiLI/79G+akR5aMjOfVIgpZPrIc04+2QmvpXUqbz2KxMilVkuqnVtYF+mYIxk5gNQ8e6
BIpJNlhGp3JKCgD/65TbHo/HU717VYmOWhyEyVYEFKG/LNmWdO89NTKoFunQ4yFOpQZaiKBNqMKc
1jngVFI1TYawXP2rvt8FKPc8RACmQPStRJ2Zlo5qIu7nz9cMTmm0ptPCEm+JCkzQEksJmxX5O6q9
+DCeqysmVwUO64+7oCs3DQfIkeKCC6He+ttZ7X8rg9Jg4aRNYUd6b7TLvDYXXYoGbTMsRqX7Q1QE
difv4ifTQVolqbZ1kTwE7HBwVBPFyp3sLs6xOWwQtVby6dYH/V2RQT0DiIh7xBVnz1/1H2+XUC0F
SUovN5tTUJSHNEhZ9sjWboQytQfULCYj+Gf5XSPXd4fI5YqSW9XU10WQG3AQ9aKSxinbSZ2GqIYw
KZm7lAMukeKLIvf0uX+AvusJdT/fMoq/kMa47s5WJ0KMUHJeD1jUQ3VFcdIUTeHCR1gWlW/iQKKj
dnhy24VNCPPf1Xg03xMeZdpme40wLnAXu1d1GxNj2qqMs4VdjmoGpqMx0MvFlpczPP8HY/t+y13S
kpXXKKA0z48HaneivxfmC0L0smSdNryFA1OF1mkK9Ux2qtOyeck8KAi7i9ceqzG8OD6QRoA11u2B
UDkMhDpvZ2YVwdQ6OdvhwnOEoCEPZRlZZ5pMfZ+MU5EIwlw+rN6ZC2nnj1ivK9iPR+X3fu4Faxdc
gCjw6UQS+7uAWSzDgBC2SjsC65aFuvcCS3DDvYtzPW4XTtJ0jxBuIWT20VkD7on8rTZPFBbw8sZH
gmyNsE5t1+22C5YLt8SC40J3YeFPEhl28wni0y5qFhg+KRE988kJEKPab9JJ5dwnciWsiokN0sH6
3VfT7EmNdyZjITJctWRB0Zq9cvs0FgDxjta3+dNh7RjrvyCZPK5zS8nY1/hKC/Vo7b/OzP/EVHFg
9i2RDrG2GGeFinsoJoeItjNeIXJ9/H+vUCUQeWfOll4JVKcDzAECu8r9CTQwUYE/X5QZgIbJ1LgK
XsXsDMuDO8aN1ZG97S2StvcohH7dx2lfEp7xiKdFo/8J/2myNQKpPOylWa6dpQuAkBEckHO5c2bt
4y8qZQWiIr9qifkZnopHPHV6XUD+O01eqI9tL2aoUeOU+eq5pPU3UWjqPZFJNBduxHfcRInKMYkI
N/stEpKdAQhIsGRgGdjeGdLjmA89msgsh8vjo/Way1JY+dkrT92Ut1nUR4KksBrZ/Pz9Spd30+/y
mgqSfx8UT+8CN848SBfICWiJZ1akPLozGETmAUAiOp9dp1ogDEU7vohj3Q8v+qmamUFYR8BG1yWA
Tz77z6Iy0gYb8i1n8YoKMz1SHVSljwGWPFHprM+k0W1vJGYQ1H8rpMNgnbB0RTe0kUGs42QISkB2
Bkv1gmKvuv+fr6KIa139j/1SLON1k8mlNIGUxI346UknfkM1FOy72dg8/LwXbW0rZNfbZU2vg7uX
IfEcOe51NnHtpYNCX5YYPwBGNJK4vzY6fHtRIbQ+EWSs/fNUIAu7+4UUwnVnrt5xRdTWj6Ai3Dlj
UHGKsd7OEdcwtf/YwCvLf4YbJVIX7lFTD+3aEPwKo6eMIae5FjG1AMR+KfhJoRPpXqoxVzuny2TS
ghFyHkDqvDjvvGqS5Tkd2bzqs1GHQAyW9ER2NHrQyuz0IkK9mz4I91KHuoJqMt2w2i6R9f3csaEU
dIR8C70BDe9FIdTzwae47DFhdbQmTb0Lm5TVFC2XqhSGJytoxzKz67ohcrtNrmRJ81GxeNiHAlLS
gdYXBtQF213pmoEtguzvJg4zUuIcSXgjxkLMtKSQ6laDMgiSyAPbM31MJBCbjvnw08ZyX8jiQJmn
17niFpMmcf6YJkeZY1zx009MDpsh5Eqc0ji2/SUcLkvpytwwb4kti0fhJYRYEuSJ3weSEB4mnHxm
TYlfa7DHw8KxptteRwTDe1yqZyo9DOgGi6rfjxbaz7AlodX800ZbymsqTFDJnta0BtssQ65kTqAB
JNOJNPF6PtshfLkCHLZVlz7Ca057K47ndSoMDh2DVjVX4qd+En+GBn+9UJDwBEnGYfelFCZzpc6L
YhpOQZjMD0CMvaBjsgg4CFONX55QDGbZIKhqmOEvEk9eFYV07/OFwOip+Q/56wu7IY5bRa+KxxqG
j/ukCuAZ64m134IMyHFGJKjinA70DKCi/L1tDm6T27GlKcRFrsmjZYqTH+8DFMJ4Ry6Gy5FrreOq
yGsI/S7hTlFBKPxi2P81y6FhqyDm7gr/OFlwHV+7XkR+BCw7FbJcw6Yj8fFcLlbu6gwcDzoznJz3
gucI8P6nWT5HpZ72VOaM+7umc2jjxE7p1NsItmUWfMC8SmfaBybzeY2FHMQ9+g2hfBTDr5hBjwHP
kgolHzOjyvx/cbNLRKNTGqDmlETuo7SUtRKjsATJq3/YfoujhVS7oic2giYGXgAlFvHkb9UJqgfB
RoV7l+4Mki554zffjZCwzIvknvvsq3qbmOmErY0ExcTd6X1EXd8dSdAjjDF7IRvmxrYnn3GRkmOJ
AW6tZzFyKVPFwqArD+5AJU/6FYpEn++yj74wHC2a4iNKdzkkyE+Ri1lCLgLexTHpMnioMBCBtcqs
+4uRNTedyYFCKa4mZXfMlA0wXStb9n3UfTPsxBW5O1ngzJMPuHxCqUr3SObLfdHSgGxmzQCN8cnN
jnP88bJ2KTqLg6hQ6bqkeid/v0unBtpfE7Z+0053wXtR6sbtg8kpHPiiernxzOCMaR67yisqkpdk
93v5gJtBRacPoIfMpJojG8j8oF123/toYuxFagyw8GXTJXZT+sJi7DlBo91zpbUlLTsSxqTmrene
sSEeoRZzlwkGYMVQXpFE/SHs64PknMIuh05C35P/yKdm8fPJzYFNFedaOyM8iyUt+eQarW0MDoPm
7XO97r/6QZ8SOmBJ8ccrbYyTQuKUI7+UlSxWTkncQj7l/EnMXobxtKD3uNv6Rg+lR35hkIMwbn3N
MHRBvBNyaPgJE3T3BNxdOgbsCj+++24k7bgVXY2mUADpoMME/OLhKMecGrndd+/bpuAraw5Yn44F
cdY/0LH0mHdh1UfKiVLqndoTt3ZEjUUPXD+Xq+ibzVD51ozDj5R5eq69PfPeXMmjtoa93z9QQZXE
GZ7Lb2x3NOejnuZvXWaF9ZEJ+TlImJe6nFETnkLKcSeb4sO/zADY82Npcgesi6RsWYioZN4lAugp
RtYvBuc7nschCbpQ/sbbqYV8PPaQjXkTCyG3xI/4DWXCE0LbYTCuhPABXvjWEwAwKYOb4Rk1cNan
64iyxPG6NPtwxkZiJLn9ruTYj6Nbbdw/YYuPjGsktIHzhTtyK6jZ/nOngPJ19fmbXj4JE0Yqlg8z
B6Z6o+GTUCCUyeHEkLiPdwpkZJFEz1CdmVWf4N5cC8DrKNH5tnRX0ptF+24emPKjMG+kQYjvTQKF
jGiGSJ5O2cHVstDEWlGIDDfUFoH4iWac8HTJDlr43S2KrLPyQBblVqN1P8aPfKcPnae1xYpxoFk4
BbmFwAIHFE59W2SXICpcA7P58ADx0iugTD9aMXDHZau35c1Jx3HUYfDXS9y8y3T5aQWteb/KZGAQ
GBEKE0XajrMDflkJzH3+/WF53pbY7rMF2HXGVmnAR6jWBOars42R5Afqig+rMe3E++YRlgVaqfW0
6WaZilHkQBKnenpNHtshPNSqk2jcgvQT2RIMj1STcb4jE9HmGm6j06GiVpxYgRCu4F4eenmKCo4r
fgy+zWgK4MfKT9u4/4xU2aPdDofDKoEc7EzQD9Q+UcW4l4v6Kdlcdy65SgJ+DCNV9enq+D/lHpDi
+SUZVaDtvzXtn1JMkpfXXu60F72iLgAlStdjxYbWljPwT6peyQx2BO1iyDQsfzKII/TKbTDhilTg
2jalt83usGfK6hiP02SHewZrKqW8Jy3oufDOeA7Tyzpnc/SqpYXCe23u10jPdD5QTcQNCkNyMaYi
4yCEbl9RYmuq71+YNmG2Lo/ALCst7KxSr9AiJsT+PqsTO4pa5fWFIS0rEIDM7YmB3kZJcU7pdCtS
nkX1MUltKRwVAmHM5LR2XH725dnzDSTymluZyZ67HxF0B0T6c8qs9vzRN3TDLvMVspE2351y1BcI
QQ022dyefTfV3pPABLJPKFiUBJ9Po9ha+mMHc0BhHu6IjBOpjHHEuirxTtTZ1IkGzx9ZnFrG5GK/
M2wjAx/O+mz87GVxHPnAD5pj2oe2Nj33kRFndxa673RPFL2sogkjb6Xrdp5k4sskeYOqEI2BqpFV
xqOHm7awnwJdv0vI2sbTqlkWHUtGajTxRZCg2LIaRaz+jXiSQ1X0WNS1JiH+qOg28/M0dgG/6NE8
KGDX+ruyJrKMyABgOalDpCk01FtUrnur/QonSwYffzw0xFAnPJTxLELj2a/8wlSQDXW1Vao0qFRN
iTQRzlKNLeMOvjRQulzTgjSwiX7thjgmar07cGAAh99tbrJZL9DVMR7+VUS6xndLnMhWXChB0i7q
dIvxOM7But//n76onXbsMeUA5+loUH2QNVkjlnkzgB3I9J9xE7IAHQf9MUzAlmVB9AF2M+hTbRks
wZweJ9ENIWKcAkflar5Lso+fIhleltW8WWiOxQRT8WqAQs7wJlqmYv9m8I9jALTIwG7lrEwgipd3
PF265gluAQVQgA7Pz9tB6x9gi97la1FAqxo88+sXwoxXB57hTJ3TE7d4XQM0I5/2wrbKV5wIgRTt
+u9akqLCVaGRrPJ6p6NQgIwS44qaW+ecWD/TsCfyKmITILJvBZnt8qE5up3l/yWz22qrUcXBQc6E
mqTqBp7qzTjT7ydC9uqq4VsPGFDPUtAGayOwrlsGbMAL40kOMzm2dTkyRNbWAfy8Fnoz915iAGK1
OLkIWLD3Vnolc4CGT6YtXwaMHZcITAHqdtQE51poC8AxlXxk3q9JCcHUtdWjEpc2Da3DwHNkpLNV
Cu/VQ0TpOwP5DrMd1YQf3H0NHxyOWomo9az+3KibkaTZUH307ND26/7VYZOvS7RFSQmFp9lifsAf
GYmN1O+qsGxHTViDC+O+HyzNzaXdNKK+/4s/hL8DFaeVueUcoPfbSX8azuL4paPy6XppqLW7Gt2C
Pkx3ZqW56dmwdn94z3Tyx/F5XEIsoPXCCDRgQV4O9aK8X8hldZGozmC52HCbGAEuKF8YfLpS3m6r
nQx3E7ZjzGy5gyoD7nEuIRW66kuA3AeW8EB7IineNVtPHq3vznEUxzPw1z6DgmHhXGaA+22nKG0L
WZ468SFua/eF0t3hayXJatCO5rQD+3mCl0I0BzN/zzCeBZ6KyqcBSKSssYBPqZH2jkUhUn/ME74W
jYZuit8thYEz0kAa2TyKOBPD+CX/1+zcz0UO4Jg3s2ZgwERxUxTzqhZt2pJobg8xQfM/b1Z9eibI
icCLtIhHqLSPEk80YN1huKgskB473Qx1HswcSoapEyBvDROgJ3riPaswrPyANdjm5cpj35CMZSKx
gCTEVF6UQz7oTKLV/K1+gURjPWZk0ZSghdMBL6VV7n+tG6vwGIyEHbgodrJlQBv2xbdCFOuIvoqS
64S/WvguBW4shqtBWa6y3FyxxHQNraPDlInDDDgZ0R2LrYK5LNcBljfK4dC72IZiheE9BKNUnGxt
bBQWDK9zKi/rpAPBE+WL96mJzwQqIG5m+nrVidnShmY5HVvMd/rnCDDTwHRYn7ef8E9oW8GxW4+6
sgTt85VZW45kef0VtUQn9t9rJuncHqVGtrsWdwWnqXxcnVfnOl5p/Q3mLqan1xalF7KcVqDztoit
xEmTEAzCIHZc4724pO8v6jKvOnxEh5RVmaF6wcCDcoWSEfdkkS8fdFc8WTV9kXq6dM8MFWtAhBcd
I9zO154RBfNoBlDEZqYnr0SfSTHktSKEKztNn/QvrXl8PZFnmX5oR4bL/wG3uMF5Za59K9pAMt7N
ZJfPaQOrrPCFrh7HjqRAwEyPANzSCtUUFGRHWC/Y3uT65EvIOOlHBaot5MYp6mfR28Nlcd0xceVL
Ftj52Jnx7AjTZVzqQN+cv44SQHCBUfEiCAAqZLIeOSNXjnWfBWZDsjr7E1UeyuSCjEO+OScBWdBy
PsWTlnVk6cWXwp8+wW11Uh58KHiQXt70Q/IeuxK5yS+nPmzv3X8+edIoK+iQZBxryWUYk1gYpVi9
gEqtsQ0xnFsSu6wCJFIWQNfknU15QdQgdKt8D8g98gSWUIIXlJzr4aEmSgcplaRkPJJgudlj19qv
6+MC0zD6/hCaLc0DuYcDFWN8LwH4v4nKYoc1S/DnJiNpEv4F3LFZxUM7pIAMzCDgaQfP6bhyiLjs
X6qeUx+I6E+Qve34s+8yvXo+f9Lbke87nFM/KIMxhZrupSI5kpFmsiZGJWCZYcfaUOfk+0BE7nym
ARwjo7zECAi8P7LthHAs08+/EDtMg04vGaIYWcAJpymPhgU6B9OSqG4OcJASyD/J93uJauCaqLoW
trRwHgAZT670XWQF9qU2WMULQknUepFRCdwKAUfrrRqEXpxC6QxqWbIB/Nd6hFpF3/ci9/6zuyG7
krAQPBReahDARgBoAvK9sY1Ga4aYraTTadQssgMU/hFNHXKG+R5cmlVhjWt2YKVn3UTiF6RkjSWY
F5VC/x+QvDHT+VJM1KpJJ79hvBsjbYPQjQTPE7gN3/Ikd2NM+otY8fqKoPhsIVs5AnzGgqNoZfgO
aKrsYVUOSdw44dJ7L663aFi/rijEo5rCliiCbLt/T78/0kJJ/5aXE22nIl0cXogcVGWIjsGIBOlC
G1MaUUtMY4RgFEfwXU6XQCwyewD07yUfbvbe48A3i49FbTW0Ozr5BgYSIbWAOpqDBP35e8u0lpPx
Rx9aZSj1tmxgU2Tz0IPKw3rUM3y6a2o7EZkpxxhCZHagnnO4c/IonV7dXe+PIlZkONJnJIiLl289
5sJZNbEI0R8SYrSZtMPAiCtyTMYQdprE6Baq8pBtR9XKGxMzzRiXO5hLbYqKz6/3+tsF2iCr/Fb6
sl5yPe5xcNxSjk8cBqoNRF5l9FA/qyZJ/zLXv4nWPaTypc4Tf3QVz0dbLeFPm9RLijH6RiNafG5h
nTI+INN3KkorryCfQr1reoQKf92ojSrpjUMiknNNBF+Su8DC8hmwtBuoLaKe8KrxFceiEQ7No8cB
r2+DTvLZKEvJ6rSH3lji+WuoK/Psnh6VWejK9qSwYKIBoKxykeYwa2XA+s0HEADSG1mbCFKb6Rb/
IIWWbjXxVEYRd6ST7lLtmnYR8h1Xab6dA92KRsVKa2YjuXkXwBDnnHWr0RjCk3fC2yEKjX2J5Ns3
si/pxrvhmAl7WMx7sgJ03NOzdBbixn+a3XsKfc3dpkbDtVOcv7/H4J3YGEsbKExYx/kN0/qBzWfT
lKtjwOzW43xCu+r8ttT8CptdRcfa45oXAghBTiqfm7hSk5M2LkiJPj1HmyNDlh8aqG6XcGvnbxC5
JomlNReTj4KyM9n20k+lOWoOkoLeIrTB8NThZBcfCXoaxkKhOKX48X/91T0AuqKMRm5RSy2wdqqY
snyuf6BiBGf7RiV2ENEjZJo0GZZpIlCTA0XltG7BYcMjdt1F5sQ57lIEYRdLLAaelB8iuu6Vg+X8
Y2CrsIcEzkAFQajAavU3OxfOFonZAtp+Y+9k0u8BD/RTrkCge+oBdGYazIkcX7JhA/IGpiMhdB9/
7xD3t4O0MT25nmzsH39JbMKB7TSQu+slZchkzNnhCe+qDaQAp+UsBgTa4LDNuooP2lX4gZJf8PGu
b3hkWWkV5RwcPjWqKEMfeFR2CdComP9HEJVjWZ4EWWxZF6M32GuyBF+xhTbykEzLvRK/S2SvO6LC
KezGJlaM3u8dB4scUN1SuKGextynKKgvcNhORP+TK3QJFMnUXmPPo99HCzF8SE2Lbpx2AJJNJpGc
7Ay8ar4W7royOoPtoBHXVWJOyESJ+FTwrVMYS6wVNYbBj0kN0urF2lNOd/mxqqrEFIMaWvcjnVrc
XI2g+s3SrO5WsgiHg3L/dSgOs95Amfd31T/jj8L/C9RU5X4967mOdvPuU3BNAZQFj73IeWNUjc6K
aaPhnPcnETPRCgRks3urxIHBMgqVZfKeg0ECbk5Op+S/xVVBHv0R2Iyk9kLcufPS9VhglbghvAno
qJ5XaQcysSOigAqCfjH11IOjBcYvvKj2qUv9co7hAWAH8IdFC41rWcIOSZHoLdJsbbk0kzQhQCpq
zHmJpHJyxJvHy3TtlQtisgXl0hK2aDBRgg3kuIVtxTF5/mM+usEMyLwyn/h2epzKKA7FRKVPsce8
TOTcKWZFKtbFR4tdgy10riRDQ3sjrlX3NFb0W/NmgwmQvdbuqUEPaskVEjSTgKxhnDaOR3MkIFLa
QRvwWOSfBHF3I/7AEf9t0CdMeqkRtIFR2V9mWVOoApyKfyVJ46TUzT2OKlZW398V0uOmVvJDSX/e
HPM26XuOf78mZBxFJWW0s0tuGsqOiTur0ngJXVGqzD5ORCUsciBoWtDnpPjGxOmKuGMWPRrb54RM
Z/Xefhm3MOeWfIzUhwl5q7TYFxSWrJcvuiBjP1Yg6xTe5JMVU0PklscytcWlniFKpeJFJ/yCA/w6
y9N0yqNDQ8WKANO2HIq9fSm1E9w7c3awx+Iw2JWsDz86ZrhzLu63HcbaaOKeuYKkEMXXNOJpDRTF
DOpL7pIuVIHhhItyujf2WsmwWEZDQSLOrCs0g4Kg+bkLMjxDLUfV3lbUQt/WrbQHSzIB+UMB9SY7
6KQHNhfvLqcHbAZft+V8L1BXUDq19H8dCIIXqhJNDpm2fj3DOHpa8r+gyXIhP5h1qj7zI9ElxFvt
XirfppNGKJeJHukMO9NOL7u53itSplwiYbbmwO69GeGxTPuYG/Nr3MRM/f2GvNhZjQsoZoQOqC5u
oPVQ3xWrQegH67YuVePaOlkNQTS1DJB8nwiUE9aQ6CGscD/S3QQ5h+qwwTFAXQclA/c0Kf14Pdr2
qoOdTNl2FhhKBHO9UkjZWHJX/z+uG7txOBKOutPau4qaW7xdYUK4DTo77yO0py8ahTwNi7tlhgIq
wSiY+FIu3M4rn9wzQtNXeTYbxay9eHVRLqZhAUSPAHmIyzdpDTHTJ7wqFSGK0YVow/1oqA8EXXT7
ZezVMnVDh+J7oIdIineRwh46kSdZwnl6JEcEcRcA2OLkqhgMwSa6wANHJSFN7EHKxLE2vt1ce/3I
ngD1YI58rpEnyLU9ul5DmyUXgXL52kg5u5Z7en5WODqltcvmIRxx1rwK0/e0pAxqtPXzrgpcYslP
p8pjifUHzWJRttQi4LdEHyjz2EGS+Vio3bF5m/tAadI50zDoZe9BClavHpWc1taRzwd9E2VObMPI
EGpW7LuRsBnbaVI523SOflIEeocW869fgNli1IUAj1WlwaSdalFJ7+OLePwM+3D02auv0PImIOGG
cMbZl7w2vc04SRsSieYiAR+YovzHTkGm/YBLRJusfYaiwYij/9tAdaRr8bqiaeMF9q9/l+rjv74W
tTknd5NTWQv6RN23YWvcAoRTMRinDfH5TziPD6lwSynEERYH+0uuZIL/JeRUH1OcRjbDIbMZDflX
1AWDWIT10Z1/sNACXteY5k2apqAY3nW3+puzAbHbMtYBl4lvB0SQplWpQEy4ZrgLjUKlFqfhdnVj
GyU887B+ZGCSsZKDHKaBV0EFlQ375LUEkOLYepe8rZWfoTF4ITuhHbVZJNq3xRlYAY2M7qBW55Nl
irSKlq/dWs9FS8xn7pfIBVkQFKMt65y/Q3a6dtFsDKQt1yeygOpfIa2NTfAyNTrJ6YmqE9WJUQiZ
VgyKqGSF1VU27jgLUZ148AFGnOr+tZTUp3yy7uMuQgSND+Zx7erEwbyn0hz7sMTxEIvqM0CacR3j
wrxJKsznVHQcWGs43s36QZaO9MX4Me//6gbwUX44pD5gN4Ii3KyVnle0cZvakPmczJOXj6yqrH4K
HH7RtGsolXDqzc9HtGv+DC+x4S+AEOtf2uvxeglkE8yGQPsXqeE6kWKZ3dRVBUfKvhZbaMLBcpL+
d1IFrn+FiIAYJHcUZrR5kSRPL4pJoLOS+PNZSazKWpkS1yG1Ejt3g4tJ+3aTstPr4ekOJiH5rwb3
8IWhs0GVq/Q+CUQDwt7ttq9Gt2Tolu1RiW8HZN9b4neeGxlA3YIJTnkBrQ/UjhC7cDRbzIZXZ/Bi
hkd0kUu+ULnamGObRMoH6z7Da64kDwpK7A3Z86OP5W4oiaprfKLImJeHLdkOiPvdYSW9M/ezzDNy
HuLMrRMP4rLteKrhZv3mdq8mbBcqQ4e2QDGmyFW7EYm13dCI2DwhNbSwR0UFRjaKlBAe5jJevsjk
SUQXK7lF3kNA+cMJe+DhPQdDsu/QL8+FsrmBtpE94Vh3xso9n9fuH44nrnIg8qIm9yb/IZnXAQ0U
qysov8Q93T1YfE6i9JC2NmRlWRosw8BS8puvkguEOjnkC5B5oHdAR5HygnBNrE+fB8ihw8cwtV2/
Bf8JBZH16XjU7ELMrYyRGXojYKcCGXjcC0JsfSjr5bE14rg6RJw+gA1SQbzOl+R9Kdqm1IkcfC0i
MoQ8OY0C1rg2lBQUY81/Ghvhe2uodPIsLfW7NQP7FBMOFtSMRYmpWreRLvDqx/twsBpbmkyj89VP
MOSsS0DDHXGTPBI31Z3bEpespetGVV+Whf/zN5D4RmdD55mO1tDgDzKIWkXc54pTOZ1XwLWG3N5H
7jnB/0Q+jBzsGq7O6ORtLGZ+Hjzen7awIWfqC1ptvphz7w8PtNGZBU8NO6g92B8Us1LPIE8cXj8b
LKcCtGoxaJZEmURuD0w87mfWHwKOUTwXkzuXm9clizcXblVWKgVT4t6jhJikB/YWsHOgZI5z4T/8
evK63cV9WBxzmbOP9FzqydqP3dpSH+HweuziGWsZ2rtKU9fTosYQ/UzfJWlebTH1gPm+YbqUYxl8
wLI/kTGuzOoUUIBwgPHHWXS2RWaR3Ge1e2namBYqSX2InyU9m47xpUWET2bStAvCrWr8Sf2rL7OS
3632C99ogYTDIfBCsRIrLQipbKhHpq4Ybq17ixzJbiSg62y/9CxZaK9G1uw4+rTdS/fabequPgQv
pQT20SGo8IOeon+Fts14DTP0ViopwMINODcFEzBfa4cVtZMvCk6uPGBH6wdAYdX3RZncuoI1sSjy
hd9uuQCozmrUqzzRJkivnxkOY5sdXAOFddeTWa9tzoYHfu8u7c0vYK/4s6EyBp1WpqscW1Kl6R0S
izNPvhto2oF3I3yTM7xO2IwLhGUtPU6ch1jPfA6kF7W9TCC2xgAh4lfYp7228XtWygUkdRpBgaiW
RmehB1wGVG7r2CxrdkqM8Z4SIEckfPz3CnacOilvEXD9UYXosgyT9fpMg/GW2LDiHzWvUX1SzMmI
NYf06JDvOzft1HTyf948SCMNMyyEky+bbo0o/u+FapDyciXw3ZhqVmeyyX/s/X3ikOqCzYPpoSa5
FHj1tdnAWrKdm50DGO0Hwlfa3aMU/jD+bdh76Ju0AzSqjvkwg7EuHxYQObpwfjaBBKCfDR6FgF3l
kU25aI7jqktjDNA/UEjQ2pqesQkv2vbexchJ5vfZmBJeQUeCl6te6h81zsg/tkHGbyvSE83HSPuF
BWKJVAPn+Lj/GUKlaFC5U+EImAAOsT7azxuRk/wuR+x6tv7RisQWNGShkhZBeqPUEPzMLVuKtZIA
0KmV9eKd2zHvcRMp5GOT5rm74t2ig+QdH88jkAJ3ZwvbjkHPiKyNDdzpG/Ffxy0+3gciT677rrFP
TDTKU9ywASqG/ACgIZBklGV4JPzQtRhkdl2o8K3XW8MUCTRz/6S4y+wsY8XAgSwozVYUH8fSwuzC
uNzJaMinqKnEg/5uIlpAozf7BL9+yzXAYnMR6sKFjqNJv9YLsxrteHizPNEaq5h+HnoC5yUdgPJY
TR/6moEzIo0EcuJ3Lia85+lxOaRdmv7vx9U45y40ZANOy6pSq0MTeI2VDDLulIInibY14LkdqBu0
xyqdY1y0x645tzv6dmy5hxsWe5cAcgF8QuSsY4IGsRYpJkQ/YaVv0YhowdRj5zQD3SNIMdCqOtYD
tr+OqvAGkIJ7FCtaKL6TUl6pQZCCKWQo4yfv4zWKoN9ws7Vr/gV+UoPJqGSK5y4asgr5ag1q8wry
sMaCbPDbzkIHtZ6eZNlZ4+XmmShAbRZ3V/rX0ht/c2ZgomhxtyM8hcffO2Ghk2pKnahnKwzIKX9I
eLoPqeZT1Gc+qP5NKoGFeu6dwGduBinJLkH6wLBduoF3vbG63JtSFcJ25H3laM5e24lZryg/Pbr8
hdiZSf5uTfxnoWhxIzmHd0C0nox+ox8VvFjGoquD+X/6T9VV6hqhf6Xx+w7U2B6hsrwdmUVQxiJs
xK8oovhDBBipDtHPZfpChvvB6jD2BT+WGdJyscdal8eYO+PcRM50R4W4zrybnXQON66SaTbD9deh
pSAv5Dmp3OxsTNdZwQsKug3ULDI5Jmev3nHRTJ3irdC8bljZqYpYHIXFLtkRoUQpMNpE2FQxfY+5
DP8P2DMCYSdjCSLGOGdMhkK1QGjajC28UNyFstu0fexzzPHf8hrZ8SeSWFvSd138fAkhxD555Uba
sIt2d3jhjlxPBVaTr6E2CaE6LPmcCXkpuAlJwgJP9AaUSmBTeo6fuEVUl6z9e3R+M1Y/4jxdoNVu
BKpqF1G/bKnUHHj3yG83GRf32SUBXc7GxrrY6I9pVanWUxsKJisrcVpDpFS4neE6lbAkqommZ9Tp
lKwWsuR8BoNDoD4dX0jqlvwcNJ1NDW4s+WlyrZpfN7Shf8Qu5Eo59ZbnSReLisLKPhcISrFXPOeK
kCXLdSJ19U+2QxRK2YD37xWrcMowMbUckRhPcycWIBLaDRcy059QJTgLPtJDsRem93BlDQ0HfgI6
lUJ61579ITFkJkITOpHrYFE3Y9aLT90L9AVfx+DEkb+eHonqoh0j9uRWuINI/NSqkzM+tJZT2oAm
BSv0V3rAcVGeUbeyByUMrmbgHE0spFwGCtKrxghgGaZux8y0UQYPA0XLzwx0FpPNfpiQ1NlI8rKV
o8mFOcJXw3Yyb3bSZCvthBuG0Yr88fjz8mTdHNbFbQrp5I18jPUDCKtUyDnAXXk2LQY4J1bU09RZ
ordFIx3MAdKSc461QG/rz+CFYoE7B/6nq/oB6DAOTRSMsxSb9eMVwOj1DqZAojcHph6FZuIF4/LA
uy22frInPXJ/Y78/qy1HbJ5vOWMsD+kYIMdv0CzszG/NmyNagU2vaV9NfJAF3U4vx6iArYahwJxg
0zdjqzHTYY7knFAyYOolAABX5q7Q734tA0Q7g+gsfbOsgptD0Apdn8sDT9HWzMG9IlID4zzxBJG1
wSHoVTak5sfXulMGi+HxaeR7YOZV4ogWlHMSGVz9L+ENNHH0xeV+oIJnsOU7n8igLiQuwHG7w11j
qrDYnQ7PYu6hyNuuhgEUWNZAp2K7clBqZ6+1AjkGnl8KcIU2wYBz9/FgTFqlaMM+HNdhPABCAeTv
vcJRjeVspyMAX2dM2uvh69uRJwTm/HYhwaYh5YUZhHcItsD6A2DP/d+sjm5j5n0xHJKy3VbnjugD
LiIqnrL0JiCWf6LH96Hwchv48m0uiGLzoSiT9R4h/axeErY6jM9bmk+XVJsgLIrYCL6fUFLjeUgi
qeOmjiLgyfQdFeUy3ZhHr/MOkByr0Zonvxc1C+AHFts2MkjaNQ/qKITMWcjWgdD/fIA81ukbcTfs
VlXYdZTGzfyXb8UhIVEzRYDzxutwYVEoT5CmG7G+L/PXVP++R2Io70pWhKInsJ1bnJge9zSQ8QBP
CF9uoQaYZOD5pe7l7d4xJwlT+maeXxLH9sDoWt6Q5DeYN79lsgtBT7tkcrC7Mk0cbKpNVycA+toK
DMgdltcj/tMeacFKoSdNUdJWnQiatSUB6Wq8cKySziPb4o2KQvTwWTD2ESxSoWPDSQ7eXf0sN9xD
/beGXWy3PZsU/pgRO0ERKXzS232SiiAto8IGykM0zr4ORHSrZiyscVaoc9iIJ0gzQp5pPwBBWlEb
pr9s7pS7MIGKeOKEnJjM43EyjEQYhneQflkoXkHIiZvUUnb2yVTPnbBT6hMxoA3E0WSDdeUKK6rb
MXUwVT4qmSUpTiQjdLkoMnnXkzv7HbP6JgYuf6pesiUY5Sm5CVxEprKZUZT0Q3kPIBTbtgq3NAd6
q6H+MYO4OguqoMiNmV3+0wGZRj3YrEn97BObyzy4Wfket8YRgOM2T0snMRkKwTTUgnqXS8/W7KZw
M4dKxOe/iW6h07tLGwD6HjgwayYpuZ3DXWKmPdJU1oSXGa9sFVQbIUHOQPEJTmme+Db50FID2c31
voHagN13IBH0gV657xgLywb4NFdcik1THMe6Dj4Lu3tO7//YXX/zbjAYdghRqyHMVdJ9BE20I22p
4vCQunnmZROAHgflXSTyogezXc7ngDbxov+Mqkn4NeWZ7amN1GnWBLoOgEOh1BoEiGLJ2Dgq9fmh
idSN29WLh7eJKwZC4QX3kQW2z6zrCUi4xVa63wSgdk27tPrUVsc5Y0OLtj6fdeQstbFTJYk2IXOy
0QwuHT1omU8Rb064UJEfBgck6YZqN9hnjpl4+dx+7gxI0lVwt8A8+bvSnhzn6GfMiTPn8kUph6jC
C83qxf2toYXkxnkKquOmy02KAz7VIlQvBJhwdPBXEV7b1BdGZ1k3MjV8va3ceCbvi9btq0PhjfXk
OiF55nI/+d220ZJNTXLbde5xs9JtSmB989x/oFDUAxjwbjLuZ2IMLGjjW6+KxFZ1gwS0bVO65fQc
ip+guPv+c3QQF94jS6Wy/YwlmUdTN13pN3RSW41fTPAOmnEptxSbNAkFniT35gHEF2L0m+b3JxD/
xb1FkGb6s5SST1O4N+u6W5bbU58jYQY5RMj/Uronl9wqJNhFFMpSkw25N+8HfOHhbfFjrYbannkj
Mx9GA1UoDnnNZGB1522eFfCcmYB87P6gaA93UrmCCSc7Tp9652fyjzWyzRCFhFrDOsGddldZx2Gn
AgfwIxxzfr4xSRxGbNPoXEHG6Ogco0C4SkgGBOs+lZaVUYr4LTO24uBB01gHCT+3cfl4sGrM4F9C
StbFF76hrwVi4YVhbNns1Dt4uR9nYHsFNYSbg8LKRBizFZKQWCVytLnD9S0uXEawJzFoXnwm/6s1
nq5WcOJhyLypC4yRLQWG+12/p0hhHBrenDR12DbvxIc47aSd6xauzqAvWzx1bZ7vONGQJuWWK4j+
Hvj+wEFG+uC18xLOnszb8c5zXHFKqkycjF14x10dnUNuy3hJEB7NIdeT6o7Ux0kZ9C6w/IV3PtHs
V8pR3U9M+g93sJfMydcbLXidzD8bxrQKi2gMEufCrH5zM6Ck0BN476J96l+3ZsTAmyP+juIhMiao
cfDAbWK/5/OwwEU2vG9toqb4yKcRbjt4ACAFpeMNByM65mgmOo8441K8Bjq8oPoIfxgEyZ4DoOEp
N3CkHQtTWiGt9pK7SQHWenRWWoXdhdwddaz15pas4IsqTxa9mazRfszR0BeM5iHzACv8ai7J+nOt
x/QyKn0I/omNPsfw00OtOQ+8fbq59SYsfpCbCY71WGreCW0PH2aS7homfGNXgkNXxoXctVzIDdKV
+kfGqikB3FA9d+a/bc/XWZICZtAkBkvMQY8gd6gshynds1ily67hTwtkae0tAy/0mQ2jtcs3AitT
lAkrMC3hngQCi7D/pDRsmg90KbanlGuZL7rhWUzg5vXtosHj2SRBEvqmhLxLTyjCoT5IEpiXAJJP
3eJUbcQQ2z6yGiQ5GRb+h4B9YmDrW1tJ2Ifw7HKR+eX4CjvBVHA6tJwyFiN2pNDQ1HTuJjwJHop/
Kd11U3uc9jx5dpfkG8hCw6zYicfSazQbw4omwvAqHh6fnA8oIM7iF5RNB8I4kJFx2W0vfDH6WNFk
9MUpgL8A5ebj8XP1P0x8qiRqyHZruaigoXTyesfszEsh/n43iI7UxlM0YpkRqUbT2m8R8+dGQdrx
IAnq17WPfh/kTY1lo3Yv6RpKRCE6T5JbzHEdk44TOyvumJsia2TSv1y0fxEWs+nK8x0dh3GE999c
UdXQZqGjsDaepfrwSKmElsuak9MhcjTHoH5C0PJzv++PjlBkZhbFCi70WOrNaWkU7WV3Rvjp1nvB
/MaYKXTK0QB/Y7+Tdw9bsZRyuUM7QPb8R00SFjZ/tBCd6Com/tKXY3MIOSTs1tSSTMsVPAZxFN2m
SBmXD9TC746t22WTcO80TQDiQQlA+zUAowtoWeZcwAnNvVIHg9hkFXuLtVrRLBX2oRHdZp1WjlXu
oL8gY8plaKaTK5CAdMgcdzEGkyTM0+NfvHqp4G4B+fzEBo4c4ii5bbLAcTpEm7FcX7mIuiH/D6iT
fGZri+Dbfdb5qV8Obs88P4q9DxIpeaDWmmqSbtaYU6yIqExqBpoo1VpUo6FykeJkmh5VsPgWBY5V
RCyw/oTysfIwsXa7I+k0lhViqxh+vP3ekEVniQbzCxOj/nsLSC7gBAOddRQw6IYLJYH36yfif8jb
YELM7y4sQghTJ55ckk9J9BiGORT3MB4mnMRv+EhIMfuw9HAjwAXXkeXj1X7uFegwo5SEulK219M6
C4s1MMkdU9o+4srIVClp6LNW9+jCtkGc8acAm8uZeChWf8lGJNWbNad8AAlL0jcCJa7PZZWxwxLd
aZ/SXIbbtchTr2W3EnMuI8QsvGVUizUNLNw8TOzxquPQV3s78Ze0XJhTUy9vSiC/5dIX9bv5aI5q
MqSyh/2TExUqQbRkVzoHOt5w78keJn4u2PXUGqfz0mbSXXWhrEBLcODV8Hqa2Bac9TiGQw2EdSiw
3UHkM9/2W0G93GjYB3JqEyGaKX/MBFsxrRpSGe2RlmqXcTlLDXmUzYGJUK3h6FFHkvUwmd/+nPq7
voqSU5sJflZe9rMUbA6+b7ZHUwN3LVxRoiPXE2j1nu7wbOLF+b8lhd6oJWZh82tIOLXzbG6JXumf
yHi/8xR+Nz2Foz6r/GiVnnDY1InQYWe0ZuPl22jYBur5diAD94rDVnTHT2WWTK3aNE56Uc1F0q98
KCwNtTCRLrImKdXkjHMVL4YUCmvBNVbgWDGWliMsuhsi0N93sorfhQMrYzQgDy6W7Re76wIPOHOO
6Ttdx6gxP2DIlxfRYbBdlD7pzo3ggsnKgb66Ah2Ona0IaUsmqaZmOwnlr/N1HWVR6TXQ+wm04iv1
GZFVVM16oFj/UgMrdQXHDc5je/EyGdIoTeqP6I8srGF7uh3nEMXwoy7mxv21MCBoL53yENHzsr34
ebj0Fj/Rh56I0u+cvKo/pAfGlWhQ597TICfbC8oJOlOyLqmeIGVr2tMyIFiLjLVU/WSLIk0pI4zV
xrn80WpdmYJP48y4ja4AoYDHlF+GB5W/IkEx9Jcjm4TnkWe0eoiJxNx/hk0QO3I3pR4SinKWkxvD
qbFcm+UI+30svHGag02IbHNVPXf9Kiy9tRs9HvgZWti7yvKmYhOi+bjJa3RRKAV5DFqaVd5nPEx0
2mr3rRwO8leYOj3tP1YVK4DdhyXzWMHe/zoqj+q3SYi9TaIkRg14g2spJhqBeEws6wz3Eu97jXX8
CKNnfkO0hk9Up+sNvOgPYTAzevVY+bWOSUrttHupS3kcRdaelYKJPTkuTjkhdPmoyR/fx+zdSu3O
pYA/egN3MSFC3wG0TqpkJZSBLUphiYhffN7HUUmForsSnBNkkbLLJolVYIndSLeEq3B7gqoyk0Dr
N7X0Zm/A3IqbICOseo3bJ6xsQ4uFS06hFlxtEhDrRQ7LAeGDZHHyx8fSwOBOPrb7ZEwxGEZvto+O
dm8e1/B/CnyLJSJrk3Bf/Re3jbNKpNGXP+bhhS0kMvHN1zh26Of9o5rbd0zyeFhevS/S92w4BrG/
qodwj7yuXCkbQ99+v4U4OD4qX36YRGSCMBImCY7/scPTr2Z0zLLiRE/P1qitN0ISkEveXQfAeur4
qU3ooiJ8jePZ15iRShdVwWsGHNlHHtUg0igUpQ3gaUG44cb3W69v1lR+8IAerSJgsnEwEWG9AC/2
EhiueowEJtRHzo3upX1rbzgeEeEP3aH3snCIlnxle4jM5wcHujUR0zr1+02SbRDoLa6AxB4pXQn2
6WHlL6KOW1UhlmCEDQ1pnGUdDkHLURLa2N0VUK7Y7TWQm4uaBdE7Wloa6rjKZcGNDsfHcpjJcoQt
Av5Kx4ClGzgoqs4XQBN11FDCEs0W8z/yopxIHG1+YRLhBrfEW5UugU/tSfsKjXNh0Hu3gIwN3vV5
dR4fAx3Vd0F9t7m6D+Rr7gqv4xHx5EpX4gLTCHxv4811bzrLD9MlqTZAaGkJ+FjPn8NYY2CViVno
DixvGD+ARnLagLRGCaCsZlL+ZhpBRW4VvA1NvbeJYBT18iSOlVtPOuZvdueDLorD+V6ToJGT2hiu
6GvsJmwSAjSBn2LjKFdZfQde/DdHizwCml1dBoOJhI3nJDtIFfP0hbRW6b3c2ttm3vtOZQE7g+P9
geLJmfIpwcvVGSuO6aFfy5ppi5RbPcTua4J7kHbH37MGfjEN5+QzNo02C5aiXT6umWaorrkFp5Fm
+uISkmvzhZlcjOu2xpsqKK+NpX8Ye1i5o1a8K2OYqPSI1YmgnitXKHmM6brsQANFJ2gSkV4MvyCZ
2AKoKv4TtuE6e0pc3AzUxquxT4JoKgeegZEfQt6o2GRZx0AcyrMPOXDQRYK6bKocN2PhxSmO86EU
zeW4DKk/5nN0pL37Sp1hW2pVvtDiSIbBkf5cScb7GzroiDBJlAyHw9HirsHrW4D2MYeMZFBSARXE
3F/ly/y+x2p1RhOaq+HCWQVvV9dnpxOjQln3p0HoewNHCysxGWnsYKN7561Pm2hG0AWmS88lzkE8
iI7nHG3MkmJCPwKw0Bp7MXlSL/cT0fBkt+/Gb6r8HF+pmbA1nkQEdXtPaIp3Cz5LmeHDlXn3Gn/B
dPtZAX57TERZCtr72rkvT6n5nWsuG/5oKA/WNoXTd2ZreQPlhRs9lSJy6iQPsaRhO07OoCh78S6M
xRMAYdwka5U8jekDKcVzRXh4SbNGyyffxfTxUDJL5cKPFPY3IIbODfHIphB/04wOINHRY+bwON3T
4Sx+MvG7+GKAGQOFPG0nqen8vXju/kboV8ZvIfE9hMW6q7eAC0Bx/w+EQDIjDXCHwSyoxN0WIxtk
t/0pAtKY3055ykYWJcGS4vITg7Eb2hc+AMctIOL8izAcVSm+km7+pbHl8/nOmje/iueWaG7hhxYh
fbiebpls9jw9WKT3zGIXX5Z32OW8evOz6IDia6fieu1QglERK0B284W4INHsQtt0faeTCJK/LiEQ
KAV6RRvVANzF3/g5Fgz7jnj3haNrXxlqFCUDBexS0+fJJDUVVh0SJQi8J+Hsp+GdmeZLhAmzShKD
HpP6ORJh/fp3B+gruxqW0NGE4v1aa19de+ZCtMrJj1BBdwDEt96MYDqvORzYDHJiZjE9lGvdGhEL
xtYlz70JLRIVZeDVIAbsRdTsD6GbP32UHGuALC7l8D8/8/m914IPSxyClw1H8zavtzJjvxYN7cYE
a1sdy2sEaIA+Mr8+EbHaRxRPBngXq026z2AEMgQsRyCRloKnPStuMbLIwf6cIzoZklWr46q64BpT
jopj6p6jTEdH6ydB4jXJNoJ1WvvNFQubHphFzsqfLB9JlYTrWx2c3TzaAio5vAOP0zg1PpKY4o9i
2GQkNsF+xcCssq1hJ9Uyt0a4CHlFareT9SmeMB+9FmPD53feO7cGfkUeWRKvx5Hw5UUglYUwEwe7
p1ZlXg8klC9cJF4iSUD62KULR82J2s2EEurAkEwl0z2bWCWRswuPCeqoZiJQbDwZHrasyhqNEJsH
aJqujkBc0RbQZDDIkVqx9deCccLH1+NaSvuraYcxWCBYewblwAwzaagaMdO8Qnhinzqb/Vt2oGzy
GPB0FU99YnR8S1bwFkMh3sgVCRxhN46Z70g9h10pW7cmy8v8oIuDI3wpa8MUz2diodTOZRww6IJf
oTvRZMZwsVVQMaAR5d9lKEegkDchilJWQ/ZWjwEzbkw06u5keeBDhFco5YDT19tIHZ7+olCndYEx
JqONCthmnFwYD2ql8YJD1bNTgSWlcbZL1TYHvul4QV/fEQ7FeeCpLZor+K83q1h8c1P/TODIk/Zl
3vKWbeVklLmOwvJbHBYpNKpjpsp0mR2fxB6uSge6qbd0JY5HvemRUW25VHlJnU+t8Fc+/DB/WiCS
Z7JFuBOwzvbPR6Vxw7HpcyBMnF6jpSS0j6eze0PyxuJ6SWhSpcRSJnFThphufsJxR+TCfw+Qn8wy
IlbeggtRuQJ6DujWPAlPgS0ZMmUksGysIZ+JPc3S7Hog6+0siMI9/2In18jjKiZIT3eCGrs8iLNu
LAw5FF6MZ8RI18w4fgMsnDF+Fzp2zLQZJ8md19bemKGZCH5SxmGQdB5699dqgk2psx6+RruDZNoq
WxVle9b0/16ATjvHnoxyAqyc9gjyGC51ZmrrjUjMaFENoaH51jOu+jEnoMvPEr0Rkq/z6sLrkAmp
ulTA3c3QAppEPS5nkazxckx71Yv1JN5/VhGfsw6YPBEGgaXndNeFR8peeOvACvzssBpAu+id4lRS
1MCq8oaMQbvWxhW8byxXa9F93Qb/Xz2X+JKAMhUjQDGGP12e8711/K4C+gCHchPirF4GIOuBAmUj
1/UrUUmd9n1RZ7FwyNvconzIM7nvUgINfxiz3ya4cNy8VZFFYWucSbqz4689UAtIejBkldTNWKZQ
JsfTsZ7NQqNkHQ7t76Hfiq1PUBXItvlNz6SwTZQq/dXxo2W4smuACC9A98uaTUtlhj1fJJYrmnjG
E/vQXim3zE/jB1ymAS8FO9SLad1+3Gi3oCLJ001IaW4Y0l/0z2PO4XhP3P1yDsC5UWMBNnKeDMh+
pYE2p9bnGusFB/1n7YCmf4NZ6hmTjQSbb3AGg3j3Rj+zZPFI4avlBhq4H1q9GNNuQm9zFvyU9jQf
Ip01LNUoMhWKk6eeP7p4iS138wHjsoD3VpFCzZqUHrMZSd2H3pyOyi/PLDFcYWLXYFIUjJLTy8Mk
BOxCBT6LsTsGopvJ3+sGQNbWK0Uz/EDcdipCN6FOW6GiXsNuo9l4+2jtP2m+qcvQIAjw1QmTvpoH
zJ0/zWq/sXocimSTDdIs6z08XGRzPMUbRrZ71okTy/THO9rbCftcF8VxVmgWwRWEyVRqtiiOKUBU
OUAPJawljfdkfUsrMFX0tfkIwMPrqZPxL03VWxX7U/hecxzARB17YxwI84CkKQTfdLsv63C3zimE
iJxAEd122L7JaJH8PcCFTA8ADGZWIjFUntYdD2B7cMFVE/+H+O+Fa0XMvEzsxS6iHmZ1juWf7sOM
euq4VafOzsqc8k1B5wCeDC5kTFvJHhMSBStoCgZPn9qOFOcnfEuwWXP0NqGzImx+2sZLAsgSA34O
DvsyTM9AI91urYe3/up0eXpdm3gHbRCNFbIO7FK/DUn7ssbzT/SARQpgKEHrPGiUfMywpZoLlT8+
q6yoDVEJfAYU2RN0A6TJaW79QSLjxzgaK38gSFmRExs6upo2crJHgk+tA5tk4hVuZnEI+QrebzFa
4jKNOf4yylWFn0vU8Flb6tJ915UF87Ay5G6os6yDHW6pqIk79M84SZOV8KLUQ96LmVO693MJ1PIR
rh8ZTX9lfiUGrXNK7cPcbnzonDgoLTv+UargjIzuBRTrBTgjs5XFqrDTsBfZsiPQM8hzo5uloNMN
mfkaDeQY57G92Oz+LpHZEXD+GTrC5ep1C6tbDQwVhndJvrV9XHtvmN+4Khog3igwHWeuF27IVr4i
79l5yY0+sw2BQ79xvrjNpYYQxIQXZruFbPIvx0B6lRxmmHkZfcQHffWVxbG1cl7NLPOxQWGyGUs0
sTwWOvMjhhgtt4swRHsaKRR+0V0hxLjjvqQxN+9bbZA/z792vadFcht7Me7STYgvkFKQWTxdZpJU
nDny3q9hX9HtseS6nRYwgrLWuQnZlox5d9q5LH/Yg68iuOhqQKpdQvKHl8uuJbcmUJrH/E3htl0C
ddXyrJJCoDBeLRiwl2ICZ764tSbVcfwNqVjdwjYtK4yplaqViLKx46p+vFvfs273nVHNjhtvzz1c
Ge7n40t7onOAoMM8RFjmRcGMNG41go675BJexUf6wXyCOyyMfUFwT9DwoMK6G/vvBL7bNURNzaS8
pxib8Nemr71/M6QJ6dYcVMATMusWLib18yWGv0OKGnAbDc5HMzO/N3cE8PBf451/x3Stnbnn7/V2
mqUVbxuiOxz2HomqlXnQvdQ0cc2zMha6IXm5HFIIFWyANk5uP29QbIt6COdpMwSgOKp9fvKfD4I0
7kMogyhzBJSl1aIS0/SyGlht9hwgLQrPpw6lEC+bOf67D/XuKgccNoTr/YDDemwPcFspvjpuXHSU
OkDnPt/QAipKvClnLA3paLkNEwWsKy7IIQuKgWXT5WbdVOhmriGdL/Nq6ijYjuZxPIOnBHxRg1yK
MukKJ/zHE1x2KjXoV1ADmQUsOYX26DWVYPHzmz72x0FkMQoQ88BCHWOoyridVXjGTrlGZznbXMDc
2DpNhORaCCzbCMTxaQT8HbiMv6zvEQjDLwHHw7jRIDP+Tz4Sa7bpUKo1E2LfYMv0jjT+btxwBFkI
sM9UJo6NYmXM4CZrgKXDqnemtsxCx/W92RjRq6TXNSvrl+GjsgGndlD9//tt9nMoYdVK+w0PWJAV
pVVoxHM64RUy/IcVliq7//+IMVXXP6ka5ogwiGT00Ql/3YH3lMjj/0/eUyED9Yp0HjdeFRafvxT6
EKWe2Qnua8TXEkul+uHkVlubFJUvkCJy1+kxlX6bejM6M/DIgDtVepnnUMk9xlzDTFL5/9EpIZlN
M8MebinFqLAAj64kztw9RBwtfcB6TPSxeXhjzlRjx50CiLbmmFx2/MDYuRnpE8PvWOn2RXOGSIcC
W5K1+v0ikIxA9RN5+JRcm7ECsnNH1XJY3HuQ1kyXyqa8nD9MB/iGKO63ZSU+W0fMyks4fPcX8Nxu
AphpmmZrSWBD/Vd8q49Er98WFA/JarEGGaix4YAZPi9OcalVRxyvuijpbx2Oz9fCXZoiOf5nmdNa
v3f70vFOsPU5VIJIHQOfOwLYt4TrOIjdbK0npBt9Uu5OzfEPVbpYWgEYbuY1ZcaBu6WmKOkiFAUW
u6rT+8xioUnn1gViZlb60WuGpWtgKEBmQs/wVaMogjvWwRTgscSmQR7pRgtkicyIhWzCkefq22AY
EwjmF1BXVVqmk5ECAqssGnr+5p5IRNTNsCOjB1rxQLXYcOQ2OGVJo09m/8LDRrs4CxP0AVqxSN8b
PoViaH2GFszRk9goX+e1Rm6XpzqNyg1qUcNnWPDp62NX/PAk3wpcu/4vFqFtgVde0KT43B96TDNE
9maPkXjLpgAQZn854WWO64CquzbZ+jqNoptlQi363w+r6kUrC9usKUA9fEtEf/U0POjnJsr2VOzX
Tdn5JHqiaJewMyz2CW+0bOJpB6WPxdyLI4hH/7lycRX+6/K6wC+GZz03UXthmPcaBHF2TKeAvuFY
uZo87HtxLBSb5Iq/OLIKqvfyB7fmA6t2RN9Ia5dCET7W3E1wVlO2hqNNNQMUlmgkmTi07LhZ/vcv
OnGzamyNrymVkihLtTy1pzW1d9c7AMks8zPLUVKNg0ljhgrZmyuXUYUbHEvqZquTCfOibEz1iXNE
ArZy2HO/p7laEiprT7TcpfFVxXRqnwclYxoUBwekDH7bFIzdYgJW9Y6T1Q788H6M7eGGGrS2Oy9c
K3SwI94t7/c26cUEFdK99jk/FH00O9/BQ1R+U1kB0BtYsT+/rlRm4PLu69UI/Ovy+AmMwkk5ICn5
ZHdat0UL1bzkjB4itUGLTkCmfYpNBdwu4QSPLoJN3SDUrE3qPWVmycHGxUbTrqwV1UXzpc3Phtxm
IJDt5hnSmpnURGo9/ixkBS4JxuSNYVH4KItOiJSzSzEDWiCDJIvxBboYNL9dHlLBY1WnGKbt61dS
61k6vgPkE6x7C5o7JpqPXfRWcVLG5U4vRX6cjoch5K4XfniM1C5Q14rjzryGZygfoYXfTjwLL1w3
1OPpe6+wQtj3BPAbBxlSWIdEUKh9G8JRsBn8xlVrJ0qMcR9QkYtQY4Q4MUTVHSa4HlzZj7cr4+lA
ih7TYq3ZzEJzOnRppI9WNdmT9qtiOVaECoUExZL342F6MdVl8m/Gxf3GbTl8PeuYk/VCCeD80/XA
SCVu3H/f1MPcke5YznY47ZmrYXDcX4SnubpL7en1UmLbqU48BzTjqcl9vpYl9/ythAWWR1ogw+Yw
bxncwmUi/KGufxsxDSswkpJE9Zhfa2XEgYv7+Mo3cWT/lcHA0y2J/x6hRK1pFRyrB3s2MEfKc5ps
4/ET4UgkCnmqiEccjSA2N68FavKZyjUOcEuYc6Nez4EK+JG8Veq10r4rS83NzUplC7FmyqqUeq/u
g5OEgSWMlvByevbgt4I5YxWWa2M2SaZtE6X4nLLxbJ8um5LoQS//sOk175pcr2R5vjUb+D+FB7gg
Luut5pQQWzWOa/DvzV2MPPZhUiVUErAS3Cf+3y+nSJeSgSI8ojpyvI1K0WQLh/ojSNqTj7XlQb7O
XDiAI/AgG0kgloJrJPXVSFsm2Ue5YAWyfgLWJJp9RiW73r/wsZGR6dESc3RtrSMWKitTAFkGg3jQ
C08kTA3dPQmZ3D4we5s1iQsaXA+aJwoBwoLJTVsBHl63xJQ2BUGMIqXNnZeJ9ek8qz4QygoiSYDr
PcQHe8jfWA5EttpZFVdp7++xIIQmqlKwGCyDQlhgku43S8oMSSb0QMm6XGU9vFb2WIB0TZKoHYgv
QZx+qdt6kGb4Fqhp97qz+8Za28os7xpNwQN/h232ZLfuHMPlCABz72muJ4R0OoFkHW8u2FynIXHG
sokBXDB4PvQvrik65vvs10U4YYnPhKgGTM5Ui/tRhR+AW/gGgAPrB/rdcJ9Nuzrm6dwVb8uJhGjI
wj9YTM2QPRtUj11eB5fDAG8+3pqirXkRvykKFhdWhPTfuDtM93QgEH51d3UrzTpRvBmeE+ika1lV
c9i1orxKpieYpFiJqqhGH81AU+dCnEX34RVVFg2oIJjIC8d+X7sSj+aimKcN1LLGew3ToCoAZJUE
NcUORFfLv6TSnw2u1hmWq9FZGq2kFqMnVlfYvvBGbSMlzH7eAGHDnDM8hv/Bza9zZWl603QPpWs2
w3m76k+PlSszVo2DvkEFc7oSZp0rCISSQC0wQ7jFbayBseGka7QSIYrXSzDHZnqp+T8gOoe9XWFl
SKkMWU4tZgdGoe1sg/8ESGUidV/hX9ZiwAZOKWYCHgLC6xIM7/UkNWwrdXpfkDsBrmwaB0mFOoTq
FegSyXcJilHrgAMEL+CkhHwwvtxH0xlM5uIgHzwC1GWKRew7h566WaP1GIlGSMS4AcOMVEgo6Skt
pDxx/NWtJ775peCfihVrNjHFncEdAue+wOqf31CCkrQ0NBQn7J990AFECGuvASIK6eABF7O2b1eR
BtK8ObHeccs16shUS97THc1pMr7yetcBGi5SZAKSTJcGU6jBrwthM3EDrdkic6fuUuLp96Sp4NCu
IQgE/KrRXpp8G0iN8T0D2diHQg1IeF9r7HwY2AndjtChk1aRbbI1rL/NSCwea9m/q9eoej63Gjk2
XCs9Xue0NhxSH/rRaAcOPS84nIhhl52NjRae5gwI+ts2omJLDfbihFA/ndmZRuTroUUGCrmMbc+c
B9CSiEa18dzfNq/YZZyscJWviSPx54+447xS5L3ZhfeodfP2j8HGTIfKbwUZKUQMa98h3fyz4O9R
wIfHGDxcvQ937weWZ0Py6PCNRhqa0mEqDlGbY+apfqZF1iFHzrGV/F8XrErTf4ZQSK9w9/sJXDmG
QggCWIeBUpQXmhYlZKPep1LCwgdyJaB5Y/zm8ahMTYbi7K6A7JxAeeK5t+baJSHnxJdmBQlr/vLx
5nJ/gR/PAZy6F617J8AbRI9o1LMZ/QjcKwgG3v8UL0i/RBt1efPT66x9/4we7NCjBf+OnfbRD1QD
AELO+i5KqKM0b2S0iTqAPb7ywBf82Nn7nXVpkNE36/yj8ILdWU9lPk1EJCKf1BJvwxeTZ/C/ZA34
XrE9LYCydQTApObh7+VFjlqmDUezv9CTDEHWUqAAYUCGSy1pvLTZblw6C0/IuJ3hTdOb0mQQvZdA
eDOeZpGrbeJOAfEgucz7PQCtT5dmEj4ThKPJ6GXvaNDQXXY0IlgkzDAkD6Jj1Oa5jv0kkKlaBwMV
0sJLuD8Yax5UYMJfSNvM/ZCPgb79s2KJisemD+Aq6FcdP0oqFRKWaDThc+zeIHVs1At4xeOR1Fwf
yuChxel9UXwqVTGYgHKEKrkmBBESQbp0lFJzh9NnwuTzlFseBwlHw/e1EuKQ7vudtQfdPDtaZsIN
Mj3wExmp9y6URKfCmRsrfwRFELT8qX4v5HxJujheXK2BjiM5B5RMN+g4x3wvQoTuwyJp17M3mBTR
02nnSDrS8WARCdFW0UhfghQ8elj5SJjK5H3/tvnezSR3RDpJE5g4BcoYHdYtceh8Hv78iciiUnT2
darAvRHcfouxcCO7RyXmfan8ayREK1YjFaXFv56WXd8w8WW9KfiN83Rd+nhhi2RG0qsk4rmv5jtc
/JSLr0xOYKbExvLGu8Fw3BaJ/fEqyyW+BAZXNCzag2vBQwf21O8CM98HXVgZ1SwAlmu1F1Dl6Au0
zui49fAMHIc9nmwdwPC11lE5Cnnjd99981siw0nIa7o7UvdwSlSh+30nNpUUdPdkAw00u+9gQHnQ
HwC+FigEQVd2xdsVKlfWOQUYJ2ePEE6iVRKtMXiBCriFvdFfqCjgWT7Mv5d0jJa7eNcBPvxUJ2gV
YkQ3pzkssLuGOA7gIULhVb4Zn6i2ZGUtWQCOa0Ca2plWRSN57WKdqYUz2s1l2jFXGvhJ4U6icL2c
eNrWJhesiYuC6EnkRoiGr0BGmPKvsuXjmbftuEam8P1rTK1C7ZbHr9p6v1uU4AXGZ6zyDyp9l+LT
hbcS8KSnk/fX9LEru/HCT5nC4UCl/Goh/0JOygAlG+G4gsqALWWlZLFcCOaHr3SXI0E4GNrpHV4R
zcNhRivgAI+OAI9xNeggPagJKpc+Rzkru1CtkZ9+bQhkWcghH3vMiwrIxR+WD0i2rMGtIQO0Wn4+
Fh9FIb8S1WB1pgmU1ComdjsXLwjYCwOZAWxxbGTM7sifIgPxCWWCuXDPsl0TRm0iP5llOS6lRasE
jF9hxDXkTpYTEcjlfqR/+yjWlf460tjs38D1A2LRJ4YyfX/hJ/dOjaDSN+ZWqGMahMIYJ06Hr2mG
eRUfKuKXMcosgCF0eLX+kdUj6V9U1O392gi3sXd7YJLHVQ/b5xp4HAAXbudoiG9x2ocBCPqIRq15
lhIqEwEPNba0PeOwJFu2caMZDRjOm7e+1FyU1JTk4zE+qUJCZpyfBFSx878nc8ZjP4Mir4CoDLYp
7jdRrmYpi4uqhapyRL5gaQvFMy/g4cH9isI19Sd/19gFB29AT0QCDkG3YXADoco7LcrUWybUHqUE
lYKhhHSrcSGdbS65xxx6a2q/O5WTV5dqDXPJ0s6tytTpKvZ4gV61uVrPZUKuI3w8AVFeAXonD/Bw
mOLVYMYBMlN2lL/Ab0zbWKtZUUVgu0UamRjitbG/8ImdvyNmW/0T4jR6B6ttd9KJZrR8iHrHSvZP
7FpbKMiUgzkhq16lvmmVuBezEhWwXAZeDmxBrOHucQXvBxXFNkVFDkrjY7GXRWohPmMBJuePi002
bxk1EiUOji5BqZAzsuNqRGSm0cQYiCqMHxdbcgfWXyzh1v/0dFsRyODfEx8vRH0TZLsvD2bhQWrN
hNwChGT+CG7Y5aG6v4JhEieS0AiliKt5XQviZhVJ/0riorc34S6ce7wpjSIFl1hbrknokyu81vh8
9i7L6QxEFGEbXBq0yNPILFmBHB4Cfz5+4r5OlzHX39G8ZniyZwQXSveSzniFuCjF7gEw9IQM6qSP
ctZXCpPvYG5znNGs0iocpJCVqmkWNoMoi9jGNBnXHjj9e5l3gPVLmerIu3MZEi4u2kq8CWu39m7R
gV7FXISVTLlT+cSrLtNcTRlplh3Ti6WnYvTXp0rTTQY4kJhHIIevV+KFzFMnvy4Af5GHAPvbiAld
sXq4GePwz10UhHsatpZVzRZH8gIjH00TBhhMY4PG2aVU/pSerGIh6oXr7qXdO2qGdeHVjSVyTTuJ
R9rr0zEaRWfSNOjAgEn+SAV8as04O4nPdhmzrdO6U0rfBDFJ4dkUPaCCmKK5BC0iG1/GvV3sRy0F
edRy8UzCVm+8KS/m03GOw3kCvCNYecKMBLpkQTjTXH9GMYpdoxG72SY08YLrd+vmw8c2PXJtkBKl
+aW2t5DglI3/VUh0bd2guxYiP5HIt7DmIEMcUC761O9cWcLm5ntQiQiOJlIhPWYr9q59Ye0WD+77
HdC7/Oy5C2kNX7TytWo6WcVSM4mGM3VhwF61DI5VtUO9mgkf7Ezicd2Z0SpDYcZbU9DXaGqdVLbK
+fh8DwG44m9hUZXUAb9ZJqSTu9oYPcIH+hwZmJsms2Cozv645go2kQaqW1D51WB9fjVuO9xpuMnh
qvi32IBsnGnRkqUxUEZGankNwlUL0ZJykYRHDr745UbN5gWYMIbtTJWUFLCsPD2+4i4+zSOBV+Xu
/i72WhCr1KD0MSHfIfFtNhbAGB6rBX/ygLpcMY3SuXMQpr3qAhD2w1p7BvoBICYBBrHrhhj7qJV8
Jn5hWQn4FPPJmqQd7HNidrx1pYAEl6P4hqkB+jgOsBaaHnXpIUYnS8CyGAmapLLgUUu/syKag7D0
fxYZOF83bBXbRzzbtEikcJMPs0NQioaIEBZqbMlVaygBgxCPWmxdiNZK7sABZu5cuEruBfCmLZGv
nypNT6YLHdNuH/Hxp4+KZ4eG6bNUh5v6jzHVuX6E+osJHNxoLSPhOw2zNn412CdyliqzMG2ekljo
M24MmbfHveM2Z5TmfyNg3dJnbSjFIfB5nei894BrNWP5ekFdP9ypZOS4BZff+c6mMH33RNjpkRvr
Jb0nnUf2mgKC44RxnPNTxpP3e1qI9jwr3ToJwIQNVauvVlR9/IR1k549CMfSM8QUVE53we2X9odr
KqDxd+DOrucrGtDs1BauD+ArowIdqPsg5iQ6d1Jg6zeC+Q5xrGQVc6N4OHGfQOdk5scQSp/ksT/c
+7UeeDkqqD9owr4J6AX5laDyeDheyjKiu/VYrossBP5I3wePUejk1OShpqAuvPMQOO+mCLktbes5
E5qr7KhxmBgCyC7p1YYKiv9qFeyp0ZQ1KGsDBLr50+bd3ec70Dqu8aDlC7/ikzX6QqLm19im1FsD
rSzRlgAOmf1AiBff0JCU8K74jF1CQ5OmD4ZrJRLVw9q5fXQtHqvEGu7LjPpLITtg7ZPwWg+uVksR
f4so6p83UgbKmH4Gp+vzXFdEqsUvCnCKSvlrGzJiSqc74avkZ/uI+VVEI+Y9ElKMRgajbzWSqTO8
wth9afrZn2kt3QQqs9bkfqmSnSMMfmVcTZh+2lQMS+6l63XEJIJM4U+iSQ9i5EcWIAJYMddqH+9O
tKGbT8hH0yzs6qhfl+m68sNrF/1s7e7GbFYtMZ6M3wkvbtJzmtyK5Pyvmb4eIr/rA3EaGmjvrA1E
diFu+Ud7iPzZ3gRzgUOD2OBBPSLd3m1kjNRKqlnXjHSBRSzCEid5IHiRniuaRCqtpJkoaffMdzrG
9WFH3W6BF+HpWvgO4Cha1dm8wNVSg95MIjnDAg+vRFjYH/EVIWbxShlpXVzJNWUdmPvy7kSfHMhc
b8uCM17vrxal+N2FEbEbDhR1SwjntRrJvWftjtfIhWGwmNvsfYJhNNK3cPebxbwEU9qTGqT1voF7
am/Qpnrckx7BIBqNFnQgWNxCoNJVA+/OxuHlEJNfivvWDzE+iWaIujViT9Kzb7Qey1O9sx8CMpD9
hDC/rfOsaJDSYvHfm1toJyp8Dne7mVmSDBqSEq/awr+fYU7qmnKojkVN/DFYZ3+IlxreQnBX02ku
DFzAKC4nuHfXSqZoYjnGBwe1Vm9fggWn3CODG5wUOq+K28GEbPyfYx0sEDfnVISrrcl5X2xq/vdV
x07eoaJLMwg3HGk+dtiyPtI0QH+jgz+JPiy2cul5q/cm8mY36VJaX3Jj3agnIbHoHWU48+QP1NYg
DDpgHWSPjTBb27KmanVeh4kjHPiQMCO+Sr4ZFqHA/8ErVMmA35kI6uR/1Bqhyz+VwEKVrv8lI5oo
EjZaorbXwbx6xPfNTOmOddrLhWpYlGZJcPhNoYBSj8s2+OhI9IH1531/hiOLa/39SF4Ovy1brcE9
eXnG2Q+dqnbRbQtMQZKaisBYrJRgF4U1w2AMmh+giZj4QcG3Ab8fPmPn8j11aIThaZgsNEvseFXS
u3qHR2TUJbGvJ4isV+xAsNWXb5W1ujzxdQVNlMJ+dARgYgN5Y4LQeIEBXqMDJavWlTrEz939EzTc
BA/VaC/2bfzIg+RCW5CQ2pwQBNi3VtqdULWQQcFvirGkneFXKp2He1YZoZndiDBYdurpGxgb1klU
h+dxItrH1kInVEwE8X+gOz9mVx8qKhd2zPlvPfVK3bDo2P8Lr3E8348dO/hdvPNtBPjf5OV1KdxX
1kbVzqnL5QPfbyOO1BpVGo0xvz65lngI4jg2uAHIZvEv55edbrK24oe1lYgNKiifC1zgJrSbsCuo
fwAp1fZvUuO2f2rxLXz634vvSGqF/D63W0vRJUIsPgiqLhBTNinHfkk08l4veBNQf9mNjgcfPqRA
2d0kfEv5XnP9y8B1aU19C6NPWIk5D/IMGz2PDOWfZ+i7NurwN2FVcBtC4jdXg+Z9Y12VLWiatu6M
iXfYD7H35muMb3D/6JkeazlgL6AP2Xq7vSRIqUxYb4uWbyxcfuChCPB9BhcWXIwCsghRc4YiYnq7
SIPg6eYNbadVH4NkEM7PLDZsB8/SW8aZwJP7on+cjKRu/qSl1EdiBHQve3BiQJHIh/d8gADucso6
sRuo585gjPwHKZidlJwVba3mwIQsKLo6EZo+B+WWq+crvCrmMUWLIzlhEHhA3T9HS2lExWWWiQJb
vISSjY04qsGKrEke+GUIOb6ier0PQoGHCoh3GxTyWlQT/XNZ9hVRhGPIXx75MFGwBAO9ddP+AKSN
3mFteHGZEe5es/106mknKXC0wJuyvgGFcONDkQGiqVwoQrAU46rtxxw7/mTAiO6KUg2BISXbzy+8
hFs0mE9MVQIVB8sedv7B2IOf09h5zYUz+JlVN3dmgVkWfoBQJ2A3Y788yON4hcNp10RwepvLvpF6
a7OppV5H0Zs7OpnLJTJRHkvlBObHcZJp+ZoHWnpKfP4/RqNaC2cqcFkCjd6w0ObgoaO2MpTIei7l
56dwpovLUDO5LuQMxiUD02KCnBUUtWOwU2wNSMLyDUOAwTYYY6fSzFg8ZZHXzigGkiajjrr8qd9u
GFX6JFf0lCcTVhIYRX6fcSHdHEa7DmrXyTqx8KBn9rBBRjtWw8BVaT/mTGKHkUKvObXdkuYMPlvC
GDmiVtyEuoaZpgmHfsqqNC81fBfjDUhJmf/UwnwJjoCh05w7GsU2iYEBwwDirtpPb2qvNBgaTw25
vamICDxTB7qmz1P6OXnOnNtGQ1liAl3iuUG45ugr96pBh5vcrKeK6Ixc23DCM6NigbAO8irbgYa3
bsSZhvsUsLBE5A3iZNraj2XwesKblW5CfuVF0uSjAzGZYlSFvz/EVK+7FoPtIGSzIGIpIDfZWaeg
1glGCcQ51IOIPwXacgDHeUvH67di7C2M6/pWbXZEvj62SEl1HvJ4yBYjcxF/SmSZPl7W8Tj7ifBl
MBt4LOm9JHmVp11/NV0x5jQGfuPwsalBLXxPmPV/5Bm7SOMoRgTNg1inCzXoyC4FK6RlG7UplSOA
+2Ko3Nmy7LXBpSDgnqp+ZbdlkacB9ehXCdsd4Ux4UDIeYAClyp3u7YPAQP6R+zKgUmoJMEb1pkPt
8/njs9sSLFnKSlVFK7a0t0OdCMkPhiTGzBhNhzbXHfZMzNwMD+khsEHVES8+ZUpeHmzfUNNDnybC
stZDRoeYdfyFfEizFcJ155RuhpxcfWUw6r+SbIWn+XFu2KjWYdmwqv2NsPL5PizWXDJqdMsfO5O7
mFTnHuFxbvOQ86JFx3iAxv5LfawQ4XfGSYIRhM4KIpLhwAI6wGtfvCnERhLSvk7duPZ33gDZMwwG
2xmJJ9PM76TZsUjrXSqBDFGavTP6lK1wuNpTvJJCIuGyOiZpEuyQX2jTJQ2Rgz+HQslvyxP2G8f3
pd2OYBj5lYTEMsE+XpSxX+TWnmr4n3kWcBrbD/0ombeVZeM9NN1mWGzrJzLdeDVmOSy/Vr/Ini7E
L/IR8afdK44R4xQdliajXSxQolI9HMVb/mM0qwy0iVdcCVg33M6FsqmsKD44ZtWWKbWYsSXzemiK
DxiHkVsz8xmcKJ7pCsX9jJtir+iY9R1aXL0ej2HdWGdWsYxCsjNjle8YY2cRngK0t8lpsgyb+Qyw
ppt3LjZhDteO+NrieO/zun1eagZB2RlSxJLXn5BTYVJIf4elGRstg04cufLvm/3HA029J9s7Nxzi
+iYKDRu+/7d/seXPH4JKyFrtXFvl2Afk0MApqHwZniVrDU8fKbwDtk0Ff9a2OYgni0OJMUAggjV9
p9V5tTJ2pRc59pIg4Dk4K9tPtX0XiYa7cUkQrtm6xYy8v/B67cg4UpUa77tYgeSkf6jewz4ETEx1
vGY7qjDMeHJEyNb9NNeeu5FNB0G+Ol9PvrxhGbmf8DnisMHiInmiGHHRkxRVLNxqkeBjLNsXNCoi
DoJe8Mx6oT8KSbGxaEiTvS8uHiXhWe1ySu1ZrZMhA+IT6fJUq8BviTzehnP4DNduxURRyg/zniAX
FrYiFU8LSkxF11loy19oOX+SYt7qmib/1j2rTQS7dMd0ltCa9U0er6bp2ULGP//r7ZGzzZfDRAtE
PBB4ufSXBdTjVvOUNToMhiIrQj3pTndycLS4qUGGO1A/98AfdZw9kml9anlzwuZLSYmfDVxndJPR
73+z8XXyTNT6nqAp4oH1OnwAUEr/bCk00UWshp63ofuocs9iu8oJjwD4hB5fcsbplb15YQh962kP
sHnSAG0MltHWtkP1/b/aShKM/7pVSo5MiS1meo9KBv9Wr3/+53RAE48NSXiphKttP+JqQEVO6Z73
nVjhV7tqisP+ODtlr2pLwmu+llPXEgcEQk6NtTsSuA0dAECYJvHLQ2qUNhooMCgtqYoyXMjg3qJ/
eFwFm8vGrBzgiaz9ufQjpRXxFru1z3jLM2rmZp9W3LaTVbJQ2XftjTpm12eWKhn7Ub5au/eMC0oh
hpG7EEnne9OGdFTvUadeyOWiJmpmNamK58HkSIHGlJ3CrgBwASEWzoUXut9v1cJQUhkioo5aLiuR
HzvC7BEn0c8fC4/zB6sgLnFzRCJEmEhUZqK9dGj2nJfTRROOqFXIGDiMxDzSpXBObYb5GFiqiELE
5Qp8TYzeflhh7zo3gay7Aa179V4pVuRhIb8aFO5Eq6CtI4bShYkkTvv04hhHEQyRPPN9miRrhD+x
Yr8CXIzvn0f1FAa6UxMWwlN7D8aI1v52OMai8l+YIKMGYUgdimKDeavkw0addMUaqfcaZKeqlHwX
uWTCwBNP6uwxxwDQw3f+kdwmlxvZDNz3Qo6IV+Qb6k1osb8MFV9BMdH9kxwpnKmM6UK3kKQSMZN/
b9aeg47tQ2/wZ3YJVMVCoOHXThePUANB7zQII+H1ZjHBkz9cmkoIhsv29f+K+Bx/7sxdseIOAe7O
uBFC7HdspFzNa0a9zzUDPhY2eHJ++sJeyIKhC3NB95w7Ah4m03cU1n7QHrcQdVWTxfEuCKCRwchB
+8me1ATtUzh5+fkB73v485/2DVw/Typ7WOiJm8hsgwYIC5Jfy1Drp3IG5r+/qLLaEcLohuE+lcsU
0X0vUOw/8GPkUE45RlWrU2HdYzg5xuAyl5HqavfoSaOuREgehGyc8ApG5ywwgBmz2jPVDynjVgfb
SVtoIRVt5rbZj9UPqnH9/OPOh1+hHrYXQqeL+KFG73NctivSGbllen3v8WGG/bsBUlfwsjrve39s
PobvW88m6vfmGiNx0ih+vgo1yHChopw6u7BXWzoqdJpcjsIsl/H/88t1C2Q7JioGGw6fqM0ZoQVD
iHUkhlU6M0SsU/TCPd6IAl0UL7plfqb+b1+sFF6nZrUVZgW5RljP2xKcYDWuhzwhdGlQu0+p7oEN
HebaOpQ0quzg2rcdq/g+4gzk0C129Zl3PbuMDeteXjyAXlUR0l1G4LJoXhTB6xs8iNgkkhTuYtif
KxTHcd+bkcPfd+nb/Gl1LoSOtn7K9Dv6WA3dW4u44KOxucvs3dkWKy+zXgQaHMjJL3wiaBVOn3xJ
cgblSr9ddyPkbIjz5PYgaTyXPbo2T5uuMpj5k0H2pdE8iCh2IsZ2cE6ALCiBG5SEmnFdo+HbQFWx
XugQ8qrlHLc9TPwms2Ukkhg5WzOcpe5k/sAGFn8QQV5RILGW4Pin3Zgg25s9SIQWViUQlWGE0EAQ
OjQvz1I8OqWL2m6iXX9Jx94K6eHGc9a0gNvr+gJj2LpILFbhzrwgtP+nQa/0WaHEqQksYhki1wzq
TJ/M9BinWLmH7k0DW8jc9AUyPvKnmcOrxS79XE1sBCzlzOxrDV9MBN4U0c6Ep6x6rCTC1clEJRRS
DJG+nx0I2b7N1uPNCk9xJeXoN7X67o31V31wvsRRtwmpaTDDI6jPJtVzr5n4nTswSXdK+tADDTPp
pj7BkQb9ZYgdCwwz3gOxC3M+CW4XKmKdWEkDI3QP+5VrJ4WMC5Gq+H1fNtZ31443/4Rk3dB4klA+
Vo9zYfFtNFjnUT3dthd+F/pYmw8/Pvh3cJzcE4W3fXZzDoWfhB4P0uQmsxmOw/5SObA5+LjeKtN9
S6McQsHQZM3/qh3k8F1mnfeZ/D4jyXzX3zyYIC0KwHKm0m3OjEoZXLVAkIO079xqjUc8qvXE7JiI
scPyYW5UqlAM/bznZ4shFjD8IEz4RKNqJKhGkA8KVB9mzmLVhFIu+3eWygIuddzBjr2TW547kHV4
P2AGhad6GVTYVw0WMiK2GgLM8BcwR76/zK/BnB7D/yCNi+T5My3aUt/upl+AeSFRnTvzAN1OKfVa
cPx1LSa5Am4nHUMHVMIHwE2Wpx9nS63mkvEeoW7If7qt/wteMRULzmmXmycGEvvYnnqg30gQEx5P
CIgYJL+eWFN3c0AqgWiLeWhdFsJEiK1V7oCQzwiNJv8Od3k4XDkb9Hr+1KhWChaBTfc1xBACihGx
j3bub5u3a08J6OfOTXDbAGBlrDHFYF/RcibNZ9/J3AyCY74wxqui5zGMPgq9oLwflidIXndPRZus
cKcFQx7N+ziGbrjxGTdF8a6vgWc5+7rs9eecAriTsBedkSounkbxikxYnQ5Mz7YnvZkOGO/FQWPt
REvd7W2BnnG022iDqo79kFmFVK12BlvJkX3r3iBE0DzGrgHW/LTw5T1azq5iTv+463JZv+YOQg8Y
HVIrBTPPNIakrbRzKEq6WWSM47h1Lo6EIB/4DyS5KW6Y3s7IDgvpYEzjHTwQ/+5UZQbhZpTVy/XD
QrxH4On3/VDC3nsUbA+id2T/rZreKp/yYAd0W68fQtbMKC5guwGslo1sMEIUTp5fwoL+EqtzFdCS
leZdTf/oRK7L3dknCmWFXjEBf0KiQlOAW93S73tZjpTW3x5zSeWKOz22RcO8tiTt08j6FafsyGIp
8Q9BpQQySGRE7WMyBcouMu9mOIIB25nc2yKC7KNakceQtVJltgY3bODUGXIMKiRzV5Kbp1RvFOaV
iEi6tWnRDeLn41PyAfkG789rnYQ+xSz0Sjb4Z/MU2CHFDWvfsqM+eKqgBNCBulGbqQT4m5810S+f
UB58M8g6Rc5zSS4vC5gDPgRrMtYV5HTpTAIpFIvEg1knTYruDCYSr5AVHZqoXHxvW76Pd9QAojZI
JEdfXNtKNmN8uZ0bZz2pIcDprJR32kMllHUi0voWfUITvzr1/Jl8FGXu9Vln6oG0bt6MdIefT/X4
5OlO2NdZ0ZBLuGdtIIerqWWvhiiGlnXdH1lZQvWkbym0ZRoVeSUyXNlcWKbovGrNjXnoy56BNJSL
RoS4XvpNxiRiOLGk5RNI9wfWZT4miRkN8v0LaRAz5PjCt/NEJjtGGtJNT+oM7JFJyhfW3oyRTlGj
nU4lmuNjugEvqiv3THWGeBXHSaNxWZ3nk4Qo9lG8CqlJ7qTqRi+iuNCfUGdxUGvVS+p8+e1VXIV5
buhKPnSbgDDKqsDSIlMrf4Ekzud19lcXYGfnDW8xxCkobouij4UiZu/Z16RXf+sj/C1HZNMmomYE
Rt1BNS0yITLEK+0PsM8qQtR5z56aOWgjj2NYWJ3q0LicgQVuf+O9YHVQg566O5Qq/4IXevs95NHx
To15ejdnOERma9V1n8h8KnVECJwifZO3E/BlYlcMNyJOM3s0U3cGjmemnrmqaFbJRNq7wHZENZqp
kjlPcVAkEfWzKXRu05/suUEJ5lVAE99mjlls3uZj9dMRSf9gQazNQfkCGwbGa3Z4phNu9xc77OWI
mPnhjqoV9NP2VaXN63YeENx7d0utdurX6trRzfLdpo0zhkrU7N+0j7HMa1pJ3OYN62ui0Xm45DjD
Imy0Aimpu8TMW1S3fcUOeK33n3Jy9Tfd0U0AXdSRFXD/RHC4DRBv1phT3MMglW8+rbGTWmSdNp6s
IH8bLx39ZMAK+56mSLMEMTMSFYhSR/kXkSaoLLQLeoalaX4sZqmCZiKulRsd/fhrS+HNTH5psAAr
7SflIgrfuOMym+Vyias31NdPIm0Fl4dtIwKTKMTpLezaKfdy2x7YgZKCw93uusmTfQlCKH1wBIE+
/dx+D5cMUTG9rrayBEumEwrExNvTJKgbYS84vmb8dzfPlZLI2/QiEAnOp1kgwbA/RP4HocN2PBGf
XHNbGxMf3ODLiJtnF7k/rOuEhCOCWvQUrw091BmEeJKp36Py5v0jJoGcbsIIC8xwwF11znflTtee
/VA9uJiuwpIDXLIXjs7cuK+iLmLJvzHFkOzvmUMbl0+2JXhppNSA/qr5o5g1yGb3+vJGAhQFwhuk
CAk0UG4PjLnML4QHSHT85LSzpyKb7jWrODhIdkbGx4LiQ7C7vAZTaSHTCd/Vws7WJUtYYymRV2qz
8vTd6OvDKiqbLpAPEq8zeY3AU/hHObRRFlLslGIjL7oBxwCpaiq8jVRkW6ujcz7Pagftl9wxsojE
oC5frUzj1WV8J0QlRDNXDuvbxhX8DYIDLq9SyLcWLLsdLZ5+Enmr3fVhVC+FFkPuMsfQwHA9BcLC
enX7bBpcpNhzyJWTpKJkLDvoX5FYPN39LLOuz6tjOB5b8Yr1TStTZ1Ue+fDibYIK106WowrxH+xn
Y+80BWKqAGPNtQfxwhVgQBl+7EYJ5lgA+QrOePlWdo6Zas2xY+D7JbB235kaRLRV7nSKYJfSF1Ax
I+5gGvCxrXahqCBANzdeDJszJzNeHMd8tdPTgLZF78nS0hIIFd7ouzogJMhC0APd2PCq1x6Msjjb
YXuOC38PonRa2xlAtUeWVwLMTwo8D5OLALN3rJQpVq/Dzu4jgWAGoi3QIGJ3yi8hkCrHFyIgOc38
kXxHXJ61jcggJrJeO3N5g3+04Rou/j8IUQ4+E50fSr1+ZcK1EC1Ryz0bcGqCax2YIlHgtblIRwg3
sHPMblDekac9yyk0wOfsTVrznfw54gq72BLVhNgi8/ql0HFNez1/+2UWU6lcoBbK4i+/wH4JV0+g
1JPdDOR0AmT15vcLfO+kfm6q9p9AZ/kCF1+duIYI8kH9c/HvNZM8GCrGHThDo/8UN9JRgXjTaH/Y
/mDCM35nOSR/hAKG7cIeXMRfNM6dgm52Lp543NAaznQ3PVsHQPVqAw/OmYSQ1KVuHtYKuKAxXUVM
/KvASKcQoft6e1D6moh902CbcyVh/PjlrduSPVMeOnd1SDv572BvficB8NZ41bA4X5hjuWsuAkBJ
cHPPIEprLqlnlN2VLlDzOsMllzF0FQ0VyQ6Il7aSalxl7EM0yf1rFz/GaVYScvWOdEy0NLiqfCiY
6/ji8yOJLCetHwdA/V281NOdEaUZ7vXucNRXzTlnaVfqKVsEP0v2b7JtwCXFlxzfzAlXByd3AF9K
/EmJyhkfpcBEQPWxxGTWqx2TSIWvlhkIXABBrLDiDqYa4lpOmRyX4ERnXhKCDywhwTt84dFuVx+r
k3RsC6IDKO0d+uEm3saoe5AkwwJNkB46Z5x6giLvZPqsjmzLsBYwheCedw2kKyOKk8OscdyETC+m
OAKh7FYL6/IZu96rr51Soxtc7iuTRDrQm3z2vhCYzJiOVDzbmZg+SimULhU2j7vPDZOPgyC5laCx
BCujJ/gqNmbLPSpFKm2Q+vcO8ZvgFf7DTHA+C2XuqtjnJpXQ/w2MuEJOgDnMPoccpRnX2Lu8AvdC
HQickpfKEkewT8m4cW9129MDI/YwJxPHjJxElC5lMoMC6UQMWOl70BJ4QKOw4+cDaWwWwQkRsiev
WMsdWXCfkPHRrlgKW7seZMP5iQag3XmEKoopzrmbBiCZn2X9roXclrM/XPb+O5/JVLXdeFicKdR6
Hm7C5PZIRoa7aeD2kCiA4v2Y6pg5innpIfTM/zNodxcap0951P1ZJRQG8CDEWNcN7SfOAZPijaJr
JL0gi4EadoY6oUfOKB2wMd/xZlRl3sjnHo0FyTsuPgcI3HAXlB1vI5hRW9pHC4bOX/BsaRLsHfOy
nePCHoPpNg6WYr/exKTOsA4KHnCWi8ZDWNdSjwIUClZ7G8v03J2AnNdoVUp6eOweePZyvqoIrkff
lTjL/s+j1ejQoliquJOCaJRVtd0rjL7o3lUThWVdocJ+ANcM86qMbRIrEOjUmL4a/mQUYdBeKRKv
d0MHzqDCuvavQbaLYVFQA2t4wws6f3oLpi+IU4bVPiLKeg7DZwzmmhBauTxEXPnIZXqmvS6Xujwq
48DXrD14lNFUiJXI/YQ/vMcHXPI8qw+UZTZfrM/Yx5JbH8jChnJ7kdtHRYnKBsVo3UteINeslJHN
AY89RBJ8GOpdtVZ5nj1jKvSaz4nTbbvQBjYw0uBSZE3x1AxiKCGsChvCAUD9csuOpTDQiQmTEbHW
DK/MfDaQOoxR+nEPGEL6OsjpzDVElgXq+iiigx4jfW14HkCAAA9+VtLOX0EGuzYTM3viPUSxHNZ+
9rocKj7kgzqFaT57U7slUvlPZreCeah9Xq3K/N+fNnA4ACNYgr13vXxgT9Xrk4BkwholmTkPox4Y
1V4XvoRe6NmYrBGV6AaBNGXow/6f1tnDH/CHMEYW3krBBlNhMD8xVLzNTYupuICYvVEdLjgwmFHt
6TXYi6yTKI3DsAryeEwL53mx++Bvj/0ghoCcltpbW8wyeR/2eB6Z9axeufSeGXv0VFfgapoDLE5S
oIwRinOT4uKgdieqPLo4L9sNVSVRtDggg6Eha6UieU71kT3HnCyyzt/e1ip/65pOUUE8ycUJ6XLT
J7vFRU0hAYpfjCZ8+ZRYPF4cZs+jTolLeIl0ORi0adwcshgu99WtjgSW62GLES58MZvJphuAhZVI
PhQZSYVkPZkezPulQcbUrwGSPSu4jdjc9rA0iTUzP/7TPCUWc75CgGLh8N7u+jNwnN2z4Dd0Wvbp
OK2RkjXZgq4Ft2DU77fVrLTgvaO3zWkitgdR3y2KnsMOb9apQOONRylW+dKAFfE6MLSYyNxY1XhJ
xrDBjoxnUIRE/H8VDbKQl/ALWO3nQburm/g5YvnAqyfjNEuXYtCU/FQJu3PqUji1KWz8/9MP0JjY
Am/PBXlRemZ+wF402pyuWKlLltBMWlw7/B5nXVFl72vHtrRhXAfpju7vF9EZsQWw9dFqgUlC3Xd4
U2TYnapncUUYAX96jcPb817dlZguQ9EOZs9Ea7+tRo/IlG2HIsXBEAKkp+EgzMdGV6ln647Ha5fp
/WIpdo0vmvP48w2jr8Xs2vDfzhQoNtPI5WqIsxoCA1MosJyftQEwX/QCjG6Gt+Cu0sassR0LUyoT
9dgnsGk+eq54kdl5qmFEbQMwqsWel5u0ErFUigtFkoC5KQCDxiIeRs80jW8uNW882DQeWXiUd5s8
SZ+fiQs1lJrfmEra/jt7X3sjo3oDcM5NTmowuMIgUHlZOCeqkXq0HxxVL8OHzNkgwlI/LBl6rCds
htM9FwAguIKTd06pWNBlpvbJ6Oocy5YgYT7Q2mWL9CsN4NUphuGUiJsuKYlyAQFmMWeal4o2eede
UDhWCegPdVdxImuzdWibJnH7Kw35U/9CKnriJVqjJIqmo6mb8K8j6FM4C0cIz4lwtUTlNUmCd73Q
/lixJeUeHFm/SVGHCvot+xZscsG1mQKaYWphzBBdTSJgmoKM7AyInHVWgYdAkgERPAh30Yf0sdMq
PZxYy9mfn1qob1wERF8Q3LE8ie9K5d4+Mm9LYDh+jD8dxuujF7ttoIO3J7WTgACyesASCielRTgA
WtQxt7Shi7e413waCGhkY1MebRSwHLy0I8AUW/UG1UWM6Zda+mkqQTXjgEx89AQXJGwpjmVjpVHo
P2/207Vy+g3Qvri8x/21AVIkEjj+/fH+pH0vkjt8q/+i4MmjO9mYQBZDiM0SNhQE9UXh/8YSf1gH
5MnZSE3J3PEt9hfrQ/VyFT3KWaa/S0ykpijKGafUWBGIGS6Taie0RhbkMyMt49at0Ci1q/nxNY1J
XS7nVcGfgVcRXcf9aKTZMfydE/T/keC20D6dD2M8YnsZAkqxYJNeQV7OT6+s93fJKSDmoZFsxg2j
KCY4wqEKLRAZUc8DGXjRgcDBTmE/kHMvoPmJ7rVF3EUuQeuonyE0cXrZ5z6bJ778gu6pWsrtK/p1
Hdd/MGz3fpU1xiqN22mkZKSN8Bnb6g138DchF+NmYTh5I7+i/I4SMAwCxNZH5i+h0LX+p1xfNcdx
5vGE/z9FA+Q+i7KpvasU1hw7GyRQiUwlPqfzKIeQV4h+i5RBOpKWEBO3IeXBvsK9NHnTHpEXuJvb
iL/+aZf7ty2ZY/nh5mEL9PZ/+2rld15kfy8ampLs6Z3g9BcJ5llhQhgNe8uq6cCiv8jtWTMxD2KV
xV41bHzf1GUKuOL8K/mnxwm8r6A+T13wdq9Q0zlcT7/iJouy4W4bakkkl4YfvNyiwTtzbN9yL00N
EfTScahqeJD1nNDYkGH+09T4GZZYrA4ITvij+Tw+Th+GHBvW4QQqSHF4nOnoellnDjBFu7jOvbny
KZF+dRTaIPqKw+M9xdhvER2RQ+vBC9IeC2/4QI/ygVRNiA97U0v2p5RusI0H4GgxAc7q8CyZJfuF
3R4tvRs/sDO2O3i0TAafEin6fNjzAJ7i88N+d+zm6ab7Grhr6j6ZG4sXcKKL2Sz9CyqBI4ULuTWS
QggftPhaOrnJrEbY1U5nJyxJ4HB1rLV8fxmjSHkuX8zHv9zdqBGjB/r1fwHhxd44rggq7q6Q3xEl
SYuVbniCS6DwkVhzIfBPhxdf3VlL7g50P/yLZi01yTiVgOO23aPek/WEl5heC56ZDjB2GsmI2MTk
g6IFdvg0xeupwt9j9sCO2+DOL3eSFJpwV68JD951XchgsR6inLpr7VCjRpPXpzxm+nLjkOZoe/Dt
0m/41dgQePEEEj9hMmpcAa85kuZS9DQ/dmF+Kx3+S9RARAqn1J9Oc2lFSgmHV6ChFswp2TlkER0l
BDwrrI45ZMVRiYtCU0LIBjsQVPNACrWOPaqr0S8e5pSfOXFrFF0vit6jjWyqKO/vb3eGdmJiLiYL
mTVQLmJ9hrqvfSRkGlIYTCs9s6GyxrUkwCvMUrpRwup6iwVlPkC4dEIoVfomjk7gTp0xXyEEIbS1
4FaGk4zOlBqQPGJ6JaN/Gk43x8PtWzkVzXf1DzB4OVWTXlJDplQ0nFZpr5K/K4UsUAK0TDij62Lo
eKw0UyTX2wpxKAlc+opdFbJC+idSTlSNm7ouL3HfxwZ8HIrjz+UU9wkqHJYmeCc9MW5uYSEDA3Ei
hEFyuLCWYWvvr6gUE/OI4re0ACxb1wu9XdnYqFdsm9RVTeVhl309u2baOnfp8ofG0dzSq5l21g8/
9FaKAGtykC0c7osi+ofktgylJycv7YUv0BqRFBSVuNOC5/lGgkOAf7R0Qg6f/3SzEcTpjFK2HMW3
cqWiXoQuX4ZnkaVwHzxktkExd3oHt8Muan1zZ4SZmpTnJAL7ZNEZZubzoo99Esisoc2ZnxSqAuch
J/HCLoz5yzrIiGLhP9V63imjdbb2Zp1sJcjy4cVOycjFr9aG2rAEqBgqh6HlgETQwuH31uH9dgHL
DEdwkER2QDOirPSviGcoTmIGIn6BzUlJqwDq6awFascWpG53CCmFFxPGhIYokLHpBX8bpduX7TgX
py45Ji0tlRR407y1N0ZT7YT66Hmy5yuL5aRi2dFPgUva9XSEVxRckMmLwSxstA6b3M1yJSo7ereQ
xiqH3uLw7g5GU50oT1CldazbopMEtbsxCYR67HOV8YgVSfA6cQL3VBKF7xkfO6xs7eEcrr3E9sPs
3IwFNGFy8SUdfARVvx6hObbnXWjZvEggEUdfiAegnIrpuYcp+vHM1KO05cLTBcFFpkwmEc/aSFJ0
Oj1lXCc6uvO/ccI6IXfgcVjkelz4vpN2YBPDm+VF7R0wYCKEOrko5mEAD31BNbHDo6PydGjSoGtM
hu0QDXNplQwEtZDsoFtJpyoeVwTJDvPaV7f4lFMTCw+7JytmGBIHXxDcqWdVT4ByWAnYDInsrWp3
e584s+cHCb5JXYQVHiSevEIIg0ox8AHs7YYOTezKvbuYfMHo6CF7aKoO4zZk0SoHEpx1aBzMzD1c
pbHHk+z6yL66AVeor/iCA6xGSl0d5yDbZQ0YGn2R2grTorVuDZYNQcb4xYnYG5/wh0QdWYdSDDYb
iCFdwNLwCOp3H3RSp3EF0JLMPmQ6fuu66CbmCdSRx9awc2iu3AiiJwJP7UZbBrzOWTN35cMe/Rqw
O7BDOil9UaPcfdDym7aCiagRzaqWjsT1fP7dd6vDcNGTe+PiZrwMRUlhYz7MdaX7Oq1z+ZbUEsr8
WWvM37q2OMJsFxptr9cVxR+zevicvP/TOz7QvByYIcPyFteYeHqq5yB9YMs+ffkI69EzBQ7XzwB9
QQY5MgsnmAIQ4M1R3fbhTwwz+QPNyczciayG8bAirbEe2GvKgPiFKVOps3fsjfXbi5tbPyteBHbW
KS8y349JCxatI9ck7eu/c891neL1tI0MdsjbquNQ7TUtUvntR8lpEJWYTSzMgGYnkOeIhu31sTHs
14pYHgSiU/Rr34h05PHPfowq2wGN3G96GrV/eEsTb03JvF68wSfE1pz516f+43+nOj7xeRTVK9lh
ZdfkZYe2DNfJgHO7SyxWkt6s/mQo0XqRFVWEVfcnVbpjPPvEHIi07JFCFdNHXiZIYXOr4DOHv52N
6XM1AEAN07KkiP2WJtX/RCcOFCmcvopdNzL6D6HJH4XBkYDvQi+do01ue0lSIyTDZnCTWZUqQDYi
8vF+81RyzYZOQZrovhKQVkn0AgHwJIj2JB0X9YiNFE2SPjhzBoMEpJTOoC1fsyeE97BHZK5iL8X9
vtdesPgAfWAsKU7aNEyPQBXjG27SNOGfJaX5aurWBxBvvCHZ4wLkvHs3zjkSHeF+RN7u5tMsVTov
WF5X0ZPSRBjDGm6yATcjJjLuXIMGTwwdtc5b9aH84E1qiQMfGr2UOT6ocHXJF2PU8uVta8lFl6OC
6w/VXc6dTw52xvqtya5ezDwfv41S6IGaTqMOCs6yolHLuTcTk638jLuWcu6Cyi3MoRRXpaEOVJAX
BZ+mZlMvxJEsoQijg+zuThMWZ1Hobfs/oFo8sKyTQq7O5FgvFhpzuYzZtflcJwTvrCT0X5XgxvRd
ljHQuzTpQlJPHS3OknMJoHauAp4Oxse/F+wFNxZP4c/9Yl/0kalHWY0grJJ1OEtWMJgd0Y9hXmm3
U5coP8o1CpIIKJtWrKQ95Iy4snYxM8RARFufd5GIL29Y1TymLPp4bbnWvU6i7wJ41ciLj0VscMfN
Wb5OKzI/x+xMNsbfy5v6VRegFcBtA4fi3H8Ec5G3kSXfIQ6c71ZhBTShqqnDt1QHhWvLE4cbZCJ/
u2cNpZA3lUmJOYABZRmZmZO3F+D73t2l81UuxWL6tF2CZF51Q6W4Sq1tk0ZZcV2eGnSJ8Bx9mn8b
5DQpjcrh4ecE6h1BLUFH5tIuBr0ixMFmKSXC/R6kMRVBLquLoXtpFDQBh1uctcLYZE5VxIQqIYMD
buT81kNLBPsn2C6CF6uVM5D2vSzB9cmyvZERDh4OPvU3Lwvag5msB4YV2N5iLKIOrEqMvIZKvkuG
9lQu4gphyM8aCyLr/LbhkNJv/pIPvAr1yiX9eEWdc0b3FTXySll9N8OKeGqrfASM2qzEKRHXgyN1
R3VItP0mLDSIkMs8T2JpQWoPjzbggX554kHnSFuQawex8J4iZFLSzbJ9sx7O3sXYLSHUf6QyjIGK
L3WiwKcnJr7PiLVK2mKGeUuMio4zC09Pu6T3CvAkhxbsQsPyCE5W9msy4mqDTvzdfwcMTir32XqS
415okyynctWX5CpDYwLgRfoLRWytCDcFNse4SxT0uOm167fUllfipW3zswiWc9XaHvYXwo6kYiYc
FkJyu3GgSyXE+nkp2aQV81naeHSS8F35AkdkVMp5ZDT7F0gL3i9hnGZOzc5j2hEnGKj3QRn7RsGj
lDSbDlThNFbbO7p/Kmsuh4NKA6BTK69E+mdLMK1SXOZvYJTtZZeSuuqKbLGzspDfhmOShiGPOytw
d6UZKAbXLfdVr5JVMCJU49dqFUIe6dYB2sPHWtBulkFClv3WyrHHHTC19+RczOGumf7EZhWrrQjl
MGcmCRuymKzF+cmc9Sa8KChS00laMpW5qkDT6baNnd7AU11rz0q1p0wiNutINHOVDqMdNV11f9th
8Z2h7TJDYpIPiSgD2ahucm3Q9aZt4ycsYSm/0gj6n1ZSnzFpPncYyQQRdHn6dg0kuYGkBF+wHTAZ
YEUMy5wdZ07RZpzSC61heeqRwId0VBZSXi8pOo6+nH6xm1S+oehKLA3ycJStGvhZYqBkhYpuAeov
2pyrblkW/zfLEHp7aPkHhsruu+Px393R32s6nTB/l1MZ+koMo2cBMbnM6waGk/lgpS5k4IbD1yco
cVOKKtjRZL6nTZzkofHppLOOEqpHjajCqhAvgKuz3D57ABkbWajoiNfOn33hLR1+8eOSz3pIAHKQ
jNmsoZbTlJtGDDB4jOeDfYAsx8VpPXSieyVyTwSLiqouSon5BhCsVCYUhWA2sTbokw/gT6QBSW2E
xc+0JhfmZelw2Cn8CXIoNs0+OTDVpN7449DaMeh6pbzROnmmZQQqdq/bOoiLkXkcAhmnGdrsRPat
OqhBy/jKoHluzmeVhjmxdtnebwh0PmM5nhtGuFFlCRWiVGbwef0zBubXLQ0snevh3j8LLZUT8IUJ
HxUVNwSKPbKCf893k/WQcp6Ri5KZEJEuUFpQqrySCTvdvUx11waNL4TED8nu7xzqhiYaJfNwTBb7
i5FcVAuYo1/kmH5LleDcSpqC6G2xw0YtoIIDRTnAG/cAl8KiiHRCi+rgySWkzWyLVTKuvs16td0w
nwwSgSNiKccGjCH5SPiVged6Ui3SRD2u0MNBMVnjiB4T6dQQf/wReZqvDkTDsepDIYmElt6tlaFx
uNsc3Txbp/6vpNhl/zR+YVEXp/PHXult6O41pgJOjbGUm4OZmLaFzmL8uLhUBQjl/LZrGEBtL1M/
02v+Bvt8VefUc7PORKK2xaR3M78RM8Cm4yRZ6VfrSfU3r6OKs9ukC9ngYhYVc5Dunh4KKR8xz1Gc
ikNnY3lE4X8m6kCUi0+np/oY+40aCd5yFSUNplfUu5v3Qz/ZZOGY7f67iW70K/gSve+ZPDMMsF9p
n14V8LLSOHE12oQezvtYMmrni4s3InFPg4flTI7IYd6VVQ1ijK/pVr+0Gq2oMd8hXXp2peQtsE4m
gl/cZV7MA9j6TCrzCasY1Jl8B0Ne1yBy3xQ7rvYAoMnmwZjrKBUZ+6NAyGyMTFTNVtpr42Q48w1r
a5CJv72I8VXY75pS0jGIOVjoxAESvc2d7f2qICbtuE9HT+Pbu4AC8tFI8JvuS490isfyBGUuYk9U
E9hZIRnr75PP2sMckO+cD2/LglcaLZaNz+EyU/t/vl0JeY2qCu7RmT1u/7CohQob5z6J5ldbEr6T
/KBQ1jRUQFRID9nm3iHvNOhXcmtiMCcWbiEZV0gVSaWM87RFF4W04Cs47qLeG8XRcieFiX6hH46B
DHmd/0+utBAs6kS27RpFY9lAygQxxgqmDDtwa1xyQLY/SALnxNNdgs+KJn8cP9rkNXnxzPXVb0nX
z7NZFV2S6oYa/0qPuQR7U0kLSJH6vJPAH+zmgKirWpsAKnTiIOMg/ErL3XtRiNxadkFXPtr1EQhe
rBqe7II+O3uBDCPArIhixoQT7cYVR8W8cz1WSd9kCgBtDGL6ew6luORlc6m2VvUrs5/Vo5syCFv1
bH2Nw69nmCKzfayh3Lb7eiHVxPhNex4IvOhFo02HH88ehpqzXiMRJZKpZc84RSDl7oR6pqaWEl7z
Xp4oi/55NEu5LjtvMHEDPeHnMYn2ipwQVYXHU8D+KSUb/JReDHHYo/NwmLibW9D4Mp2q003ihUIB
INfHbsY2hIgPzglTHUDXBTMy6BP7dz6DVwSpV7scvxb1bQ6AHIlsn795J0a3WngaThOv8WuiT8Gx
fzBa7sB6uqCGEdW5kktgCfG3BJryDK0srKoW4aJcAzRhOyc+6Qgnl+UMk+GWHmf9hgj01ixQVQXs
BCOEQ7GFG9fZXIjcbnr6tzqA4fqerDV1JRb1Kp93DJYocm59W23qVMo66v9qhgIMgI+nFa+t/hEa
/IhyIZpyQlxXK4W1Lbu6uQrOyVdLGpusfc2FpKqOCB74TUyCuyRnhOwUV/A1+vOm1LDbKmIyK5NS
bqOBKU97tvaAGhBt0/oRFapt8NeUZkNGJXjLFu0soopLenXh1ppgyMglhxXbKpnfZ//ezhbMOmo0
tOrKr/4+fJTXvIi8ijQru6SfeLkEahWBT7oLKZdf2kGrTzKbeue40TY55BkFb7yaX+uMuvzuQY4P
Uch0nWNncdMxBCnnvI38ZovvXyppu/ywPHgWqdk5tRohRL14Vzij7rS8glVztusCfyjAxnvkm4cN
6TueqPsBzX4zdt4DZ5yI+ayQabhEBkLKh5Zdu0H2OA7KxU1E/sc8dIbI1hzllfrxaGEhGPgkhNWA
S01FPaWQCngfMJgutiwESPWuTWnkumXGMmJRXxAF5OjWu3zEE8FujNKbdpS81a6A+kIDQBFrX5Ke
GOACo0kmV1nDcCEYZjXVbCYzOvoRHASe+q9VbSCWTLLV4CxiUwI9q2QMwBPRYxBI0rtpBZJdZ7TI
WI6h0fWc1BnuYKsx1ECrQBX1KIuBAgQnF/cUjsALY8cBK+Iv4853juGKVx7wcFTQuHZUo1s+We+f
/5HDkB1MF29szRBg35H7Ij/LzaK6UCR7LkMNvHQDIjPrcSEijxDdj8x9aXjBBknmsKZ2egb69MuU
2n5TkVKLIHls2OmLHW7AjNrBzqFblQp81HZ2clfOgk3A388kunXt2Xj4o+s1tgYK3jFmVehrQD5a
BhMuUhDue4aPgCCse+5gLM6CWPcrn6ALX3IXQ2XHTKGsbYuICjoynOwm8TQvIkRlQYRHFkMb3yvp
YO96kz+N7rlb+73sXgDD7KBb/DZyR31R2PrbdY1DDbn6uXjILJQ6biYb7Z5AG4/57PRAZJNSLjJr
orZBjZ89NY3HGjyB3fZPZVqdUZHZVS2jY/20rdkEdmcK7i8Ikx23H0yc47dF9ZlTzCTZ8AWAzFrQ
hukrw1nNE4V2P2q0Oub23GC47fmobx7kX6YA+YaDeBRNCa4pKEWDVwHWp4wTpUsjyuuffUbwvcH6
aBGM3Q5zyqwLaYFvSQXOh8jw3W6Q1MMjMUyrvvRZMzJhOthW0HyVtUGVtyHUvHffqMfGZ+I3wHFB
jy7LR78Z/AOrt208Ln30P7iFF8AnyJJTyR/NJCs9vyykt0caSnIottfMBlE7RxWYD7OU9YqjqoIF
F6dbP2WPh2GTxZE2ytpdR25AfGnzKFjgBJItFfnjsZS5Q0egDxDPtzhqAv3AixWI65qFjdeqidYg
kuXHnCS9TWGrk6FWV0HmLP/71tat9277Cy/43136Q+VlQuzTUrCkxE2YKwto5uERitiwQrStDe9X
mSPB64Z08E6vAN2uF8uBhYbZqPpccXi98YaClFmG31UKUwZZuShtwGsIi3dmZn415J1AhdlsJ4lP
i3eLgDfZkwq+XGfGPHSpBmFpZO65cJpQrwKhfQgaRiIaN7Xakwe+hiBX823BwOuZOIvwQ/ktQ1Bm
arozAMm3ERmoXEVqbiycLloKUzL3g4FSwNTPjFAKjJMw1O4fiRKgJ3lTZY0jlNqUttE11BRwtPpE
s/rRg5sm/oYzcqLz1t2h8MG+9SspXTos5g7RMcR3p9x5DtVhLqmrJW4T07EpR+67AQ2YDFmKBt/l
QO7YwDfxAtyTWx8UZ/MNFNrPIFdKBTA3OnutZH7+Oy1wAyx220hDLyFZ5rJi1xf4g+eapoG/9rgP
bA8ANiJXTnS7JfJhyJKaBtmskdb3LMDNM2nA/wI26CblCvRIKsW9Y1qe00r81jAdhxVJ2RIzcUeQ
19pYkRC7tB1TGppJWT1eZm/c7+ADAaqAsoYlAdvxaU43bSjZ0VvAtEIW0s5eqmHdDFrQ+9K2Shhy
iaAma+MHHcF643mN4dN+jxnLTNzrvif9nH4LIkQvegh3F1PugTDjEH+4ZUvdx83RWL22kSFosKM+
k/3Gn694C/Ma6KuFrFUb+5wG046gh1GXiE3B2OieuvK15R1YbtdCaQglkp5FoBXglg71nbDeoSxN
iFNh6H0crCGn3tLebaNUzGqgAJYdx0v5L18SmMr5tAC2yGh2mzJXWKWrc6BbRCv11JbLitA7qmGD
pwMlwW8Hj1ZBdR6jQXKgsMCUmFbrkSShvOZ8hAJcrY/gnnilLar85hXf5cKdGxbsBszUICu8l/H3
PaC1+tfvrOSjUwA2k8Q/uye71rQJCVrsOKRJRVMB7H7vSEbk+IvUosOU3ZT0LM5+Vhjr6j978sOe
sYuvdEjbF9EVQiecaEo/vbSqc/mXDTrZLF2h4/DDHLZheVv11iPZOWOT2I2JGysGIERK/VNkkQw+
wuWQmSI1hFS9EFRjbuL5Y+iZFRKfPS3yGjh3mj+Xquoc3HxMOunaTYTzX92OVcMIoJVPEOFp31Ka
VI04AF4hNTspP5PxWyUnSE5o/eq/CNxNYaojdRSf6tM2khyBwn9OIK50Oq+ZXGMqAyO0MrhBQIFM
GGVMUp0gV2/afKCi9zxEUCBcQ6+SsLTCa4He65yvR37sx1EXsksqSPaA3X9t7egP8jHWjGHIYBAU
uElgZOAA5OWtMOYyBiIFnYAAAAZRJoJDNu2PhzXU2yl1ny5HTohaZziJk1vAkz3kcnf31pZeQqbV
FLLd5DqSrVln9nmpXtiKLO9w5Yf5UrkKwz4o8Oo0VJlmwLLz2F87Ed3VCZ9hkHtK2CJqGMx0rImB
3Ne8Xfbb3Jd/Can/qr3WU4MTdMfXj5fYzynSsxRt0XD0FxIfWHVDroKRlXDTl1SqxSmW/OH2IRfD
zx8e2HkCUF0txva7eMzrthwB3WVu5jJKtpvdMvaouvwFJHBWQXQk3zKId53D21lVZ3eAImqNvaWm
zGiFpg3FEworYpL3FdLh929OmvSDwYUGatmCxSijafQCx3Yf70EdoIvGW0Z/7RD+Dxtyyyqlk3Al
8u9fLYiMbF8ifoo0wFPPjsz66f3eK0Qjqho/UZBSfDLMZqS0PfairxfvG5VuoyfygueRsuUuVIu0
ETyt5YxA0qEbUn/0JnTco0lY9XejsHdkta6lz2IG7lTgpeBpWUVm5J8xRU53qBvcuojJ2bo9dXtl
12XWXRlK8rpsz44v2F2ROTnfzTk/nHSR5PwqzdGmdJkl2fkgJkR+fMbxposISmtgiuN89TqI0Tit
ijjVnnw02oMRLZcnLh9sitL6bk6c2AZuubz/HjGX27xDyIXX+O42MIvOaTfN+zfCr9OJuQyIS0Oo
GzxE8CPV8rPufFnXUCrNl1v/dmHf/AmKbgRQC/XWykryH8bXU4ZrqnnO0+kmsC7IFWXLi86ycRjB
Al7NXRJ5yXJdQqSWHSMv3jciyPScga2pFEmWmzBxTcqN+mY3CIbgWQkm+UaWkuR2GwY9f1EmWv8G
RjdFelk7RNDfQmjZfRY67VL+7PxNSyQ8jx2iiBNoG+Aywh8js88iPCL3qlp36YoP5Sx6egr1yV+c
PVW7Ii98fraJ6mgwyCndjajGzhH/zVWXeeM1Ju190FLxKihqxS9jvwJNgmvUCKoXJhCfBQ3vM6ti
CzrGHUmMQFeDoQBWYdJR923glUnkuOvbiJLUOxwn7VbRwLKTzzKuDNRn0l75Cl+WQ2wAK5a8RBcS
7+vfdQsShQ1brxNrZTDMy8U+zr60dzc7/Zu+SletrP1x2/tYqatCxCxabg8CbSljWoVvHLbO374k
pilo+5hMYSSHMF9FkrXTjK5ZAogaRE0p4poYxSaRoHGBIw99QqFo8u22v0WxUzdkdtD4BNH3fdju
vgVweJBUT/ud/0ofvuzZBkmRPjYg2fADQrwOmFazTJ5x+Km6kN5dkmQurvTIpQSmMFFMqoQr0e/u
i2+7DJGfA+ntF77LAah5H+bYJQOGnNweM5ICEKYvKmXx9huw8GWr2LHomzCLkti/MKN3sF84Woxq
ek+6yKn2oX0L8ZbCx56RlCv1wwgfGTnSZcKEsJ0Fvk5hRes+ZxLmo4zCq2MMk7Gc6Q11cIuZb9iI
twG8+0qge9unMNgz5uHAUGF4eAjD8zGoA/D6f3ortIAjjCCCnJkd4q2rYPcja6xpRvESc9Inmm7H
TpYFMWVmEqrT33YUmyJNScsi7xbPdXULqY9DiaGW2YfFFvTLg5aacWQ+/t2KmnDRwh7wpPEWG8bk
mDZL6nkGZOC+lPTnlPhPTQeJ+mWFXtTXnko2Bff3SYpkrXyNj1kPSwL8rGJR+npnxO0NvjPofepa
bJlKgwsxPUM6blhDqj7INAPWL511sxn6CC6DVT0VfYYJvEWWCsSgnlWM31753gnRb6GmByce/5vW
gL+zcckbHnMOKWajO5EJKix9aqVaXaKJtHocfb35oV0Xya0uF8YUTCRJnqHtU4M7yEP0s+hBILTa
3kY2Kev8SVeZJk2E8RIdakC1iB4OyFbE+MjHcf4at5dPL0YktLYATXZGKHv6aeqGhFpwBzmL1vFv
DA41nWyBctSSgz5wMWUQRWf6Md6J5IkGqvBSuqFqTktu3GYdPPHEVjFxUxZa6t7X0FhuS5+ncids
w2ZE+Lfs16lVNtGkfouV+1Imec3Fu5hn66kucKddvWtuPCkS0a5Bk9ojEpztZ5kVgXpK1ayhLSE1
/iW43X0R0YH1NN2iDqcpwJhM/d4ixwHqA9LLTgxEDpTVa6jD8Xg7aUiRmUt1L/+CbL6hwp6RE0kA
aHMnMW7SmnuQ/vgX+WvGEnahIBls76+FwhKoG7Sc39KyLd+YMPT4UupkG9JhN/c+tIRamneh2wN4
pcRS/nkJ1lCQkJv/7rrNBsgRUDopkPpXo8uoqEo6rJgdhQcPx+ITSzbTtXttBiqQBrM9Qc0GbBA2
al8Ucw0dpbVMQdVfT22a9zAp1LRO1JPUULZubqRymPwd37wusbQpvfoCgh6oZv3Kv9lnHRgmcQZU
keztSLU8JKnhX8Djn3Nmrn6qnrJq3j/Z6Gcd7nymg5BL2sg7t4eAC5yDc5kdNVpY37jVgfQISGT2
be8R+HjVvOI2rrRNy056Z/vbWQselgnYWVWhhxOH0m07VfKXkY5qhiYQnS8jyMKYb5iB0SC3HEFJ
1urOOJi1SDA+DHbuW5vCaEEEVdPMYF4+0sNNfmx0AUrihb/7a+iF5XABlPgq+S7a0t+nGOgzIh2x
R5uOY0yVv1vJPUAqYwLOBod/OxT/0q5LKwRNFFi73Xw90pWNRjt4mYSRD6uMRVTQ54HKGJCF24hC
/GIhy1ImJ6WwQVsmdVf7HJVjYbKCnQPqYrwC294ued3PVh0Zu09k3cCwiyoht22J2u4+K9j4YQOp
bv1fkF4jW27MwfWZA99i9Hno3D4Kg9rJI80/uMDHx0jbpB9ezx1vvMbD7sVnwyeVHIq7gLgTk+Hc
t3qCt8hZeWHhNHmHBJB4i8OtirkYVp4k+gi/v7WBoySLxVWH7nU5/8ML7kDH5nLv/IS3oeONftW2
75OzEzwT9AjsvDQ5jn7gck32PfQ4Se4TS9qI1HBCNCEOuBjaPxrLjX1ht2OJQEtK7fDGFpcGNmmT
o1P0esGdq34HMnyRf/NKXqxznSScmaLiQb+fHyR2z0rqvBUoaRiytFkiuqSf7CTTmzZcI3makrT7
7kDtS6Me5HJBqkZ8Asx4PiPvJdVZCWphrQtkpdrPAh7MPQmikR7l22uqLhhBVnomKznpHu+oJT/M
I8O9K5bnCpjIQHeSdt5fd/jlx/+c8cxM3Jo47HSULOoh+7HXHSlp5e5pcQpeDy2Lc/mdy7rnmS8d
Z/3yhVUOqEsfhu90IXQvOEo8TVIeRj3SZQdaEY1gFQc6l1s/UCW68/1p71an9cQgHQMfWk77jdH0
3sEudnUPbzWhp1uktsn41cgglB+egl2K7jyz0hOrUd/0EjDyUGmMFIRcVSVMmyUtixQ8XMdvZizE
AO2Z6sDX0X7/WyMSxpJvruzOriaV7LkDLcTT0L77SgvvqZiwJzCCdiIjpo/QUCFf1L/2kK6QgD9J
+iTTCtpdSk8ucRoHsohFWSEL8sjQb/mcigyXNh8+tCAGN9qm2h5FJFxdDsXL42j8GXn1wm/79m77
t0el7b9AJXpOmu5iF94GrBjxU4hXHWXC+Q2l4N7equLTp8poN0nGNYlYrNhmdZNvqw/8ZytCE8ow
4R5ZxC4DF1BFF1TGTsRar87ZOby3o2L/IysoflygQ0ZS/4VxFCloaz/Bo1yyjMlfWMXW7J7Fe0av
e607VMl0PQRX3K/3SUFqgV9y65FlagLCJRJ6giY38UY4e9a8CT/YiY6FbG8CA4vnEgY73wez0Gt1
DRLiydOkodmgC/Gqjxe1dG9tBT9Mo2uW1JG2RLn4y7gcN54l5s0+LisuWY4e92+WoIOC8qaQ7xgz
zzhRzGVEOC+RZqvuj6PMiRTFqYKQ7KL72h1ZQRfWWkyqa2R7Bw5Gz8CawSTRYlSlFrixW8vrqW3n
dcFSKkcv6uEF9YunSC4MTP+vbTlC78wiGFfsaoveUd0ogjfcaJZijkyl9T1r/Pgv4tPQ1Gar4XyP
FMcPz36L5KaOIqRVEdup8wwKeCzjOBfR/nSVvpTNa7LuIJg54UNgZmk+ECsLJcbaSlP/GesOvysX
05vgA7UQIxGH4MgJBXdpnA9ivAzKpep1IM42b0xdNSTyUqj4Ai8mJgml+PrwOl8bvv8EYBQVC23v
i8OLUe/08a6TC0j8SSpdw9SDQBJW4usFdfCUO++sbsIPCPe2c9GePR66yZpMKkmbjn1mLGL9vgz5
tYQAYtJ4r5+TaCgLJLciqxDqU9q9Gshzxd9wVWLV+4S5IFFp5l3uWWTYKZHSMvULGeQWe7v3pzyn
bTE78vbto2UiHtohfz/DkBKhvEz6luGZSvmU7U23RgYPvDQcCfcwQxNF6/RMZ9tFjmTrMI7MM4H5
L0RdNcyt6bHB+imF/609lSJM5MfdSVoW8aHkNbt6xNOdXmtia/m81dvNjCil18Eva0j53wKbQotb
nOAepWa9MO6GJCE+BSyV5EeQL/GgPx+WpfWl2H8fMixJV6FcreZ6hKJ/y017PXdKIsjohtG7LxnC
0wnEezxseCt1R4mffjLlvuqWQba1LIhj6neetmL42OimRcomnXq+pEALLV1QYH/450O4m1i1QzTg
u34cvOLrUTLYZfjBa2oKp69VTYmt+CXSsS6wGTeXoNIfDne7zuta/aDHbIsPAt3Dv7ijj/X8HudB
FWMXFAlKERF31X7vgr55X4ctwtTR3B6ll38MZNVioG50pVPRzoLBZdXuMd3glP0DT9MpSeuJfUF/
jQGZT7RwW3n7vqH04/Mvv4DeuOauvVZU3dwhE5GKfi2BPeoMzhg8/cMrdjUZhob5LOnJQVR6Y4Tz
RymXvB+lj+Omk/ksX0ICuO+uLafgeVCySoO4H8nukGejRwH9TWALm0dxZ6R/WvUQ4fo7Zt0+HUGM
JioGOgRe3WDSy7UevypV0PEkMgU/YklGB7h3KjxTSk+Z037mJ81+XNzM1C7jv7RNYVZRKUCuHJaZ
DpK6LR/+nF7ydK+YF5Zbb33jJHdo6aM8vIMXalCbJa/zyC6GZIsHIxx9H5RISriAE6SZTn/4Narp
x1dyfaKfhhfPLCL5Fym0nm9A+bXWOXdpryUY5XPf38Hs0Z653y8q45gJK6+vw9QGUfuKGfR5ouze
nJwKdpgctY5/JVSv63+1gK3AUAP8404OFVsg67MWMg4IQpOxZZLnNWzr5fHZm+zWh2lTKVmSIejN
EeQK0o7MWMTASlNB+YTgEIzS0av1m/LjGq+Qkv3V4lc8moBphenXWMe5OcaizSa8dTSQA7ZabVBO
14HGQdpVxNOY92LrbSsG+gUtioCIqSy7tYg1j7MxGK6JucWcB2f8JJGgRjifLfi2W6tvd58wS7MV
+HPWcySEaH77/4QuKVxulzjFavwecnzBJq4Mg5CFgG4kBXH6nO7xeAy7nXrbhLdGkV8XeLykbSYF
JT9haUwD0Qp6lx1sigOHX69Pt4BtNJBTsHS/acdwD1uAGK5YPryBju4SnwnT0Eo3cEHWZ9oHGmbq
V88/+Pv9vDuIt4jxkgUY22rfth5bFqW8sK/vK94SZnFRRwXmJeLpagRzZOiOeSPuY9tevfOs1Fcr
t6nLBUpI1nJBH0MMjBoPWypiw/hI6A+uB+mOi74WE5ZyuvYKg44VjfYHYVEDp0dvuO6PxZJj8uim
Jmspi73ZNJ4wwQbZR2O9OIkin47nxawD4Sb4IZoCYCO6jwPrIjPB2mJSxf90lopOD4kLTbYDe8cC
dKAp5ulcDyPHp+MrbEXsxuzHSTf6PR4GuoBgvvOiRFbqOlDVwamW6LEE/hRB+HRwI2iTYKj8KZut
ZNmd/txKDFvLZDyusX5+a0PYl3kFRxMmgcynRFjR1j7TQV42VOVxt0RXvYCqZZf0IxHSr1333Zqc
X5vV4rPf2bhLPK3vG8voM//11Fh5sH89udODDx7P/y+261+xRmE5N6HTsY057jvLK9SLnJyY5xsk
VQIyniXmplqsbg+jPRaweJalTaeFY/a5BcdPLe4gmC798iuD8jRBDxXFR8BcBiuPl3feYYKgDglu
97H8FMJV+J3VMTBMWnwcivnogbawZuPKR5BcM1exBkrvbUgJH/f0t557Kl4Ypqq0y2Eu36UQU/la
tyszoY+LCelaLlmAp7Vn8TuDy6bk24LNGdJBEc4CqZIBXKn1xTurZZ89Y0dHeeGpMlt1Qm/7Lq3y
spVmXqxgqA6qEIQPLuy2r5FDgXmKUguLMy4kzCL7MEdYaEJONAuv+fgD22Ox03VOfpaqD33+5HLl
sThXmi6oEnsnILLHzJ4sHOd+s9KS+eTarYyOl62CAoOlh2NGA6FjLDlSTj9yC08GeqT8pFYcO8bX
kIkzdL/ZNMR0/FFTnzZSG0EWUxF0tg2/8H4QdvvzwiRFngWfBriFfIn+t5WwlHtzyZcuquFDI0Gn
VqWRJA6XLANXtbSi70SBBSsLO67lJqj/M90C8glvFM2A2j+RoqV/ELfGV2yM/OI99r1jXBRwWHJD
Kord5rPELvAz7bHAWZVTsXfrE3sz+nuoHVjyQaMxNy4e0q5rdJQ0sCXrStBRFg1Ap2mcbYaaYrEF
ISdq4axx7zd9AyaaM3iVy4RwCg/kNycK4gV4CT3kywkkQxnmG+RGyc8p+YPEBqwxCQRIstQP5TQl
NzIRTDU3EpVTRTh/RT/Qa0NY69RMvg15g2HBcRdiWVxF50NX0flLk9aMSp4jKrdxbi+9+KhroHo9
0/yrcvlQuOdwALN7aoJ6L7tfScke/+UAwMdptU8AFxXcBZpDOL3VKi48KtA81kAJjhocF5pD7nDc
JadsSbOz7my0sekHSVhTT6hTtH5CG6Lk+kVPMqx7KfJUBY7McX00XVwFOMswk9D9KvfRtCDzplf6
fjhyMZXZDauHRAK6X5YG9Ge0slGCoHl4YWQteYYJAiI0c62MUpbU29oGBWNP+cbkh4DDged5Gw06
61M1AXa77MLgV/74j3rrK9cAuoGN8INMPt/xhRuWx0mtZwcW8FKWKxBcQJ78jFTX8kKtGtYc0Sow
1WGpdKGm/LJ3i7NjXEY5WhUa4CpwdgZhosVAppP5cGjqUz18HO+tJ/QqfZWYucbliO19QOM5sV0S
wRtEgDdRU/DdT0ttMY1uPJgipfF0zR6IbqTH6UzGaca27oEOcIxIona7F7KmpzjnGrTAEN2li3o/
LvidQbnkKZ61L1TlVMkMLD3dslHzde9YfV5Ah/6a9d3R80TK5f2ZjAIBMUfAv+r/WHLBrsCQCnSo
Zj8yd/HGIEcfD8c9CWcI+sFkVGQxt+PkiCJvdtQ/qmw9Ln/ov5t7TBtlxI/fPXiNGQXA9h23BRGH
gUcLFLGKE0VHpzrSIDoAhvTwCv8j1AbEFARTQpJ7OsO+p4KhqvyMkeh4fk+9c+8plWp5QMtkCDvB
CG6nGS+F1QrMMYTTQP4VjLIoA6rMNg9hboGKuIXxIlX21KHRwwxiNZwOOh7ww9H1P0nDNvP2f2Ch
AZOqHcA41kOoIPX++Wl0wvVH4/oZ9y9tqiEq6xbAZcFWU3JItnKp2cGqcEcp6ZZi1GmjrvvBvq6B
+zSk8zXR1ctq/DDTb62GwL/eXPpigHO6Z/OQgVs1imZiv8m/CzluBMe7X1bo2UQvI9/f28Lkr4/n
jqgZgNYF8Xy0gqTR4y4k9RRM1yD/Do2EHMapIWiDfvfhMWJGW+jentd5cYzDCVswRms6+LZxXNH4
vgElW9IAQu5N58xuK5+f5WDhtKHxL2HCfyM/3KvJlAWE2dt6CdX+JYxJh+id0OV+57iWbgNVZ42S
dMU+Qn8Ox7Q8l2NcLBhwsMdI7ir2h34wgBtsenb1BbzR6rGl7YDfOTv7PaQkWutOm42pgm9X3H1C
4Sk0+e1gWEfbaub2R44wtu0ATvj2DJIxs1BSTAv9AmG8et2Z+uKdUtyoLx70m8tH/aMUfuIdSJQB
E7LC6ycU9H6x5WWDbMjGbWHDK8D+PS1qkV6n/L6AUX5cAv9Tl+TzxP3SP2kXENiKwhVoRTHU56e+
5JCVtOHDbZKU1a+CPzqIk3XtVQ1Y8ATYfh+aJHlp2+av+/8tzWlIJB0Ar/Z/fNLZfCvAKERog2Dz
gCD3qYLztFs87zFXD5V7SHJ1wlLDuEgib4UNiqX/XG79SeVjwfIHh7scjKGYAwUNjOB1dXb2gHWL
J5X4gFT6CUsAn37AqE3aARQTbln/j61VqkB86zAS1nAnEFBqcw+3qUGxVNdo/T7UXXwukUOeYhYB
dF4taq55bV3BnbphoC7QRG4ghYfMBaAB37KH58IbN5UktL874OYiodW6lESE+NRLC7r7PjDNJqGr
JgnIEQ7qcGMeXgkVEv28tGqv9HZ7ITjaGqMxz1RCSmYj3Fv9lI+Ju04muf3KPA3Z5AZo6I96qKhg
QeyU5krxWH+etOq3scshbXvqq7CHDXh11e9hOgQL42tM/5QNiff55TPFTnX5UhbINSSyaK5qJthw
HOw144xiDLCh+I6Gb1B3fCUF6gyQCqTLvXWKazvf8s3FIAjgcgLYMmdgkp4pdCmo8nzFetLaL4jx
UOza6zmoUAW3a3d9sw7ej9WwSlexoqiwotcaQ/Md6RL80Gr2epuN4qnhhTNgzM7oNA5n/zR6cz+u
5gQeB3nSsjt45A7iEabJ4C8XLbpHqFphbLW+Bw/vG1e69bByroU9QOFd63Tlm45DG/putwEE825S
ka66hjErsKLALWq0L5wETkOZGfTjRSa26VogO1QHGTZj9D1onxUwAnRGT2XBSD8c4Knf4iM1GiCO
L8RvvQH7OhoR/0JFaPYIHu0YHq+PwxSYnZWr/L1GJ4pQXGNLgXFBaQSr2xDjlOoFxfkbniA5CDnA
A5N2kccRVlfwUTfpkQ3uijbKqR/oxJtQzTwHk514espU+4OhxhgqvBl9TCQ9DvwiCQDwArY10Hzx
o3f93dmKEbchVMlSEjQ07u0TxjRVL2LqZQ/mAt6aGojcPKTtri92/3TaXVmp3m/4GtoISHMlRTJt
G2fDaTFi6Z+Dmbs50AG93dwwXliBhjIC9RV83y94FGgI/4Ldd/BAWVJvkwcZxL7Sf8nba++DtldC
Xa/hE0M6SSToV1NB6YiCOY2cdvZ7LdK6eYfqcnaDctbXXAgUJbo2G37sqKmglhzeHMTjPs2ydFHC
cttWrd9Sxx92HZw4lOsjmC+c7O0HWCx2T9ehka2qoIQJKbN2kn2pKaAj7Uj8nJl5udieibpu3i11
b80XIQEgWM+SDm83TQ+hs5XugtsBBCdIcZEF74uyOkpGMtglNNmTw2wQ/i1SefOw0zymMysiQnd4
IYIP1vTeGhPEvXZK5vk63OInP1w9rw8TF48Pr7xPtUJths0CTwnqTNUff8Ef6vzOvnq/xp7iL045
MgJ4eCDVog4ghiV23NaN3g/R3ybdXeJbr3HbYqNEMc++JCTsVmE/jlKbppWX7qHOpOpHOitQYWL7
WXJSfH37Ilw1f8JOG8j5EaTggMHjncy7rZsrmqUZGlW+LrE2P7CdBq7o6uCaUxzJuKbhzsZ7CaI1
SgTJ9NB7yQLl9VW7Gg6pANvONARjIkphA9GEYxKau3PqP7qQMDXplD8zaYytqNSwcuNAK3Ux05AF
JCHTSkLXoFsfio7RB62259RU1e56qW7xz89o4njC3dGxVWHiaC1ZGqSTPwUxwG/vba0o8vYkbQYJ
lxWPLOmZqWPha+I/dMh03YHTj8Ar5HgDG5oGVHMUOM1IgaWP1Yxf86cIPhPralyyT6ihnthPhW9R
vPtgnGFslqFq9gJzy+irC+l2cEl4z/lMu5ypq+yC1XgdROSje1ygW25qG+BYGf7eH4pJ1HE5KuK3
90y784EYRo91ei0PUouAQqwf/vdX6NWz+8phZXuxMxntmLrykwLkyuHzb4t6QPhaFjPo2huTTc4X
iUZsK7ZPPgia37RJIn4QExeGwN+thFs8cHQRaLW5gnIPaOPEW/+Zcr8b85k3dKrRqeEt2k0dTljC
XSLTtiyBEY9wM+0/A3Otd38oGCzx54Sk/oYxE2VmF+3ogEbSm93htOy9xZ+bvEYdnyJarNl45EnO
EI83W7vged+rvgWbG/EMKti1l/IsNnA6yJLGW9nGC1sfavVq9aH6Xy5cebIRkC+B11D7M97hzBfZ
SqFsiVssmd+S/vaZ1s/4T/s/1SecC1BUedPbDhNO55vWo7CBjiYC00N+hg9HVscubEJ0VyT7sV6p
SCUne3s+7Kc4RBB/vNejJiiAzekfwXKp96QKZ939DmoSuXlb3btxUeaI08EzBtPp9EkwNGtrQbcv
IiGrf3knxKktvvLtxS7+DqQKB31cyt2I9o7X07POk3rFMcS1jTh4yfcKavWscedfNJU29UXja+tj
3Wxsug1wzI1vEwxAyPYDGOMRwM66By03I26uGQe+lb3EEnAqBlSR7S6FEH13KMnHRnuBSJk7OhyX
15kIVZS6tRXqjtZ035f6uGSkTbbN3qtuC0Npg20S9JAMHfGtp6BpBfdIrWz9E3Hbbrsj9W/nu2ql
y9HIDnN1xW64LAjRlnti06XAbq6dBdT/f0L3BxA3VD/dh1D47OKB9WnJcsv0dUCz2Ftdl3RHpK5p
EbooUpd/SIVwBZNlev3awRXWtuLaeS3cTzecSXVWCM4tPI717zK0Q6446c60oiOj16Z5gLb9SOak
M3zcMEXwr+tB5brm2S88zrhiINLNGJbEOopZXs++RvuHdBzkf0gfDxzlkMPJ3dlu2UlL/WXy/hz4
vWz9u0Tj8Pg//gkCn5aodOKCTqDoFhaLMC+X2rxGchtaozGb4Db+peQM30HgZQ2wxpJKmCAH9O5K
uUtjvugunrIJgrBg6z311Y4TtdrijrRZ7mCCrKfq3/uPDBUn+vvxetjK9PCaMiJEgDRppGWAF/po
yun7DdFAeGyxl3znnAr4ZpFfLmZyk6VZ3kxj7GFfo+A459l5pcKz9KMn1eU45kKTkeK7kKIwHcWx
Lca/NaPVP+ENkPF6rXqSHgad9HB7gHthgP3RcGVh7hVLdt6cPBCpPb54WWLqXt7A3PaX5l8Fpnkg
Lz7XDf48vE0xe7iP9s63T36rE6UPVBvfWL1UPUQgdhslMZpzhFTGkHYQsodklvpurRB3yzp4OW0z
JPf7P9MYKUBrV26V2nNLExioz1v9ggzYWWilWPLG4ZHaaLoO5hx+4Gq89LF+S17LLATXi7sh+KNE
irE8pKA5jBBDlEHCO0CPViDf9eBLWY6x3NKI2/OctjTH6aL8b6Q/ybwPTcgRRKrxP1a0p3+UrWGD
QaGDBItZLFyDvwsU/v/0niTMGwyS7cZnGvdyevLWeAbpY7EHlWBgtfyeneg9zmMfK2BC80xttXT6
JnvdyidtXYOZMHvgyxWjlTqRSyMgGApwfzZ8PoiRtSnUEhuEYthOAJTMZjo2s66E+cpSFbTIy+Vp
49Vfq89S+qRISrjXNR+lev8LeKJUhnB5mvQCjHFsWRCbsQnfo6otVUpocxedYivfAQPodzVcRv/A
a8qDTvX1HY8KqIpniPnLbSvk/uXmT7xz1Vy47ATXf7xF/1WhaUChXhUtbg8x+TS/73FRLaUWdNXo
uv/oZWgwdMznz3osVOj2ALfi6SUZy+ekuz1mbG4DvtDrLUfqcoGLQdcnUb3bU1hCPMX/fYQwsTaT
TLee5Br7d49Ev1Pq/q8Mf1nABDmFL6ytLm2Van+VEqk/EdJXwosCftUKS+Vm2fM/E3MznX1fYjPg
j4BegWhtpyrQ59d1fS1Gv06KdvQSgcEeoX3oP0dsuwyRb73wqIUY47ik8Bj4xFHCctUGs7CR2ua8
qa3lsFKKuJsgZFbRKAB8/3roIWdCrNjq2ZdJrGsWobnAmDvd5ThYABubbkWV0BRSkcM8pIsWez8k
67Qpn0jXXVI9zgOhpXNGgAGpkfTXZZvimStCLIyw+HjUEheIAeWesLxWJVGbCzrsNfHWDR2dKqv6
/TvNmvPvwvGqL3iKUSRtbD8G8x1F/V53CDqmaKExXFVPsE7M73QQwFxYahP6XoRfy8anZpA7KP/L
syoOWWra/znXlWis2Q+4TU1YPasr2uHt/KpqJirPv4GpJNzlMJc6peFKRLlXOPr66K00U3zZRXSZ
/SrxX+40G84R9GfJSy2Ce/jFLeGODjTxc24w3IZMDZKHMY2E8mOcDaLCLbGnO7VQuhGtHnNRef48
Nz6wMNtWJF9NPVWJwnrp4ItUskVMhIWz9vcr3uP8wkiHbNjhM87JoOndaKftwBvJWFAoPbMTBYcF
F1G3cxoZUe988O/kf9KrwtoZyDkS9Vh4ZFCfhemlD4ggYVq4o5+ckAnDJSjf3a0Oc9m8ukpkHd5p
phqter1Ck5zQ8zQ1DPfUSyE0RTCcHcLBwJKK1r92Q79C1VHXyQmAzSaHyLPsegmsF4iFyh1OzlYl
/dz2WY/C4tYgU+sehWe4yP/3dMAAOfEesZXrJFQAlntpPQQ761o4tF7E80QZPWJvjxDuxs8gqGSb
yyDOEiYKW8N3xfbcSVyoGwQN4xgK8LggXCYHL2HnO+QU9JugD9vWV2FH9rV+kVxOQ3lFcTF40WZ8
W+BLPoIk9AjOu/JlSV3j4F9pf2zpu6nfGWdJvqmRBTLR2hm8tjb85LsCSAB3U1v6xLf5T8Py/MTI
uAXobGBHQGR+juRYgG+C6FhkXduW6nRWnitH7FtaQLFtlP+HVwV5f7dy3qu1u/1qMF0fzSPGi9X/
VGTvRQX8RPpRaA7FYxhmgAyokIwU9/wTi3be+jZSGzf/nT8ImpN+NymtALEyu1poqJkeJLu5JSMb
WJqpUTBmc4qIEat343AeyaajNYVrhB4ZoWyysmX6GvcOzRkqY6Frrr5jRBd0pB19dAD3zi1g7ahg
Ul8nuZ7kfWFp/DG8XOVO+w5YRhMi5BrqC9rw5NC00CGT9h6GlmWs0ffudomkh91BvMklccChOJiy
HC5yDdn6Qd3XxMj0nFCgsPgOZOV5ox7I27gw54liNqIK5Rn9vugMilnzrflTasxrBGe8UZleHh28
joFmKbnprVkOXD9AoYfkvYgDblxTZBewUjvnHm7kPXuwqELWBfBl/UDc958RY1xy4v18Z69pd+Pz
nAdXgZyFL3eTi04/ogpi+jw8ZyjBjWbQwGJRwALlb17gA332GDoOrHtQHH+JsNkUb2z+GHETDI5b
v7RhSJaBDoMsL1Ok47ylHPlBUVyHFJTjvtA/xLLqQUvkGewYroAOTiO6oPQlivkG+KWvJhj2Ms0z
81WT+GrBLfnd8Uy8qKHWxHn3M5EFgWx2edgyxz5f7kHc38/dXtEM0Sk0fkY9Pjlxo99gIrLW//MD
+EPazF4vnIA2hthp9mlGes674x1bLxBMv9EYKUAY/wph+iOC5dq8+4Lak8JKcl6N86PKPleWze/n
GYW92cQtYmsTj/7j3qPYuZJ0A27kESOavYcabA7da8dRJ+gl8hLz1yO5Fdtqjb0GttrZgupXlbOf
VB2dVtwDnmP45PlJfBSUVjNtPKUnhtpahpfdhCbm9UzoqpkT+OvZlXrHEltzoygPKdAeesjE06f4
s6rxEw7E+WEqKKFZxjquz//rHHhJygeJILUT0CTNVayZyVobpRBV+WlHZznn4vQuAEVit70OjGJ3
0/XPDR58TNY6zJGJblr0JDq6D90VDhJhTL3R+/BWc7eKgkBrIRTo6T7lI2bmI27cgMy/iSBVsF6N
2IaPL8FoHjggxlwt7Tq0+4XkcKk8PdHQjLoFyLzRiEtxrsG7+M9bQqI9vlS7UAOzmNZIXRrikMvk
wZY4IomwQ/9mf2y4xo18gfR4/xr8RqDKQ1sDjjKhoweACvTkGGb9i1AtxQC0XFwrQYjgKqfqfZ/s
9uTTuW84FeZXaZQr/U5hPByvFSqYv8+TZi1KUzStUplQBAL4pAVHwotsI6G9FJmGnh8X9WFeZoVa
PT71KuGfxDHce0G0jzgARJ/REYghzevTMlmGEjkXESkF8Eb+Ixll6AXUteis57KeH5VXgfturvWq
njzTZG6Oglov2BrhPde1J1VRbbHNyf3LSbIYfsXMKKCjIWWBKi2TNl+F//rp9Me5uAbRypW/mIte
r3dTJriLfQzeIdDDBP0mfuG9Cr36LpdddcBRG/Wi8/O6KmF9C5s3xcAYqD6ktf3V2+jLLFhB0AcS
Kk+6OgM2DyfGthEJCz5zesxTukC1HGrHHSz4OuwYfblmu6fZUBxkXPgZNcjmpJ+PyQWHT6O0LMHr
jmJByOrDDIY4V6kaG9xPqllMU/+n08unWWGUniNJSMph5CPDsKPwFu45atVIbBADQ5QDi504O2dN
aGclamZ/VLrSP9ESpjUYiC9oDhMpAW3vhf1l8ooyCOJ5tBV3OtSKk2d6IPvHoAU88pDK48A6ECoP
AHvi/oXoxyx0c3R3zgrFI4nLeKPS/kw8Q/KDtSbSLYCW1BKQslv7WbQUZxGSivrhvMkhxlvjIUo2
NymfUO4v9Tm2LmPTiHl0vGb2NcI46798T9MUF8Qt71CdIVSpG6fZ9Q/2uAaOFURFlfCaRs98Kw5s
XFtyHEj+Up00h1MOkmyA/+WTYaM0romJCfuWz4IR2uqx1Ru87mLpmsu+DeffW817NnkRLi1En2US
1UGIgomfIYtMiGdDtGrdhW9B4WK1J2iWFaVrJdo74++4E/IhUoT5wBZyF/+12fIh+cCqj1uuT+Jg
HsQO2ahkkCA6dHMd8ZNzcTNhZtDxQgHs816Rp72ejVTtVqkoTG7jVvi0GNiQg/ouHubjgxI7u9el
ywUgSKyqRI05MOVROc+E2eF+UwUsyITjufcVAQtA4aqnurzpeZKKuasfcZM3l/p2kZxfohmS1Vqk
opfXXFGQsdg0z8x/6G3r4lS7xYA1f2blLh7ZcYEBy/m7ST4BVMnXvxijWMnrkZ/WPGIWZw2Q32P7
6ukgSJEh1n3RWE2NCxGNFSVMWEV9rJTY+2jSSH7pobFvWKbzh9//DM1gi07VOFPj19YTSi66nNNm
kD5skA1jupKyteOBpt7RcaPzkifeh+1TJolz7yJM1S2F3OF4FXEqUn91ZXAw+2E6KvlJem97CX7l
RT2Km1TByrvW3ZHq9Y7yWgbwLvtfEeS20LcFN1Pyy7fsN2v2iwVxz+ugDtE/TES4NKDDvJBX+kgj
dYW/kzNT3d94PFCG8xKG4JyFICvDhe6XCGu7SKxIuHB6ekLNa31k71KE4n8I89D6sPw2nVE7DiZz
BfeN1E5VA4axuTHmWAAbTvolRoiET1+p7OaiKRsqV3jEM94HI+pZ4s4uxtTRRCA2tHEWcXxLwBib
OfxN4Bh0KMzIXV3qOdLC8BxaYgVKDK72zQiaF0pcwtviVO1M+YMTzmi61TvL/98z9mL88yat78UB
XI6OHdkMBsPvx9xkmCtjZw9b22sKNj1bMRBmOThazOcWprAGbDjsfbW58pOkcp+L4CvJia68/ZvH
gnMv/lu5lBXLgew/dlk0p/HFZe+uAvmIXP4hOC5FbFId6Tvv7o4lt2aSYG5ljuXdjTuqHa5CYQOD
wDYwP0GcQ6dt8cpGw4HMKDJQ2lByyH4nmF2DHyjKLb0wpggWOoJXECYtOXTMnDMNr1QD9QMzNFcZ
Siry8N1tkExRvBlQqmRdFurWKP79HoAZl1W5vLXQzpR8e7HtEmmDyrFFzqLtpzDxSiJOBsE4xL3H
/JqoVo04yIM3ONc6bvUDSi/BDaQOfGwbQlHa5ghIReva4xF61Qek3u+E8e6A01hjXbY78AeThiJS
weoefBXgZ5CPE+se8yPGTbcu5ybI6be3iVqNWKO6bA+Z089UWPem0sJyk/biaJpNgxo65tq1kfMp
0yhLR3e4iG8U306QOzem2ySzNhzCPfZduIXGSV6OJuBloT8eXLrDjCjnjmAdG7cOry5ouL2W0Im8
dW1gUOA1Ai2Q6aTGhtnL1s5QPfJbE4qOOq5hg8kiKqPSE46aD12c1fjjdKD+GKMFZOCua7Nsot+S
C4JSUgnWuDXDMJAGFNqGsSKxQspAGOse9839unqq7SgvhxbGj/q0581nAiU3KvH2CtKDPQKLmDQU
0R74wIeW9LU6qb4bkyUtBKlp6s4j8oQGe+DWokRWz8CpvYplaLyOh4KPFy3wjAtl55YL3p9wVPue
DNNVoFmEy2Ac09slZ42ExS+lxCbW5NgpRF5oDn27ESCL+y/OpGgToXrYuPV2HXoSYB2nx/xOBFR6
RTBOsvJ8T9XqMC3AK9qnR7lIo/jH2V5ep8nKci6T5EKgs/iuGBO+ay3/nxz7bJYzZn9Yn3xIDPrH
BQzaeEbZ9gcm9isgKmjFlEgQWAZde3RYmabdJuOWhsSYzXf13Lu9peQJnBgyrGwp+d5tQkGzZiyJ
KT75xndC3pH3Da8pf9psqVUbJa/DJLBxEWJHK/D1C18ZV9qd6NBFlx0EE4USBxV4HZkAKSZPX4uo
UfjUgf9QCtiXH7yEt+5GQ9bJqKWdINsHDoiZ6TDek3uL4EOV+0qXwAi1/G+cQ+8BvsefWbx7DqJ5
E2ExuefIF4AjZXrAWkpL1gqs2mwCe9CY1IZVwxcCa1sfDnPzJ/asr4Sk61PimpsfPciF8ZHGMYot
5zpyIym0EHYyrrLPLsGh5AMPZi7D2u6YJxrXdoDWlFDizqJP9lQ+Eh89GGaG2mR/Oa4aavBrhCsz
ZF4m28S7noq/O1m7nLqELPN5uH1GsuJpUUzzuob32Dk/xciwOj+jPDUTrbRlRuJpbRbaqcTovBUe
9K1VZI1FFVr4IwQo6VVjtkJp2akxM/+aMQf+8iYYwuvjdKYjAjTaynm0uuodqJexGETyiptwVCaA
pdUgV06tNiNn7ebn+ZFzRhyCiwbQ3izZbn6cOUuPIhskBYm+zurX4lMoq1Cc0qsLFvaAWYKdxAoL
/SBnrrShuLsB3E8nod2bGCbGMtKh9xu7s6JNLsB8xqi4mp5BgQTl6X9UQJ4okeGSAvpRd3iRs5L5
kLDNiy1F1sshrlb7TqcC4CImk5IuELOp/Wu7fxR5MOZPNeF/glSmxfFU73+v87nIfTEVbg5b9NuG
p3tHs6Iz8ZDuSwFm07a6nySMytmbpjVOLlN+3vCwP5Zx4oG6C1kFrOKu1CraocY7+g/1c2Kfreut
KdOMMczP2lXbNL/oSPvjNWWhCTbtdKid2kYbZFzAO0FKWZ4RdRTnY+3RF5b6GySdU1a4C4iYcI/+
mj0bjVek1baDiNPjlcOQxlYC0py1QBQygOMhWxyIiOmYgxdD0As1yB1HRRDaIsspkxz8aQa9Tr62
3bxecAdwOb+IO/CGUJ9GXgGwg3+23hHVUiy2kV+FrlFRDBxI8CLPGEdEjQ5GUJolLGfx0+/j0CsS
HsQ5haL7hL37GYBoRcVpBb0fQjazpmKnrGeN9TpRf2eAvdgmVV4DBolf0h1Jmsu7j2xNLd7hpu2n
GyPKn8YWClv4NOOlfOyPfworLHovdZMa/XqX79E+xyF+ZbmJWvsu2EOm9BTbEK0c5CXX1z261RSG
QZ4id86LpW+lzQ29tltUPhyAsp6Mhal1YceFfAnpBhoaqqg9qp/2Azz7nW3ECeXHyLDkVBrWxkE4
aQ6VqHVtSyzjbes9UGXFrnHJEWtb2U/9DiXJUwyn3M4aiy1qRQbZbq4dLX/mfBzBxBMG0ZuNCE1h
jzzfc23FpQUO9xllLEXcnsJycskw/4k5xpvoMm9o/y25hyce/tgtIqT90koxVY5PrcSjPZtYwbs5
g75VIfWhFXQH2JSB3lbPb8jtRN5HnqMyLIDnpZqocQO3FEDac++hVNdsb5CbVWYuXxlOJ1VRQxpE
lYKlf/kkfZCdFFTqJT9MhGWHcgjg+TjYOIedQimzEe2hlsaoW360BSXotHjEnubmxvrPL4KE/sl3
O3qzsG5iZzQ+GoHBF8RM3R06Pr896gJFYJyY80KQtP3A1x1O29a0Am13q2Ykrbl/chNHd3YTc58Z
B5I8EEKiFoxpjlwmrHVlTudiqJUlB3e0SM5HFeglE9ZxynDp2hT/gg77BeJ7OPkA3/TknfeEZGwD
EQBidJtklSo2RXd65o2GoAOuF3pN7Dxu0Pp5vSImOO6sdMYlgDDVBJf6BsY5hqWiVlxSr0I30z1u
3GeR0Zpx+Umix+caEA0bwmxLHDCHZoR3gdqIp6FzgQe2LSXGujeJj4RlSb1cxqzOeJ/ZbBhQ+E/S
Mq5UawPajD10hoHa8N6+80QV7b1YKFR1dG1G7/dB9ysl1bY2j+jNNaTGCtIrZaMevdjZUodVHuHb
3yxsIr6u1b/g8DoMvxJKPzKE3xwVWuH8xEF4yrUc9p5TS8ENXOqEq0G4dEkGA/GrD2nRdfmrHCs0
hsuqjn3k3ybqSFUG4xlFZGdL850+uRUBHbvdkG2L1vtVffAKZISJutnS2CNFKXnJ2DREfCQRtWyn
MaC1q9T65xvxK8r0E4Hi3+npwKLjkqqn2TpN6Q6BXv3tQyw+do0iyUFfI1v61wy07ebwjzMk/Zz5
vZeb37B8OtrpPH5znQ8wHvrrr3zWgiec/x2PFPVZsqJomH4MiVqKINTQd8Cz2eowTjSk8WqQFrZU
hsNzUshKyjkMg4sP1Fav5l17z1uLw7lOVN5GTnRCnTSwBE4yvWZtXBANdOL5tGioORmDfJsYTbeT
xglTPW/cFxJRl7Q63AvtK+6ceC5Ari07rJOnFgWUabu+kI2wtvo9YK9cdKdOfQdl07RajyIwg9TA
PeZ2gbvwGuCjv2ALiLd+l4pdncRYaWTxtGHgYKmDOdK/Q2/2EYhe1UxV0AqOX0bgH5VyPoatjzLh
bPZ/kTPcJQqdj8GmZi+75YDciJ9C0ywSLW1mCEX8oTnuet/f/0rN9ZaiOVLR7GPY0Y9poWI29uuV
MNE7Ml7ai8o6WMWea7j6fY8c5AZp5a/jVHi7HRqGiv//g9DJTPlqkDraDhy/JKLIMZN6B6JG+ofs
xK5ggxXtrfBZjq/HIUArLA/uc17vvB2nZGB/Ta0F6t/0s6l3r+2EEs3Jb36yjzN08yK9DlesELPG
uMiF6Tr2v4yjhWzcF5rnZ2h/cvXWAyq7PCmn4yNZhPpMlIvQ56DDr/NcBIsPJFzAI/zLUNifkqJb
KZ/ervz4QQk1dmiBZ2dM4tWzCq4hSgCvMj4jVU4uJ1nXftwnO0tWjl6cKz97s9L/A4fkpGXWO+OU
4ofjxwqB++3w1F/B3Zsuijk3nVl3nlrPT2t3wFSiNgr42btSIXLmHpO2jM05qyhMIpuu34sG2g/3
DqaTXXrmi0iAfkZgEEjYjBQcV7dUQEm4kMJxxOOFtZ3T2suyjYgH0Y15JCcLiqvMp+7EXc1ZL0M3
wmpPpnoQ/vDQTukm1L1TC0CBECMmgVUvfBq5xOCNojCQTVWlnV6x0FxjZ6hdLcrX0266UuZ9DLYq
A+rGhTWKNm35KsxyY/XvXPnK0QyW4QvoWu3UtISdqXJe+PDnbESG/Uzk8B8ylvgJwZhrot2YVD34
AtTQU5ajrajZ35O4cNrKraLX3KS5F1cKiCDUazOGIVUqu9JGdxwujA5rPtxH6XuYkjC+NXQK6Z1m
yXSA+W9eRczywSYJMOAImFmRoeNukZkW6cvInn2vhUqQgORbLt7VBvqC58yujLDmx0nj4aPYTWQC
eqaR+a+5XceC2IJciGeoSdi2C17IB104uBvbnZv7rZVzbe5Wi7L5Wmy6E0PC+e/zLHnNSWghmotp
IAeJOxFB1WCVTPGCwuletD8J3f2mCdPm3eGAGaI0Q7RurmC3e6D0ZZ+xfRHmc77IgU19tPsEJAEI
JfcOkJolZD9iubIJO3JMZO9JFIuGSUUpTv90jQPcsb3kkKGWsG2YBILqsjm9zSd1YjC+IEi3u7cV
/pDfbZqfaPmDD5eHP/uPn6EDuoB1h06dztB7a5Fph5c0kVNKc4ZoPIH1N+3F6sWHFe89y3tLGJym
5IWbOIl/kcTB/kWob6kwWWr/aJgMVXUOS6EsIXRvkX5ixTnqCdYlAqgqg29MY0a4kaNzrJp3ufqG
sGpZ97iJSIBZrpAwkj6XPN5NVUX+HDt4536Ei0vvDtSGdnF4Mt54HaRD8BxliMKB4db7GvA2ooBD
zAYPc0j4kgVvPd9xvl+xD5hwm7a8BayfG9D39MK/3HKpnm6+D3qTHaQ9EdP6P05WJL+7QKum5dil
3vl14zmved3y6ZiNSaRI/hLJmCLxT9fGSD2N1i7i3avQqgaN2AzWDJ8oO/qIIPHBgoH40frhA1JX
H+z2/QQqS6ZvGLh/MDvCEhmeIPX59dn4D+TEslU2pQ5CyBNYA63LEw6VR2vxK4sQJ3lGGeEyQbpo
piVlwDSG0eYdeG+OgQ6Bbomk8yOoTf6TEGrIUcIGr4qp1nOXOhjdkc3+GezJ2HzeeECPXIlFdkO4
zrgUk9o6erjvTqjm8RUpAvAAdOHebd3hAla3NgCulfmnVH20x5ZGXoZRObuhXlxKK48nLB/UDnJ/
WGiZ14w1PzXE1OIqWvVzRi4kMoXCKnKyVcQhP1HhSgZoVwd9zpBp9qVR+Or6HCwBtHWPZzXelVNY
77BKFfTe10erNbJfKAeFxBYNANPYnZxfs3gBnQ35LdlA4zBaNd6Yg4FqT2lRgzM+lqdF/fo4La66
SBy6qnRr1hSuGaTNt37+evu3PhJ9RmIv6FiIm5mJP5PHuXkB5ToSv0kzMkV1dEKdOH5Bl6zYplTq
Xwo4H1VxuUaC5rtTv0XFqjf0g7PkF9EpTMLkQffpeYDV1dTruRBQOClXOuW3avsJMXx82Zgs6uVz
RadgIRbRtRd4CHU8h6K1Bi2BekGYb5SUVFZvkIrk0WgTIOTciwsQKXOpuDzNB7BusMUQo6lngCFC
cxM0WB+T3XKLxZ0EcDDFEGC+Rn2mZWGqoGzX7q3xmu4dlLaTDl2FcLPs5bO/PvML97QjBjJx4YwS
a2Slo471JJ83r8JA0kI2WGHdsTGBF2xqXX+hhBWJzvq5qYEjPJWJyYECFUOypk/urWAYMhlnOTUt
9b6wmOTW2Pv75dsKXKzFuhUZ+UunOaPRl8ZArNcdhrBcgE8syyKf7shaMI0QEqQ9US9jhEFvZwuM
FCvfl4FoB1KHrVEN1rp5aPn/1gF+X9KcWrCYDJydHJ7uwC9U9HgggEqmD5B9qjVBIkRmulAtjMIp
F8arTEDKLgNQULKYbbS2EfAa98e9wQFGGn+d01e4zt6Pm8Uo9yYkZ0qHD0lSydDE26j+9ioT8z/u
qYfLd6rxO24zqrftT4E/wZZrb8haJsfSsWgm8kokcbvS3Exi+tons5/4VoR+essN18vitmfXKIRZ
iUpbi2nqSvk8GP0vuNK8pt6MBtykT0/DZ4ZzdMFramS3xNnVJJ+ZMXHQ1Wo8V6AHmla1T7nWZ/wx
jart0hJtpGs2VsPw4AVPnYNo8yDm2n/gz1K57RAlLIru0LO6V0LmH34nTn4SAQTEunSUNHk94tDH
P2kCgwWdICNxLGa/ej57jK1ngo0i3a9u28v+dOCIWEPKPr33/tgSqVOrJkruRasbpGQx5OAVt+zZ
sUhERD+ep9bGGGmnOYvuh9mUDr/fy7odAoFXHT7pgJyebEpcCLyntof0T8+0Gooa16OtnPhlzV+r
ou5zZ/uPbCcerWLIpweOo70OrrIeWD7VRUWAnVjnHCCmhVehBfEDMEECd9ZJPIrQegiLpPjqAB7Q
6Ck560eCsGY8OigGwtROAtEnM9pbWdO1Jybd6fBqhAOhraPNPfiZbSboCwpqM5DWyNCosyzGYVkY
nvup1V64Tj4yOhtLQp5a1baLHBKW482pfkst0E58PiPG6dJt6jNiDPPHTQv40gkF2RU4pU60F2It
v/t15sJFrtptfM7zU0nU3FjwOR1z5K3GrqF7mZcSzfIJqBYC6zCjn7L0jYVi7iifGrzbQoVubEg4
ZvBgq9WbFn5pqTdFJ/m9uDpLP98ANOFpDx8Nlxu9i/WBATH3G5UO3uKc5N0uHpCJIHsRWrJU01da
UxMDoSNUvHEib7rn8X/u9uZ+BgKDTZMYuqCVLZkdGd/FZX37NG8sq/GtluxZ0sWydyq9Eo72do4k
/dGlB8PMyjxoKPmNPms3QI3Ospc5H2yzeSD7y94YqQyRUoQ/3/AMZF2ekaG+lYhaZrK4nNQ9qCWD
AC5w0Ji0kowdrTiLY9OUtMynyWafQkII0+ULqaGDNmRKXvp2jM279i1gT8247qEaRObLNP3WiCTt
EmcawZP1x3CTed4bIToqUI7LF7G4ZfUfKnr7FSyt+v82WbhCdWRRM3UcpIcWDym5Di61E8XkK0+C
wgCgbU0l3zX+Q8dLdB0reZjuBj5jD9eK/pP7ImV1HEc3NfgGVvWR6+W1kjstZ9FxtySHTVlLBLNM
fjXU74yvvORwEpiyKM7Cmen8SvVCWkmBV2TOtl3UXzLdhqM3WYLkLu4UGMNKocvJ7SFyd++EgGbH
MHokU0yhUnbj+KmiM0Wa0WCs/Qx4p7tvn36aKTA8S/XiXqPg11k3UnYiX90SO+DMDKQskLTh5WZd
PaZ+KDkX3diX17RWgJ6zRdaAT9185+DmzwKTpp4QPP5ypxrhZNUJiEjxVdzZROAXX2UK+8p3KWTn
QpnBjIIvyaej3nMSP1lbBwMgxNCQCoDui12JJ1uoR7GVSe9T7G95NJ3nUnpDYAzsDhZVMuz1etXG
hqmZ15Q/3QsBEUoR00z1r1yt730AEFGkUfs7liHNjgYSCNsqm4fSFW+2ta0lxM0pQkpdTOhLp97W
bVrDayh1uYzgETEC8mLz55uToUhTmatmZmZxllvPCtr66kLnkZUrMsgcOM911fSBaf0jh46bcu3J
lFBMyD5ozio6EJiafV6+elNxFB7b/bDGafJaTyNBmUfPtcM9HUItPwe9Y9hMW0UAhlFwg/5GpguH
9G14qU+SsOn1PGDXX7DRE8OMHsVhCRPm39BTGNyZPLS4yxdByYGGF00BZTpqJAMJWiSeoM69zUEB
XaFSumiCkVomlJdzBSgy/7eHIDPpdcVUtYkljhTAQES20ncjA7y3YbGmqqNoTwYwwAjNOoSGb+/A
Ni+eLtJmoA95gUVW1nW3yoHwIYsDv3sOQRXFSiiAXLLTmqGUe4sabJMYbjFykpmFO2oyUvLKxoWh
BDciHWjwt4m7qTw02H5c46oY5yb8bUP83nwdKqOqw400V6X+uzUeB8d0ShSp5l2c2Fkfy4LdU9tD
JCmXHZCnFgBed+RImdF65CKKwS3WKHEeWzYhJLb/hqTyY7VzmIHdXtzkcz1b29pmarEqrBLHTu/N
JsOXP/uo35w77YH/Ey55h4eHCoHkvsCklpc+pnTZ9X5n3Bl5XBeT5nTwpwEOcqza4lrENIK2AA1k
hpEoonp0R8nQgFEthUKcpH2pFKd1pfAzfFOG4VM834YA5IO1cqDkF/vze/fa/8OGYUBRfWApuhKH
Wy27ee1eBMUEVkq8ep9wtzY32Eh0aC6ZerXQlPRxFNCp7Xm6RaS739SZSWKVYlXqq+6NgemyVscg
t3rLpub/cG9wQiqY/jRcFYOxL6mYzjBJNxYkzGWp6e1+hBerzBRkqHm/at+wPVGi7Ri/STdw16Pr
Lh44C3jyrfJ5/GRUZTnESzg6SQ6ym5q4hIeyvQk+1TsxEk1Evffv9eMflrqBR8VS2kk8ae2HPS96
Gh+IrEYunMGR9o4H01YajOU7ydVeSjntArrPYrHuUhKLc3KtW9Dv0AUoMWf9c3uKbLKg0igsGc6K
X2B/PTPvqZYhyijZNNXDOBXiz9EV/wMbvmxCmqaaFxYuU/yoJKj/GpjqcqSehWKvm//WFyOM/qpR
NDyQqftDMixvz1W0u81M2UvZCL72KBc3YO29TrBX2Y+lXHtaDpW8rUZXVlvfz755f/ZHE9HyYQD8
/EMEp8dGI5QwW9cwwYiO6Eg2iaQixQZYoPlEmShkT8jDH4Tl64M9WvzmTS1LuBKxR7dLW/w8yIv0
LkD1kaAqt+UDVeN8idvQ1lp1O6sbPkhxn7/XJSNQ9nwaIMwg4HgFoQWEGERaWU+ve4fU+traJaQp
L9c9ZnilQZivORgAxorcCWUZ4lnL+A3huSYEIUjzSlegRJmTeo4zCriglQkfhHZLLBrtU7kp5dG9
Z8XXcNT+XxGmiCp6mMYCLn7hwOX5G1oXdg1cC3mSN4e8IMAc75NnqZNlO+g/j5/qic8ncXquWWKy
yRx5d5aGLE8j53jFAdHC1sTcv2WiYsqpLoUe8Fsu/idbSG0hQ5ub0OASddTH4EViNbQRBQZVee+S
ipbsf11FaPvwxv2vSxF79zlUjcDFmfOalEhkEk/w44WW5Bi+XHzZPyUN5IxLBq7AQoa7V1fQDoYI
f5HiEzxyE3nKp11xqfNmZ1BC9NYb/uz1uNISJJEPD+NfbGyokX3+4BKDJSmiai9rWZeIEblerRuB
frg9JoLDwaiNudsXSoPGypLgnN5MeDYx2ZcAHIeRT6BZU2KnH3L/U9mEDsxggMP2p9yp2lOYIR0V
hNdjXIDnd63eY9+6s2LlUUDio+Jnoj0bGE0LSODSbGSTa8OUL7LggeleHSFddT3uBqaJUtexSOoW
rzFacUp0YuLqfF98UCDausZJIHAU+XdmvaM/HVsQ+lfj0H10iqQmNgx3HRK1/L4OJTu/3+pycCNX
1EsmxTrN/+srCDC1BLX2iZhukQrj3y9MMMvb6/IkXfZOkxpcvb9QSBcQGAbhna0XGlDwnp/9WOmn
od12F6fL20/aaZ4wQnAnZtR7rNAlvGB8dfBWBk2njCFa8GRx3CZ14cPX2N+H1Tx6S2GTIvR4WldB
fguL4kMccYB2snP0ruY5yGwU79kBXQ7/8B6BtmIePzLLQoa4w3rSAbBVXJ7p3FUWZlUlSR+RNUaU
iICFkjHnmuNhj09tJeCfZo991vBf/3fgr/BmByxPvgxjwdY13Y2AhR0x58P/Bo2HAaBmAmW39I55
Ib333lEhmt1BK5w7qyzrAgVNGQ2NJsOX2e3dgBf/qZbTisczzx0WGXAfBF1ILIpSJM0hfXZtB1o+
q9RjHoxY+Yp5hQLY84xlAFlX62NL9qQTF2PFN4JyYFg6mDv/4TEFglJO3bnyrg7IUNT2fQNYBXZ9
L96CiwXioBWHPFuO6JT+XrTGjHM7khVdoRa5XPWxi5YeWJ/kYQWwHVbSpdHawp/XtUVAilBvFi8U
11Bf8RXJ/RN4uo91kSfduYU+uyCHqjSBICH0S+hyWd1cJ01flAHMjVD+i09DxFHCo7eA3utxP9jl
KSntsbvV8ZAcJ2eFYVVcJJDFy/oShiC/1qEga2M/7qqHt5xS84F+6O4VZ3uaQ6BNfxz0EnnUS4P+
YxuLzBB5Hax+9nKNmpMwynP0nJ+yXwmQOLP8tPOWDCxEx44keUeUp08AlcAINcgXPlCe2okQOLr4
18x5wpu4qzGPhS9q/7KueayOBgqhew9NA+CXYXvA8/SWGG1OWOXPkpI2GrVhksNjgYMb3SwNPe9c
lMw+XnMIICYzaIHp/Et7p3qn31kiQkonf3BFlBE5hIAN/TfGnIcj2E1VuUDLE4ALexglX6LAeH1l
DDXoY8TQE5UI6+yTfXSHw+anwv0w4dnr/Z5FEC93vOu2Ms85iuW6vwhaoCbXL1olPsNsV7K+1B3o
zFNSgoLIOZP8Pv2E1/Qhz9gLMk9zIQZKzHyraQt1CQ/f+NfsUjw/+TU2p4of+7U4eizXoA9GeIoE
wTfDJ2uGBAe9A9Tk7OFHnW+y8zrELBCFHS57U//Ufs5e7Ve2wZO2FeeUeeumarzB04eqDJX5EXp0
oWCbU2ONtKHl96BwsX/+7jp/jqfcLbz8Y58vDJ2m43ecl2ZDiP9O+TerFe8cRzablTluraUpb+0F
4fIlI3kq7uoeyCfuBc52wSajelr0yK9JPZtH+XwKRC4n8xftmTwQjciqTo0rOpwnC/8f8MVpyNKZ
xL7scevCip2/eZbU44PE9Po2cWvkNYlFm99aN60EX/Yrmw4ATFXzL9Nf0wR0I8JMYTomOTTjcJQR
gf8KEcCD4m7rkg06Fi3D2EwK5GTcNGDyfCvmK5rprp1pTKb7X/52ixwDFgH/fV1dGjsZnQMf4/h8
8ERYpZFgYMLan8OUhUuZwMnfbdG7Y988ZuR69XY7BO30dkZg93znMHz8RFISVaBlKU+zR00GpgRM
I+sxXsU1O/vSaShLN2XWs7vsBjfA7Uy0j1kFAvUnOjgh46AaSTV5qp+9oolI9VBUQFf5iqPGgM5a
glwn887w4nrcChCeCmd+uqDug2tWrCgWr/i7VQdsC65TRrlZOJJzB/EJ484k4FcDLK/bL61oPMcr
HFrUv9K+4NQv3+RIxdDIxJKBgVtPO3S9XCwpx9KMHqSH9Ix5N91ksSYopApHrCK0kLoNFCpVoLhs
RuOZ2F/H9jBSv4g2BSqhmGbcpVfkU0WHObD4XErtl8FSUaJVDBCJUs/aCE2Nvy1FU6bQPrSeMhRn
YMXNAznDkuZgm7gVsRFS3Of4HD/grBkS88rJXPJrqsWMZtlYzFVlKF3g38L8sKOiyrBLIuLMQEUz
iWtPm2D9l7B2zSkuSNOXQCAVVuIauf8smZNSCR286V/5Up8ESdD9Mlz1PvUAMDZh1A+r5rjkk3dj
UUjFGPGGe9cGefX6sglNmb9qwant+V2CfVXLSrsZUnEF53AkQyrKSMnhfIdl1j9vVfl/toaS+Y/l
mxIR6LK/VwYLgn41rpLf14yBtyyWkSKZSCIKnaG+yDLf9lO2psbSjeb6y6PJrEcp3+mzx3ND3Xci
40hVptKgs4H4+/4Kt8+8CZCmEat6yaacvnB5QU2Cs2+Dxij+gDyojclgHvKlW5jW69YkfkKbjdwf
LITblODVhIaeqfl6jmI1ayX9zED02+EGpRFlm3KwUf8akJzktyuj0AjoaI9z4wix35bzd5r8BdYf
m818l5/M0nNPtRTOXo90lK45Nxtg1YZYU3com5aJVkqs4J9CoUduiwwmL70iQccO3Kj0qxTgC2kf
SHykKSL0BU5tGKJ2hOUDp1YP0Rvm4PaynFg//poVT7VUewkKsMnPx6GAwUr8VFHeWnzYVpGuJVAt
eMbdNsXfcrvuoxQd0QvOuHylu8YJ4Ig6gyATTDmejHkROxGScPHxJJpqyeg1yka0RgHizLP5WOum
vuSFUXNePap/BTKoDZJaV1QAcWLp5+TPLsb8CU2HAtqWzrhJIWlfemJSDeFGyT6o5skgwFGtS4HA
2+wGG8ojhy34dIH4MpLKVsFU1t33X021mSatHEZ3W0oebHxaW0LiMvQrzHhjG11JhGH9UPCb9q1v
Bco6rBZ+TO2uv1ak0V3h6O/F/Uj38KBs/cd0W6v1PCBM8eVkcwzPoVsQeerJUmv16VRYQxAYPE8T
APB3krrAWEfBvOTMWEmXOGBoavZfv93pMiASlLegbTEpoBcOTTiSDoMbId5PcpNT9fKNkeh6qPLr
ocXYU5ZxqqSwLWc+8UUK2niw+DzUH0X1chlahOp1l6PmZZJvOoGcGDKSxjmu/OKCpYwg/jMgcCLI
kSz/7GO5uZ1A3RRF/jw2eE4qXnvql6TDx1JMpFry3MLIrZynj//R17KAmqycgDceAbkfHWaAz0zr
7wij6MTeFcnATU4KAKg1qrtpP+PL0iVkolpgHh2uZ+Fv6lnvHYnv0ASB2Sut38t2KiAZi2dn643r
Xh4kUczS6lFoB6gpb2DTsMFg9C3ZkyPPbmjPuTuT8Qq3hodK1Qk7IAlhz+GH2ptjjzwGSnqF6W3k
BZU4A44h0s1o6CGAEV4bmNZ880PZ4OWDf3JzosXd8u4IXiM0QsEqB6kh1eutk6+u30FZSq/ByLU8
mMHXYFa+jijyJxj5/+Ew1VpQtvOa/Lpo+KoeilNEpW9ymkru+Tyhpi20Np8q/0h8vYWMNqCnfsHa
UvOEFhfja6pspDIjuGJaAa2NSH5sApJgFtR6hsmwQERn9fz+CLJDLJqZ++Zqq8Rs2h0a3wQNoWgi
xVGTEz/RrM+3im8rYJA+KcrpK/KeGcT7/190pr7j9T0MN0dsRw8t13E2gUgfDmJ10ToUuf5y8rF6
NEu92Zp4jIpUt5Ni4nGUaUaWh7uR0xxi1E0Jhx2sD1fQVDR/v7MiszGzfhBXJexLKQM+tg56ROSg
+a2DeitsBxh5w88fj6GB4FNhQLahS1F9aRqrq7IL/kBgCjgQS4JRuNOxc5U2E7u3IcS7hSAYZi2U
PlFgxZDhtP1twui43LnsQx5TI7STGjFuAklTlEFpDiNmr3CPJRZ9SNKj4eR1IKSX1gRfn5YIh9xQ
ZQIBOUk2w0hTLSScKPFP8Y+813Yq/HniELQ9P+AWESdHs7HOp//ulCCNIps3tLFkA8JGDk8uBuu4
Pjo7ruLTZRovtIJcFlRufSHQf2KdAvlu4YTMbSAG3ACbwYJiAfDLZbVvXyKaVcSwpEBcm/DpbARx
5i46TgtVB8h5tq5ZYrbczrSdMVqKMnpDOy3X6Oa1T6Yd0bhRfoNpyEHhYzF7zGDhQXSlutWUpzuN
3qM/l4E4RZdGFWIRyC+Rl5mkEbQk6nHqEwsmnfJEVvrP/gKHuS2PY33niPziRQ7lLGWh4ZVXHIAn
sCZRh8WeojqyWIA62no1mGSJufJssSh6Ae2xEGrpWY+2uzJyE15zrQfKPGJJ5EBVcWcGs3xdunGB
r+As5xUJ/BYLSptbGnpaJuEueNM06dKoGgqogWY/iK2D5zhZ6umB2o7+Qod9uyfxKmdVyZbkRS7P
V2uHbQONDE1OqOL8DRWbrdW5C0ssXEkFmOH+F7jjC1KjMI0xdS0PCUj64SBFHmVMSGJZznUM4Oji
Y4+c3/Z3EZLGiH3pRPPTfmexB2Jh2PvPbhNyUAZUu6dRZv+odTP7uFy9yQXfAhjCjxeE7RQlCLmm
YxvyZHjPuAoWGqcquNTMwAE1Hx15SfyEkXsHmiSVwyDnoP6zSyqZ0ihOPmhWw7G+e+qJhzFS5UmW
7G6zx1ZFMqStfqhrRzrMnwhrnZnNCk3RKStua0nNoCJGFDaLdSJKXNmYJ2hsjXHuYMDDIKFCC+hl
fxp+KZsrcEuCqjE7XmQOZZjGZaRlignTV9CuMUWHSuRCWDeBb7SvripiBW7ZWSGbFBy/acvf6u5R
2LEGrDIdVYAYr52mRIBzMPEGthWuQtuiIM+Baxj8xzcF0KvqaZqV8YpGc2MJAukHCOEE5JnS5JfN
HN59tBUt9/JU/+sGAgHdA+Ax+vd5ISWKydyAOzqQr3hq4I5xZwBJofPBt5pCQ11upV5ONgoGrw9s
XdeM2Z4uJwVPbxqEaIs3EvjCmwuOM5YL7N2/LqBiSm3COSTf55P4rI4KHOaUdmmjHs66vg2KAjm+
8L9uwOQgw902CLNyDX/NaFtMJS2oSAvbz/bH3xsg9favbOrRE4B7K6IXTiFkVC2ZKx4+6Z2xwVsl
sTBNg36lyklX8VJwBovPPdElkUZyzle3vbJJMlMq7jGMibI3mB/VWfcEo/KXFQScK91SyBWaB0ow
/SqKV/TMDHU35KranI5ou2euk1O0no/RTahDpUW/oLapxv/yvpN6smR0fwmB7n/0bOc+ET7w9AVw
fMYRam0PiMRVd1pNpgUhTvzQtVGuVouIu6M7Uxma5wM4V2m0/xunFQcHsdgYBYDZh/KDcyN0dZ2+
F5WtIFKMfVkfhEBxfdZJDJixfSSH226ndGidSH6+swrpVn5/mnwdiJWhbuvOtedhetrn6TxyfDoN
8PzrfOUIzyEFXq2AavGcU5+SPQGb01ppzQjSN5RbuH5HOxwiSAO+IImP3JfdKeiFrqUftLjhnzJa
9m8KwM8WZn6T1qjVThsabU4I90vlrasLV/53Nq2wXKuRE703GdPu5QWZQfsapEYBx6x7xefAvIvM
JRrfScF45+DqBoGeAIB13/eFAKG1VLX3gqD7tBDGXSyph9idgDfscbsuAxjG6IsdLmNJyBFjXTDq
sZ9AbHVjIrGauUm1irPCMyuLahtwuVYaT1w7gGmdaCKofhyQveRqMMOu7OL4MmFk9AojqmvFgOAE
Eo4lRTdZGYvFWCQ2qg230IVguaBdimEKJUK2ly1un5r4bIORZD12EgFYn1N8d1V1bnOGHd6I4l/y
c/eFTcuDYU9tg7ZbX0GlIt67j1WXTfxWjDK3VZu6vyxWfbyNQZ+hADmYPmn3Lc7ye8yg/Gx1UkXX
/kTKp48e8ra7QZ03lZGw6i8plxy1gtb8w11anUNz/iFuI7BJ6dilJ5ImKHFE0dXxauv76OjXKWjg
rELKCmAy2bsOkao1wNV4axiRTMnfSkaxZISpObODfnw1CJTYmbki/cegE2Sl5cKEL9Zvos+cOosK
f4gBwvnvelrKMdXO3pxQ6yuxcBnaS1KSSQTWajeb7ktG+pzJ+dBz/af+D97KtDk/2BtUMjka8F7p
daA9K6LmoNzYH8IHGuhuTRjDtCaB65045lWQoEzweqprJGeRBX2N1QnA6fCQufnd9AtI9ukJ5IIj
CfKtOuKtAqUshck3zzHu4MEwfD6HIpOfb8qldrVaQiEm6iVkSDJOyF6M5NxwmlYdelW7qx8HHQgG
l1i2lthUxYVpVT9sjjzdSFbAdjfItlddzP9QI5lNYmJDs/6nxPnThLQnJFlKGPS3HwUSHAEtHkGX
nbbhGh2HCXW1bUJHwQz+nvbSkr1VUIFRZYb+wVrJ8yy3shuOPgtCSd28GdGYupKcjk4Ob7Pcvq+x
2daUFrhLvuRsA3hpBNduw0hHRsSbaf40WuiMYsCHfkecWp/w/9z+U8t5PYgzEu5YqsgV1JENsOlF
3XALjWkXBauAUAKJBCbn9Ph9kfTxL/dZgbzZ3toUYSCBlfuwW54CeQMby9YH0XxoQO/c8eO8hrmP
D5T8QfXBrtq1yOsuNKSM0mw2rdxg6Ns5FjRp1Tsy2isHoQTt5WfPuIjzNdHBtPjUCrle/0ZCzU4e
s4A1WvJKVl26Xr/FAMxDY6NNIrF9bJv8CeB77M28EChnW3ImhH8zG1/i7tbJVw3DtcnE3rY8qPwj
dalqkPnTL8aqoL9u/QffiaznU+8QVoLfMMp2EnV5idFejUf7T6CSKk+aLxQfiI5QbsEZCxCm6Knb
Upz3wvW8KLIHeDR+kzSPP7AIcjnnyAQ3D7bY2o5L7tRuIBENwEKMQLut5gpRj6cKXo4kozo5LuC2
UpH9hYG6YVXf1dgUf5NJeYqWW9mY2/aJ8YwOqFjPdibhoRuENNkeq5rdEQE+qhdnLJNe9exOPFXq
1//gWlKXPms8UVlW88HAitNGWxtZkQOoUWOT4cJHnwrHNA3lVIGoApCCN894GpA2ltxv9A+7G7TN
pPIbFQwKWmNR+IYoM6fZlIF5PLtb7G/qXckOQjrovYOgXWkO58j/3as4/kqdxcSeP8Unh6KUuRub
c0NIumR03iRgREWtvIYoc3T3NcYaRMCBDN5HusWaS6p9h3PIx8vPjlUqTHOmuSOn8+IF3ZO8X+aM
E9UHInYTFlygXUDsX45MOSrHL8sSKmA4sXkhEJvO3+54/qNdWhZP8C5vwuXhj7+D7b9syidS1HBE
x6DhYLWeZVaayKiTs+AXpd2eQ3q3dKaywt0WAsjaCMqUdts/suKOI9FnzzLCkCjNbIMaYU9dKiLJ
bdSdcOfqOOJQa/fnKGXaJErmJz4BOtikdgp9qZ69KWs+PkMvFF8S+RI2T0k3bh//anVel/lGeY2M
z+VltVgLiwGSqba7/9Z+Tp8h/vB6SiagFe+V5uKFS76G/h13aV/Pjm0dduQ4NC2777uS1suGK4oF
+dOHkKa2S4dPHXQgJOIjyn8fqvMbpprc7Vsd66STKi0Os6C66Plpd/3nnfR7yi0W3Lg0Bk4mtZ5q
WJ448/nzvhEnZ9bXhA9xiOcA7ylarG/9gutTbKzcHBZfJ/ebqd2mZByU2ixVcdBYdgGBxwnVzXIg
8nJhfOYUDqNru4adrYi9x1u2QLVGpy5Yscv2jxuOg1UiRfkvaFCNH7O16bn5GIiGe5fhRaYzgbsO
5NjRhZejR9JCdzSP9+H6WRGGdBf5Z34V9sPVwCjvw2OSR3PCxn5uUYw18+FTVnoYXQalx/8WgzhX
fkUIJGdiYIBQCyhC7ym8CLzzaQukfpbUQ1PkACRW03CjoMpI+aXJ91Bt9pjUXdyOJDHmslVVjEya
M4D6HMiUWPY21Zpal+sRvk6QytLAaY33KB+BsNElFPnUPnKtt5694j3U7gm0yW9BS5ERjuPEowVI
N5yIOecXTuQmV96Kva9RnKyszrF9QXPhvfm9+VAdh1ZKNH9O8+AI4HY3fuWHROglArr5mypfD9eB
tfB8V5ZnfYkEWbIroZOk78gQVCC4gtdyHzfFLrjrtgD7jSt8L+gJaV2gw34P5oxrxsiz2qQdgQ5n
96uZr5CaJnHvwC8+0q6NoPO95/JBV4Mp/ohwSdNMHUfZE5jqdqzms51Kd4J9+vi+zPwXbUTlh7gh
ELnYthP8vbiKqkXZvv6/S0poG4bE/WuSloWx9rFA6RIR5ev7zsBhAnFUl10tHwvHJQP1zUebg8J+
BP82TQlyxSiyLKSaL3g0b14CmxgVvd2G3WlMDHe2cxj/AZx9g1SKL74bMzuF9IOWz05+sCM3a/rp
fBBmvThz5uY0A4JAdMlHpKZnXqKkpzBgABW2kxxzoun5aZL/lz1Jh3chHlWH+vXra70J0D03K3cJ
uHFWvG6yTQkiOLqnVIw/jC4cLCAsIczUJT5r9OeSGCOmerzZhFutqrDNp9QhzwF/bKFplMEMpC3s
yn4hWBFOYknGqoGnkjnRPVk/GwRLHZE/L9WCHBySrLfm1bHx4G1Ka+z1qaPpBv/YUq0vEjutvcRb
czU9oI+q9IyZr/FSp5U4BTdZs2rV1rohz4GckexwMC7d35Gwrdo5F474Ue1QQ1OZBHdl9mOicNIh
vAZtScJGtzzi9S5xflOVrXm6NfrxDH77v0u9HbSTyJw7ORI05J2DBqJqMs5m1EGPaRWKYwWPiZDn
0+gt2qSBEML4QWDhSYDYPJkDc5DM/mDwfjOsTCN8LTFWVYg16vOlB57iMGDoPbQYOnZcMiCEU1t+
B9cBxnw9I+QDGpBJUUa4q9eFUiUT4QNA9BMpo9kLlpbppE2pEQhem7haYPujA+0hZsCCQ4SNV/SQ
MiKsV6MsZt/6y2oTKOvTgwOFHvq3hGrS8/PXw/lYQbGMQCDEvTajslY9c19wvzdDI+Ot+FHoQuws
ENq8snYXTrtEPUhJ9C6PMJtzel0uEHK2H+/ipsrWi6gaGkmvM6Uk0nf56eMs070/u063bJGrYQqx
bNn58g2UzvtWnM8TVJXm/8P/16o4/phM4NhVCBZ3nswvAEcmGv9hlnVvs5q8V9/1W20Fmif05mNS
4bzpXfW+dWGYN36t+ITI+/SNQp7Ssn9etOrGdJAf7vnw2RMkO3DYzmzgd++ItS0fVJgUvbAI6V3T
Po/yEbe8niiFy1eISn5GSU8Eg93Z6duCf4y6RmPLzct0Ra8Y0DknsvyCB3EcsEEDXr0YViNmTomD
cgeJA7WbL2HQksGEJGwhIiafnFdBkEvZf+8L1WSTglPNmH/Zjkc5wKb/8N6Yn4C0u/bXWfgVQTom
ZgK3JwR1/VWt9AVHwEwws5EL7VKqvhUZ7LhcbzW8sKl4gT+hPqDAGR7xF1/XeeqVGUUS9ovfBFIv
qh2AsBnbhFJ3Lsk86w/81DmHJhIzYuHBVJvc8xiKdD7v+uTva9bJSgJNg8qWRgRNDZOM7wvKyuTT
Z/MuUFNYTG+/VJ2ltWJA1himoUbSfeOtJK0LI7lkEL6zXuqp45/LOBx3XgQ3Ywr571rlMFYSd8c8
MxdGhkk2AmAnsZMiD/Kxp+xihp82KX1CgkVpHRHVQmAfb9mzjj3XO0hVeGmnrn+eiPBIRVI8+kgT
fbRdffLdWYA6D/h9eIjTMr5pQ7lBZMsPHMy7xbaNcDf8a04wSr7C4yJ4pS/TsfGkuh/3JsSK/JeH
ZQnSWEfT3fM/Q5DrO7Ofo+hZThe7nBFAXUfFovwakttqGLqEgunocjRt8YsVnw9CqnCJeNpgtJZ1
lwD0XpHuRm57OIaP8u53+P7fQCZ/wd3EzEydElFWUnEammHdoP0EamTz7PWqYV1W9LwLFfu6xIO7
e3sloXVQo6ivxqIJ/Rc8fq8fX14xzaoKW1zQtPyDnzbME0UvxtrWfJRDMmk0zVDfOoGQmAv1Ry7d
nomueQJlyCGtfrCVZbhUfRkK33t/ldBPBL1khGGBz7rtn29E6ahHy/XQiPMM4SRl+B7GPepP6zZA
yPbmk0SHavo6tkAOXLTFTxrgxmHMS3nhJs6C0veoC5vPtaUtUwwHDrJxf2UEfAvzvU+8osXwPd3T
3Sh6TeXiQdCD5KfN4dUjRzbRaTmVL12/RlxpixKogdxKtO/8kro39hsAqtJNvwOgwGW2rWsxQkg6
hNJ0003KCRG8PVNd9p7rxSvZ8bs9gTuhlhCxoszf+XoG0S1G/R4jCLUZowFQIiwYYZqon/qRKuWU
EBWVhagNUzwAx9KaBpNmzE0ahKluamnzcSSk2iZQp6vPvIucudsTNqZqapox+1BdSGna1qbCfQ/5
j0i/yEbE35W9hAhhFmrfI+5F+Vuqc2iuOUAvyKSJ3Jw3TJ0adoVuOY/B2d38JuGlisSomxmcpel1
G/PtdrMLXOgAJ05aLVT+OfRrVHjulIYm/dM0yghG6xiZA36KS0tWqzkMbenpWPQtGLojkTD8EBzl
8eVmgT2yxp22+gClKuY7puZsD0WyQhCQ+61m0DAzwg8ECZJBPe8aF032FwtWwR5AataCXHDqmbcv
y7XPgVCaunREgj7MFVVeblH0ikRbt3AFul3w99XGNmiRfa2my9Ac99j/uZ9yVHc4DCLv6SDsw9YF
zuWoZ/PO6AeNPYzz3xPT43AyvjObRSrMGQqqOODLcaqvCYzJlGpnR14aWE+4aha1ZUynHkJx9ZPe
WHy/7APt85kBIH3/5299nZOP+WnfrWKX2sWzJlm5rtJrCLy1AAaaGfUkcY2CdL9O0Nvl3w6rvGKq
lEMF3VCprpeNpm88UqPBACuOSAJc6B/QO0RwZEfHm+m+PZ9HRlOkgek7dpnCBl7FnkShqu8/vK8E
ilTzh6z8KRdr2KzVuCA8xETzxFbkPun6izRW3dtpHYDTHPUf/auknhjT3nKOs6W4ooM+Z4lY46mA
6p0hnGjMUnTM5Uh8XEuidli3mXPGeHmnOcCjnQXqMC5ELVlcfcLqIGv0/vYCBoTDt8C1hQuLMTsA
B3ruKmJTOLF4MzQlnWy3CDXRHCQvyT0rrUhb1tviJ5kWmHyqfNu2FaEhrqusPOTaiqz0BCbbAVCF
oOaidXmQz7XHTQ0gG66q6/L2c62+3vhbIWv4fnOz+B2WSMXJ8sfpct8kXO/vzhNDRPaWB0QJvPhh
oAfdQ1bXoIdzyUqIJ7aHuUTFUgDGo+qDYOSlHmMr0hzQOE7MDr3YDOuYRFzaf+r5EiE0YZ2f/6Xl
bwm+5UJeNdNXZCSjQsIg2aJF6q76/t62Vxz28ylGzVWsbtXo5ZDCkHgGmd+YGlIMO44ohLu3V8fJ
r6rSYs8WonDgJFpqPcOC1q1B2sepHfctG2bsWESLo2/xwOZr9X487W5jfXt4k/XjmUNMMcxm5bTq
gsJNdj4sG5FJFWbVtVJ2I0fq3rjyXYWlQoaDbD2QIq4IQ0n/zwbkjTcFQ7NqU/p2XqSrN9VNhZ9S
vCZCTRVUb1JyeYi39aYzaO5g3i9RSeUeIcwekguwhplw1bJXrfo3ceocRQlugftCBpSDv+rXOcDt
WOOxEceLH8jzuSVmjjrgz9/0HnF30j5K39VL1+5rRMjs/ZDeFbxMAYydl2FU6/ZD+p2YfvQUTMFk
n1N9RZTqe+hO758K50zFtrBMJCBBGDBO23j1sQCcR3hmlBXsIdFrHfw4wgOcgI0tF5NuWYBclyAc
vqmEN780+FSdLEgZhlYa0BAZuGD/FwdtSO40UKDyNVBTXnnmCbCP67ZnCFvel3/o0q2JSw7zewgl
wxBm54JvWTtVb4qoILsPdlmwlZZayESbv8SVR04b8Epq5U6AAky7GHbDX7YMXBGBqzPtYUVAEpfb
QLB0nL0py0OIKXYtZoRkXa+RwBbDUmOJfJ4JSuoeskRi7SgImzFM01chp0OZ7Qi22/36oEiF37nZ
vfMLhwKz+SY9EqzM0I1R7QcPE7L+6pP2C8tB4PH0qGOvmLr454n/XGUeJnTQim6XyJSfPAw+eI5T
hOfeifF8qDeiXNjZUBekkNaJTEMsNwFhQ6TJsEeLLJbXcRN8wXmYj3m/gWY1OwgUYPqmfM0nMwZq
QFGx8D9dLCvRk+ga2Z5WCsatW593UYfy55i3avlcxWezKse0sNxMGCF19x9kMl4ppIKwhu7i63vg
vV92XsvxuJqq62JfWM2kdPw3P/ga/CybT9i9QTeGoXHwH56wr0zE3EOXEIzn0SoqKbwadpRds+zA
N2e6RLNFjCavdy5Tpz5ckkNmj1FE2U2erQOiI8KL5MTsquWfSZ3+qxOLF2eyRcmqqsxDXIPhaEdP
FTv7geo6DnKw0QldejNoshumyDRGvvHsd3RQBqw2rAd7tXnRUqxp5s/+ccEzWPlm1dpJzF3wMC/I
GdBPEmsSx5Exfysd5s321ADZv4SkWcfk1w7aLmskZGXZsyI1Zv+cycAPDu2oOXfeQWvtEzQDg/EA
ZLATaTKY+bEKcavvsvyHLPvNwmAZxF7AI7btQZqJAggH6AU4XztA3VBfocCwzE8kTil/rT4tt70t
YfmzMnmGk/uoueW9jY3xnqSHYPn4JVCYOunVmzf33BffSgu41Sx/DQiqTH7rzJ0cle44PXD0UZiq
vCed6XszYf2Q1ESQ4+rQKvAAPN+uttvPuomDi6X2/HUHxFwwYBZrHa33yYaxWC6h9AEAmU8Z/AV8
9WZsdo5VVK4jmCTH6cZYze2piXWfAiZc/C9kOwratuZqRqswzoQvI1Cs0QMZ6M/H99LRWOiULIQH
/Joe5w6FRWoDXx/MkrYT+XFbxwkEC8fNUwH50WlNJl688AkPFNFPIWUsW7zSGwTziIgOaLE948I2
E93eeThncxc/e8fIKS2TgY1gk6EuspHgMhnvnfaBLRi3gE7s/JhePyLxzYN1H4soUVdwbPmsO/oM
YPMSV9UZ9ppkrGvW2Ca44ZWdZV5kOI71isqYKo89EyVPRPDwzQWj0yHCXiUisbf1FGBCf8DQsqij
Bl7V23hFzZE+UosAD/L/kpWchounOBkHpZOXQLvJWFpKtQZa8S0jGVp7+ATKx+M/Z2qN1eUbTKdw
ZzoZ376615+d7q0/U9iinDnOyW+Yxv5A64/GDdpEXi9CdMW+U6mzH6cihXKCDe/eSz+HR+ca9ViL
ChnXCPbBGB1G8MkUHmz4VeT+Df3mYJ2Rx+/C0pEutlQ3p+0mfzdlUlaG8QOvOT0vEh8hDHWIodCI
lJSyu04yffzqQRxTl+cVdEhZ3A1Xykz8K8iGyHnlE2Xq9TKCMe7XfzwDWZcSAoFrGTuVAQkhIN6o
GZfytCfj7U25v94UYC9aswRmLB7pWbU+3+/0FnQw9lhxZzmClMn0aatHKsbuX6fMJ9W8tOdflrQX
ptCr88PDNelT+dH3yaoVwPVF/sSxfiWQMRmav6tdyuXcO/ebN04cehuNQQDYyYWfWM0VOj6WgK1C
gTQDbYcqehMWqgw9m/HZpIoGuio3G2oAX9m/LSDbs8Qt0ZXFNl+UkTpu3rCHmqmczZGKQ/vy5kXO
IDWt7S/IawMG6M727mK60jfvk85fkzHYk10nQs7/rp/v2LJStED1jop+dv0eEPQESE6T4f94A5kl
dujEh37e0FoOuLVZ0inqaaWeji8lnPB78bAIf9kZPMT+rnRPLmsLY8+tMj5D38OkkeVoejm4P8S+
6XFsdeRuWIIuKyivDCM0t363+t8o6ZW18zy58pAWWKhmuzRicgrB7Gc99mE028SxpRcxbbLFSzVk
Fk2d/vFt3t7atN5e9yFVpOvXe3KlxT+8Ew68hcqYuyP4CA8dJ0mnLWoAeYdrnMqXeltRU75jLjgG
w7IgcG1m/NfbtpvaLKpvcxJhhtMIv3hvZi5bhJu655Q0H/jMaoE+qPQwsBXf/vSeoL/aq3jblJg7
bl4ICkr2h7QCEr+UqJQssANPITiscf+y8LelJkDahCpLs9CqC+lSY819ApUIzLBVx0sdn+ILBarA
dMIpoKUfJA5KUAF0KnmUQj6UIFnsjxiPyNvu09wkispCjmwW5a9hLUFJKgB+RGlX9MDP4apmtB9W
XaV6F//ciD2ZvtVfkJLjanS8dH7krU2x2nA2YhDEc9a1pWHbrUZjnK2GzeqIds2cl78zk/jMiXfh
4KbdskN++vW1v70z4r4ERBO8pBl1uf5hkEB3GzxftxsF67Dc4URJjbaj8Rr/2gxwEo6vg01OfzxJ
7swlOSR5XiMmWwKfT/FpT0wAXWSgtEHTXt6n+I0Df2XdyQ5Cv9Kr2NINkYG9BmpSp3R78+Y+7/Ll
/sClG18Ol5o+VDZ0yQq+7G5hoVoDhtkZ5Hj5hXtGz72vEPyGX3LR+8IwspRbOFMAAFdhqsw7RHd/
Xzq9Sk6okpZl2zdYcQ9zrDzfCdqaqhyvWgmLWBIowZ7gt3LiNhF49+DMYnO6rGFYCNnGYBL1y/7U
9RJiiSlFjFgFMxt/H7RAZRY46YYUT6chYIrcAqgvns2gpw9wbBfJzoD3iPu1H5WLLeXoOzNKmWLZ
e8vdu4IQ2lBjRSRvxjdzfRnSWOSfZQ6rPNa3cKn+ikYXZEdDNbAHOUW47JNJ0YsK0Ddzo9XNzqpz
Wy2UZBhX/Ydu22DgTae6///Hh3c9Q6370zyImOOG0gmTU7rbkl5sZo5IW/R/b9YIZ2v+0rCxAR1z
MOs3VoHEpXVjQ54NqoEWPi8sQRp/UASgKEEhJA0yvp9sJyU3uy48ircovYtPdsPUUTpvNFDtj9jB
qWHPx8PDsY2vqXtSscMYeu257qIMU6X5ACJAi9Oo8SvsvvCyUpgbkhDajrhh8/ZR30Wdz8veersZ
sv3V5pPlF0jlgq8HRKSB3q/Sdw3o3lXZnIMsyH5DV+EF7vYCG16KQWQGV3LNEcur32xnWDBhyrGl
XoTzKfPAiwqhg1eU71ouhEPSw5m02Wo3YsRFzusIc2OVZxMtwxHTttoMGKLUlksrSI86QAfPSiCB
x80wypOWRlNDNkSBlRvUNpwjEEqEwyrsBibkr6vhWNJvrFO2rZ1/syw3Uq0LKngEbjmqaeDpZvF+
KDgBU8C4fVOh3NwE+OFJjAUN9blIkLiKglYqyHwK8W3PFTCgwmLJg1FNa6SX+FAHgiUbgiZvqn/p
vEKCQeAOakGekouZWIapiI6lae6gYM6UNvifGPlwcPSrhZJJIBFGzMjJgNDBP7qopQUeZnTpSHQ/
dA1SQsS/jBpzF7vBjAFGToV/jVSlPSNMFWbB279GmWaohRzY9Omk1y4aLgUW2PobiZUbZH1PKyMn
Z55cZRJRyqaVyYyL1R/r01oC4VpZ3KSz7bwbzyqaDadx8kX88IUWFjPGBT/EOY1axcahu4TXRfnq
aZl+UUlkXYF3qqXKr7YAJEg6W0HBMD5WuTegV/e7dP7/gLIokpW4w9pFazmIhM7VRWu3vB4FvIQX
XOc00v1Yc133zS4LQOTeMbClbGM7dGl0vSY3dU5Aexuw3SfcDkyMzhs5k6wtO+NlO2J55jW2pxVQ
4awTyDJFq6jCvXN7z3QmgOEvYEaJDEtkzpsl2/J0APByZS6DRDycGLyPE5LfuOWcCdHzZiFtG8a3
eqGyTrlYmFUg6qUKsDriq4ZstVZ8o13wZBSqrwcpjMJPtUOfYHr3HIoqQuROpKsy3Qop5MEdZ5Yb
DH0HG7ZJ7/1M/exYEqbMTnMVMNpW3FMNxBN15j/7doOOQGY6u481O/MbqxDzAJQ2YVV7WX2hHN0f
BAgTKpZt9wIOnxc/lrOwBUHc/C1qHte9h1F/eqvc7wzwFWvO1JvlQDKk9Df7wuDBzrwWCZ7h7mlc
h8Zb6w2KwSLN/NHF4NR9cdW0xRaQUs0N3+LoFeFgXpsN8/s03wV2QPPEmnk5TifnUrAVaNHoLyJ+
yPCfq82cG+Fl/iuUoBHozqyjuXysc4hxX4xHokIknkudR9s8qp13xzQ03+FTSU+Ncq7aLyMD9V32
oUHHfrp9D/U81QGaHUVycHRHRcSi+UytwIFVYEf9OmeM/+Y4Q5MnwGF90JVEHu+kuNMGRifekQD6
6qfMK5OTP22jsLmPdR+xb9irt1zL77EnkZW38Uztx+uVQlm/zSdsGJKvmaAm7ZjlUrJyoqHO3ibm
7jCZk3aLs8OxKRRri/ZXu2AEroyaIsNec2H7GOCaTS5/O5G8cu5OPUGd2QA5NwIcVC6SWHjWADby
+SJxNvQap08K4KK5IybetHgn3oYTU87agzYlZjdJJAPcEv4p4giFX3McVlRJAtGd4gWkIbAmnWTq
PRfR/tnUr9l69KacPn7+Mc4nCaxGKA0lvcP07l1U4do/PZIe1PLQjg4PZOZDE0kchAzTJoj08e7R
5ADhI0N0o8SuESQqbmEi+bOkXNRq5lV8ZH+GC0e1R4H7l1TnXezkxITVPAfvWsE1QHGhYVsuDwMR
wZg0jry61eZx20OwopwCe3MLangYFCcsrwhteEYI3qU2YkzcTs449vfoF1piPnJEB4RFyWdcAz7I
sltl8CRs2BnFWnhxp7BtodComOY9BCWFl6DYHjOxJjzD0PVIsp9RISKFPly+nS4Q3e41AbzC9lgD
9Hkj34p3ig6qUFQ5FDwU1pFuyFJre9PCdY2ZrQnVUU4BILyL/al4KqSzTF3xAmqbwNk6TWpZ9JJ4
A0cntf4e/q8zhvnMYBLSgqv4B6UwNaV9aGzvCh0Qd4Qgi1qxaytan0UL/3ZJxLGBEpGCPogiN5d+
UdaKytI6iYcXxxsxtpCPmuaQsD3/E5PSRYq9K/jupxH/V9QFlXv6uc1ifjtmWd90IHxhc9hMuo5K
rtfmgTxE8IhwDogzcftFHZ2qK+np/A7AEIUbUQ9dWXozQQPc28ojEzkzxt6kkJiWw+WLEpA5QCVr
qHYDZJYir7uBkgzx67Yg7dToadJNAANP1cdRRq2YHEz2qTUev+aBh/r6YkUdJZXhe5a//1unvEEY
1XxeyI146abxoOkb/1JcBIUayvjU6mnSHYsRqQ6HUA/kd83A3dIFff9+0QfKuD3pZBRJPbvCgDIh
XSwOElQOAgts2cC+1n0iaPRqFXstX3gC/0tDf5SLHYkhDNIPajtclsEbFJYbpjdXb9JA6tJtU7AG
wV3WMG5yl79Vp5KR+1YNzbFQBy/tNxwODfImHJbm1j2Lyxcbbqy7mpTgPh0gbLtABWUHBeHbYW+y
GC7zTab03Rn7BPVFC+SCOD0m6AVzKg3NprzzW8gt4/2o/vJQIpH14GkTV6JHnA5tOV8DoWHwlRda
+6Gz4wXZNrFMZ3LM/sTSrWnENq+r8e7GVJsrklu5GTogxI64KRdXKy+0Z2bzgLffbaKyvu0E6X6H
h2Zk4qEdaJ8oLxl7J2XASld1SJjgH2uoJeQSw70/BN0nAmBf4VPtvXJ2Qxm3ZyBsG+qk2MTdcvPh
hdFfdh2rpyAFM3EOdd6F28GdrgkfBWfph7Fv6ELEcxHUhaitFj5Op8a6TWtp/cQtYtPLtuzs9xHt
hWCJu4UOu/0omDqBi0srN0JchFKCkX68xyYPDAcU9fWGshux2Xs1RVdEc95mKUU3s6Do/RncqUrV
k4NCUNN5w0XqDlxclqsMdFT6RlnppPwl/ba2cmQitpic1i/gVX0wS7dUHazHMnz7zYNW8lzdmvLv
Pf53+Uoat3lqCcZfR0FSuFroBhehSEo1HyPj/ipiDcQVcK16hYfHmOyrc9AsWBLPhDvIc52Wg0UC
UXcxRsBq0ICJJDVsHqNFtKziF+ftRbeQnSUS96vxA+QWrPcwJxwlS6ylLXbWTL4qqtZslDtq7d4/
yDxzcgrPvrg8c79EuSsxH8zntJ8YfR7vq4vrBE9oswGr197QtuoCa9gtO6aAA48ftprMqJntAnBb
6ekeV1r8jQFSMPw9EV6vmcFTyzu8jbrY/UXzlMJjZ56bpBTIS4fvvYmVF15ql1jB95VIoZf9Qqjj
6pbro850120s1J6ogLFrtrKZovBhoe8CPoCri7ia29BdIlKZ1BN8N9IvhQ2YQCbUCBXbLyZ3OXoZ
5hCPXAMn20D191KA/GFlsSnIodts5qn3H1/ki0CmYWbydTSErkY2fhlASJdjm9JfJ+ZhuQQQ09jn
ZZF1TZF/XIt3PrB+rtIVLK6t2nYTzilnzkoYljumBlMDNiosj4bH/9T3gcB12Yx9bmuMuhKbfHFJ
3z0MOwaumDbVyAdTVHOKC3OLf+5Ott8l18YjeI6PjBonltlFeNExIx1v5FV+7J7GREXLBBTDd1ld
n4io4PJCZqF9h4+HnD4UgAwpocckHWGAaAEvEAI9mSx57PupgDg4bkuM6iSLM4wdXGGg6pynh/c7
gGIhJHXKezfGaZSUCHmFL35w1QSWulwbnyFHVf86jZd1yybpFzD/QJonj0fNVdUZWUwH8Q76cGB6
ET6rlR0W7+5yrz8KrZ9PQEqG45oyL/LcjuDj9mOqrjTNL84RPH30FSy3NlkAk/w7YK7mx5CnvD9a
2n+BKyI9V6VPT1AyEem0DNVlvNfnAByilkbmLOLjsDsb6wsRnPYe0t8C5j9KpNs8s2ig+L/5bxRU
EOOj9H93vZJOpsdpgGkDDcSzyOUuEadwAr7Zo27mIlvclaR3s5orcbn+8KqmvuD3MrWCmUTnmjky
coyisG3ttX2Goi3in8mM1WPda3mr1D94FUzYbse6IEnZuk8Rw3mC+i+iWxXJrd4wG4rR/bsckFV9
eirFqXTI1bWnwx1Xl/kbFdGpBtxg40mJ4Wh7ReEY+GiI2Z8WvTcRFMeqnNzrMJMBy72OM47NeEoz
LYV26i/MtHw++GfTNawze1vz92fcZLzg8yPp8U8XiVoIimOvtfZkTeJIVKO8BDLbQRPm9wS40vqY
L1dGkW5VnwYjwRh68HYh/wKyqPhn7L48gkCOR/vFDqiNuhs/j4szQctEqVzINGgWFc+pwEuyDUW9
zHK1DTGn29GG2RDabBNayceBksVOdDaW6o6RKNMeZ5zzKF/C5N7ozC0X6Sh4wscBCHOJq8Ri0+ps
V/GI0Lir1YhU0jJAMsqbO/KR0v8pWqoqJWnwTc4SpRlUd6MchMWXFBFHLMvrlWnBvGVXAycQRv16
XjxEAOfc5XlvVjmydmnVV7fCJS9jKA1MVNrSpYGarQee1ctD9IKsQvyO+ce6VAUF1G/cy30soAH6
g5D09Wu2IuBSU7fjQO4bXLtfVSPCWpp3elKwlyD5HN596neyp1diOU4owzv36gSrNVzvV7NZxtkY
VAdkZwO5Ie6BjAwjPgwe1hMkmAHVYbKt/yHgZYjXrGPAnaZOq95Qsl9WOF5dFVcw35NGj8Ccb9M6
qmmWyG01DQ9JipiFJYQ947fqyQnKEOuDCI7GDAl1IKtuy2igWprf2pDiEoR+bIPUZrrNRW5/4lug
1b1ZVkE/zzf6aV+OOWUNUND3TVxjCt1hAjZgzRR1KVOFL49IE7mu3+eplwNAgBiz1MFjGf1mATkO
H+Glmg6MUtARSiPBLY/VZ5YLkYdoa0g3i1bHzDFvd7/EBxgrEbyhk3kaFq8RPw/Du9uc6mQUdzQk
EqvSnyy1Fa478GCbq1UK6LiHr7X+rXVOYXz6Dyjn0uRDKmgQ7fptbe8m0Dn3cWO7UQHzfdeUedt7
vjv5prPzD9saTZMPSoizkiVhtbaCliA10prySQHbt0jIQ/DbsZCOOb4NsNHNQsil1uaTfx1nhpKk
5yqNCev+yA+m0QVoRnZinojbkNgCS+pWY35D0ojbolGgIrPRjlSmMmxvDSNBTQ9ohi64l9VufFl9
FYnJB/Jb6KjZojwNxALzapOxvev7/l4HvqnTTynR8mAq1oIQdAp2pbOOyLfLh08kj5D6icD75+Yf
+aHKZMV76Ya4m0eqFw6tbsRxX4htUR79ucUoXt6LgOhmTjiUV1dqcIMNHELoj69m1ZtlhmbMj3fi
nHVWc3C5q3wQYoEAGmTClrckSOWQUaGVkv4UZuY1/tAlYLVa3b8F/h64p0YbSw7W5QqYCnKHkGkT
vNENO2rNgQsopjEwhSJ+cBnC7AqUQRDqEuQPSRO/OxJi2hdOr/rgZEL55UPGGBFHtbKAdxet4bRg
p6G9VDLtPTrXgfz8bh+4/3Lv9uh3IkJrzAqSaQpRJXecgzyW+jTJMS1tMB/EEknFYaoWvtZX59Ux
OPMTD7UpSpI1fkpVA2zgw8kJYc/Lv9RDBZt34UahuREJ0d3eB8zlAf3JavwIM3RX/hdqKPatOvFS
7YkYC6H73+gGARufGmerweQ1wisnNDp0DvVbwKBxbgxtSlzmbCKglbGr+MQP0znH6tpQO0gin/OQ
687OdcAGf7DRJ5zA/UitB6EfAdqTL0+GXh4iZvC3R/NcYiKkIVOBJlWvHlqNcFennOFoU7NI25+B
qVj5ANqFNQT0TQU9z3CF88k6I7ssUimhNUV8Y7/BgDnvJWDEDDYsvfxjzbx3oZmisEIvucSZMXVi
gI5PXp7d1pw30WUjGbnjSMHstQPjXIK+qaId3SVm3hAk0Uo7rjPdscH6RmYu/TWQDgNbDOV2Vm2y
Y1c/lRklQdSnGpnXQ07+rd4nW9sRzB6KNJRw1ouxjO6oGYcb6Ni18Er2GA999/jUOVhluZn0lEGi
yva1xDPQfaURwS8pKyMCy3cuZEjNIgDlERL8I3IK/D9NlBIXIdqkOXQsIPiTXEpu0AFnCWtB1x88
rY4ObWUoNmTO0OsNrGW9+NJDyMdvuF8oWAoDjOU1SZoCoVdLNaMpM+06siKtIPS9M7Gi53+Ty6cY
l3jqg/9cIzF1oB4Ika4Lac/m2RPG+ni2GD1F7N/r0XtK0+L6qMHyOuPEtVsO+k/U6qsacjnZybhj
RbeEiWhlPJYNGuM469gbft6q44b62Lavyrut7V/il3lPrM1RjHraeDpvN2kMo5yohsFuLmsGS/kV
iqsPNTQE9EX4QVTDd3MVpLS4H+A2RweJITn8vKmVYtjYSEappIY++eVUbmNQVR+42gBONqk/s4Rm
5ldgT9RyhKi3kpsrqTxvHfBk7M3tIjoz0Cv35zNB0HIufF9OwxC32N/kPmjiYS8Upnql/yy3uUoH
8RPv7pjYWdZAyOgEVN6C5Qcb/dk4U7/66TCB7bbXzqCcCOGPHGNj5VH5vqwK0AoYkaqfd2a0VdDE
VnldlZa+JOkZIvSzmKmxmGczZ0h3MsXm7kWnhKTG/BwKlfh1HdXbJGrHYaG0GzX+qaAxLBuXOvJM
SZvHJESPLCJbjW0d4J6E0v7D5W+3DDmUdZOabpdLa8yGa3i+SIhZnFXegjPrui8WXPE4eB2HIdtl
/j2tmq4Jq2AdJ2SC+ovFSbf6O8kI4wiEAnFD1XkpV0rmtuzJH8sdaHJuMmV1YgFw7orSDXIxgKu/
TqfSPfxAnZLoh1F/FTbK1RQy2hjJ5BHShHnIvYlzXpbdZ2BzuqzUi1Vv6+U6HTpZMd/PXNh2UL4E
RvgS+cy5XL5GtW/Tc+gDwdIzdKygI9KgsT2ODZHXg/DyShJMwA0O/XdPYuf5VbrkIlHYjPTpBMNZ
3DLZ9+iEnJmitaCztRQHGkfPiER1Hhi+464g8ioWZxifnoA4Ob6FNDYd8MPnmGgSAisXa9m9KHAi
YyjlLIRcQohDflIYMmaF1X0lSiRgzTFucsOy5bdRkn5ksiL6I1pqk81tUAzyzO8Vw/zUcd1PxImF
VmqDXNGAnP+zdb+/qIgxrj0eKd/ARUpsQDWzf4X12fO2Oenm5KPMImVeU3dN6ZxX3Kg4i4StC2dG
tgRVlQR53IVCsDQWgUz2+ldldwp085luWoz8iDeiRV4SqAXUchbBB63BSscROlqxznEQgULZyAf6
bo5L8F4b60fGy3DdOcq5KtWUVEXAwz3IEo9zNa69tgb8vim2iVu1QhQbb/gnXgmX9h+6NKIUzIXy
60DhvXdQ9QCg82/Ry+5xHSmQoV9iOCKJdGetU3X6wzVTt/S9h6jyESUCyR1lCDcTccj0GD+xp1W3
yRN55GI4RPA4TOT7ujE6tXmMqRs4NWb+7uGH2NT8FexmoG6zUFV5Ic77pxOWcDees3qcHq3OTcdS
D92FcePbPFDgNB871rGEwU7Ixk7UBU//aO8hGTpwYiyZy5lQbw9xcVeW8txZfRX/vk2kQukarFTL
a4sF41IeWlqz7FUoCyp6wbCs/MvC5dAlJhpboqaRVfO0XBU3kQljzMdnWUa76LWrugTC5YApqtYE
+s+vcJjPj4k00boU2oGO/F+oHLskLOH/TcVJvBVerxF/dvCO86ibll+ciU5g+bPrL1gCJhPyg2WU
jMcVg4LeT/QMMU8jjfgmWlNVhjUQxryOwe8ZfvCcDZ+5zH+yEon8PI78pMpgHlZt57FGgiVDB1Uj
GrVMIe5/svYIlJsEbLuFbjmCdBnYp4A7IUK9d3iAfqbBuQfLmoW3CirEiSBAxRch82J0rutS+xv/
W1rnJMsQBslGOda5hyqZjegbkdf8R1eh4FR4OKn31rbix0/zJ7hzHWFuhSY7+zhJXdiCq7vzFP7F
93uLURT1oz1DLU/nHdyk47u9C6McXwPeoLEt58oog7qO0pMd5EWjxn66fCc+aDN1Pg3X5KN5Hlwg
U0wdFpCBjZeuvLjJa3wIJeNLCCwGIZlWNOQt/AxDRjJwn4y/9N5WaIEMLEVdGP6y2QTQkoqVBL0/
XrK1DuYWNbpTItfjGzQNhbQNMwI+ZiwkBdJR0g04HZybwrO9TDmMoDhTTacGBIXMW4X4GvoLLWwd
eLsq4X4//O2CiwW3M16aZDcGjau9+B5v7bZydKPGDKht0oSdXq0sC9dUsOv+Jih+NwdLhY2sgDNB
QK8Bv48NJsQmRBnaPbahRrvVhEkVYJgZh9ztpRQE1E8QJACvGTrI8ggNB9KXDgK77cquqF3lClxX
BSyYBPKpf1NN0hr8s6wLuw+DqsHxBp7ljY3z6uC79Gn6x6dfCmcf71js6N4NXX2OC3AdUDWlAEkR
XlaPwGuS806C2E1xZdvc1Mltb/GUUmnD50k5PrNINbHOl+EZT4baxqQJLohylmAb9ZGXL8aqBkjg
19dEahyvSAtxjEyrDSXx+oR7xWKNgnkK+DbrvK4dt6q72PLij6TxcJb2zPYP2HvfFEtA5pK+6Wwj
nSX/XAWy+CFGY3QBzgqyxV07iHgBQPKZVV2xHn7LQtqGipAr4dMeYwcZD1JCI4O+XSTekNyO1KhR
YFkaAMBS/KQPyCYGsRVJzIEeZHWuAU4pd1CjvA4LAxZjhPUx16wk8uBKKRNZwuBvcR40IRImEC+1
h8dZg7QcU3LZCD+rk7w7mGnHllIkQTTfSsaoz56wf9aADkll49UfRYSlIFWTowkf+reGu5K5iJWF
YdJ2kOTAX8HR7Au0J4qVTCsbcB1DDSZsctObapBjQAdInZdzoz8TsAitSi2xON7BFO+i7Mbd7pVA
cbW66qn//CEkzxxRSUtfp7Gt6L/2cdbvqnkFCasbInRZbhm1gZNI07Co30vEl5CbstauKAebCDe0
nULe9qvUW9fGthep9a37kYncvfk1IIFO5F/cam/MnjxtuqzKjF9+PwbfZLVFhbKhLhwSZL6xIIg0
FXgj6ZVKPdXbwxsII3G16bhxx/NjE0dfmdstljof74IuN1B4dE5NCu6Jf2gYktua3Oi6MbrNw47e
P0X9bM7sOqcIluIycIi38qVI5a6BlJLezT1TB//mpHN3sbbOKR/6upgIhhHlL76XBpucBtcjz3eT
eQpjWmFoYTVvcRlR0KA4fjogUubDoPcToN51uYl7nmbTdzbWV46RniHHlDE7J4VpZKW2diiYSvbi
9vnnl2DcbOKeUd5jJYqOmoFMGVcayR8F3eaiY36pH5nR71Xg42OpXA5BMjH96x0Gw8DJK6KqE2AV
0FTMgV2tdoDnqrrUQNFHk34ThLAAzztT/PlZcGrjS6wkSVF3lWTJMU34MNR+BFQWoINfd8xTzj+r
P/TqCMFOAxylQfG1XZH5MoyCYNyA80zH9KvBRBWws9GR2EAPEoN3amXUGgO/aW32xWIOHbDO3nKW
qx+b18hd3Ee2Ncwlw8mMRAHONHQEqnG9ebNxluXq5/TuUp9wBldapIFm4jBL2kQsenC2W4eUOkat
9KocFjWgrAw86uXCbvDnt5x8Pc2S33kIW2pUSZGIpj1Eoub4ddZTu9JNCs/kkhWGlCJOT1spVvaB
6ngJucYHtP8tbEAmD1k85SQ9xJYt4A6yZT6W6Av0JhWCDvtVWRWdtN9av2MYpQb+o0DzQgEOrNeJ
G9AFLlbjOssaGcPRlLZ9iJ+gm886mZBqLIyZkKuMG7gii9YQdsquXYcZd150IrrOpPdGHbB6sLm9
6bh8/TH853iLIQP1qz5I6MRG2m6V9goBsJfBsybYsAMJge0QVL49gx189rybVelc7MNtFGJwqLOO
GQ8C1OwcQ50XofkiG1Me8TMdlbXY7QR44MuQ+sezvBqNwECQS9ecD7AV2aKnwl+fKPMyuh2lEb2r
g+1gGCwj60/kCL4R3LOHtILmpkxxKLHeAX4rxoX6SChhFfyjbc/KRyQ/cmsfMBtF3zumUeH9HvoW
Jq+PFsVHDXh3x8MrLP/nldsoDu09+/nR7BiDI1DWZMaLaXVOjdVprDn8YJDGpxk5TNyMkJvPBLx3
Rzymwh7PGs3wAtt1QKcDSM2wcpq4PhXnkoe9wL3QPAXlMY664lg7D3B+HJdW2vR03NTWVF2HKBuO
fWs1MJkGvcM9nGd0ggNvycNcVpt3NRPW/iy9oFcsfxM3NsTXAVUFRauno2ge5Y3k2J0TnEFjYoTQ
6IIIQ850JDhZGTLISTzZX6uiAKTbudLRROjheOg2rj5aD0QF32UaWBuvhDpNeWM2iWEAi3BDDjIQ
5D3FnkcjJEPfkgJmZMO1A7FYgrNSS0viB/MOLG+dp7skDH73Yqt2GMbwLfgS2iXE2ET9QSLRfWnJ
lte8TSxgU3wFX0gVLuYvHG2QlXa/4Qtmb1w3zqVQjoLKxcMaAXe0XZLCNueP+Lelo3xq123cbZUV
pFuuHSBTgOO6z4dP+rS21MTc52KT4sM3ETH+PT9l/zOvKlwX+TyE3DDFOZspwoh1EMmgptSQaVQJ
x0YnhPKPZEhp8rS9Ovfvu1/kQA6xzGmFUlyD012AQsdSKO2K0T21dNHp6fdybwmTnnuf7HsSVhps
hDezHeqFNnfvRTORnL/AcQ7CKcEDykiQtD9qqVJTpRRcw0CqVf2vJuEJJp5fAJDTq42mS2Ha1ZPc
icA9lG+oBZRqqMaKAu9MjfvHUmUZz/wkiJ3I8Hv5UZ4XnGtoRc5i9YRve/yXLMo/mXwwjL1boX4M
5nmDuFjf2FoB5LbY6iplsfjmslnYjNlH2oO+UiqVw+FSJBcwcxhuLk09l38wQ1sn7lRduNEz4xMe
xSf3RGI/05LlwwOa3gWR2sApCbpp9cObFG4JFUC8prQzv0uDz8CmFUdbRxOKXgZhtfPTL1AV1IqM
ju5RXINEFuIApyZulHRQcKvk1WXX2HzuFt3AYF7HwrTCYmnvJoU+XLZgoCYgABxiFfKiQrixKLiO
hzqxE5rncg5WSnA8R6SIzYeH8sXTxcmWAS0/1B49h2WpA8oDqhjj3JaX65ov26Oxh8ZYS1b2jgGL
mteX5+knK1SXKgYtTzOiAydu+R0Dq9Jb4ICkfYBJMQ2FhNfSWkGXtnuEf+CdRpDQulI1zHkK4xVF
CnOTcu12vh9vO8mHlfFtYEhyAvuqM5Xt97UgkeofD5cto4MiSPdoMhftMw2i8QshwfOicRVT9lJa
KUHZOdY59MQ31XqwKX0TMGoJuBII5LNHcHTt9PpAzJnxwWITQOTrRhDUkVeyyyPXZYFBjLuARbu1
0k6P9Bsyf5/xJyF5ZRymybNCEGRK4wME+7GozxvEq4bU2n7oi1e3qDKtmGuvsPoBRMJjxndmaYPR
WM9GMPkGaEhpbKXm8cMwj35qRxptCSwo8g/elcMypjAwqnwgQRWMMrXegpkbzsDDHIgva2aAENdp
+Nblb20ljbQR9l80zN+MSu+g4AD6YGzI7Kn6yiqPC2O1z2kfC16N8woMqyj2lFeyQxe2x1LtysTp
KfHZu4zBKsDZw3PKD/WHk8Gi3xznsccVuM4EzKSH9W0qbGYx7j0Ff12nebAhJi2LayVW//D3udoP
lMod3OHfjTnvMlNl5jYVqUiTCwHS6SygMQdlf4rwdaum4eraTxSHttaFzx7omc4aBAT5I/UmwO9u
AfrsX58bmeNDSuVkSN+Q4L2JU3XYB7a5lE9qoj8utA6872PO+stwtUJoX08JpHAiU8wnqjzLLiPr
CcF5We39Pru7hRldHwMkA5UvYbouh9aEAP7yrQpjlLBAyJKeIrmuv1FwDi5Dcy7ge0tKeoJIH4Vx
S8UafKRcMmxOMS6vKFIWx8CG9CiwKOEr4ExvjxdEBIreZcAcujMVdHsuhaBoI4HIhdV/DDhxzSaH
LjT54rBMIOA9Z3agkxGPiS7lgMzriklYgELoc+WqATxAm0fIvptwiY9rXNkt1qtK6WNEMq+vZQNt
B9IYcQtMuW2GuDpFYN5yYen57AkRozXurBYbH6YFV2Kby417nLItlEP0NB8pxZ11LOBy1OCnehr9
Pk9kEfB7kbuBfpdBQnEck8f+1omGuNfbotMe8+VGv/jlupC3XGJpeoTzISsp/XOhiIUSgWtq+iY0
cWZQYO7H8ksF6TNw6x0bhFBL2kVnnJ8svB17leFNSASXwhOjX9eGFx+m7J3E6HvbqH9PksavqfbV
E+cZT2Qt7m18ecUSxcsRQAF8hj25wHiAUC6t/5Hlbiagi15WllIBXcHq8owgSkoVB+Cd05dK+JHg
Wt9VROK7LpcfANKgY+pI0WpPEXSmcRCI27L+aepnVOGr4eA9RKLmknZhVlXlAyE2Lk2LWmXLyZ+9
bjm+VnutjVf3ENo+ZHmLFRFZE5S2Y5eMWYnco62cZ8AhqpZsVO1eG2PC+aXVn7FEn1MMkqxX8/VZ
4cVN2rQCEm6m1HVt/GxTsf/l+oXE20dh8X4XD7b6vzDM4W7sDxiE8DIeQgjQl+eCAUB8XMfjT6IF
kjKjO8t5J7ePTr15/RQA4Jt7V9FmMUXVvOsxBy5coLqrqUjITtRE5aAEP6GVYXcaDPFfMGHo+mNf
/vIFiluzeWaGoHB734DjYnwnVPGTSRUbi7I9Y/5A8gH8697GM6zc88sOaAFkAnM+ifuiGJqViybJ
xXD+DTk4jOP8ttYPMpIzgPsFwMch5UznQnAUz0cFbAho7VY36SvK2NNFv2yatNb7wsKTZL7TXSgQ
rxJxqBCuvdSB7GU5wt6CTJK2KlCzSo2qzj1lYQSEuEc8n13OGr2+NBFIsFxSCe9sUlF+yAtIvt7u
LrmMbPBpGBbzOqLnaaby3RpFJs/haQnJnOEdsLhduCg/SwhpCAfpZ/MJzYIA3zEZ9QyC9Nw5GPLI
wOE8p6vJuFZI+1rxhNuPsTW8k+yS+utbxQ3WGLEMA0weh94CliC3vA7uk3VD8016vd5Pui6rY6/N
vsxeQpUeiEAMxLJt+qYLNhRHUlZ9d4myls9KL3uHtF1rfp5Nl1l8mlarvaDIN4aQxBlmfA5Q20hU
dq4XvsnDMUIwA6lRp8Ml3KdftwJuECy5DcrWVyVxdba8QUxW2Qx9bAYkHuLmJIV5d4yZEHe30H41
n/pd/Z1+m9iCwXuMklpt7oRXC2L65z23e1Y5/s+++/8DQwxfBOccaGx1rxTJegIyzoxo4DFAcqyN
V6v09pRK9KfjPDlAfb5Gb8+VVUx1l4iTToMEd+INjUWgBQYckj0dygeo2998tAJp2beS0hWFtNHP
YN8YFiydRVsGt4E7XhuLVs0KuT0d3213gQBYyl6BPafHed+SgLUdUWLXut/0Al3sb+bX6Iu+Zl6b
u1YMx4aoc51yKgWJl8tNPD3Yg3nOLh9CE+mJJGmqRfJon83Yx8Ym+BllpdqjRCSvx1vQRY4ut5lc
FC46h2qh9Figmk7CsotHraXmT3kMyXGOgXGzeuQoNsaTf3tkXUwxSjSAPbEEHuWm5UYN9uwSMjTT
wJQ7LVw4hpTnhLibTuBv7CADzi66EilqCf00WzuhxaUTjfnGkH3Si45bmxM1wKmwPjOR2yIVTB4+
KxGVD1fENlkiUwMr3BgQ48GvhHyzZ4iiYp3vypDPhpmxRdMhga3Gfk7hupIdxMQv6VKoBppKgWl4
oVO1jtA3+EBCdSzkfQUVCTXVqg1lUSf8DnzojOmXoYXBb6oo0Y/cgLYbl6OjdNuG2S/vlpFkjdby
Dbjha8OPnGGPE/qN+tnvnzeHtlqDYDQEC2XijLQgl4znljjIKgZYKYfjn9izBLRwkVh8LxDG7q+0
tcPWBkZJZVPqLWK1O8OaQJ2E0cL2yDfWRyACoRhZlXWmQo0muJRorAC3eLj/ozRTWxbTlDEqWMSm
9tnuclXidUkDVrI42TeORfTjBxqBSRucUrUKNrOUPfFBZ8+TNxMTIxq1B5hOhUU/CYNB3yCjmPgy
tWrRHXWS2Bc8m5fag+jW8Ubu/QcH3am745Y/xWwAhi4JTNr+lT+76hDTgViVnSEtoOdwtJjVe+Qj
IYFHpWFhZVFH3CA0h4gA9Fza6t1u22HjZsSY8wlShiHxDrZwS6aEMFVe4iE0ORNxq/Y5neNdE5Oh
7IU3kB3b4t8a0fzQTKDujRhyC+DRdk0DiANIEQVuTkNX7SAzJGqvB3kBJDpyizLgfF5D/zKEWLwl
flZx17xNrMORcaLsagG32YUbVKFYWqEHaX6xR5TQR7w0tibJDhYY/URss+SQJopSj0zAiIXjsGZ7
j/HQgTxgM18NIduYFUdGiGPTEAZ8n1m7sQktHA+vNkAtEC3pEtz+DjQjkB6SKOdbRN+UjYxCn+im
W+tydqbvW7/nMfJhL+YT/ET45k7QVYpgn5C5acmFpSWvqg+h7gXHg1IweM7/y7b8lgmNjqANVEOi
I2VaLBeKG/2Kal7HmeQDrkjMyZg/hRLj3+7z9rBuM8mIYlC9sU+sC5gEbrNoWB/ODt0GVlY1QrHc
+5NAP17YwWRAD2+YPLKHnvnXnw31s4OwdL0ii+rUoisnHhT6Ofn40/eaHaaEGXHpbC+KalxwwqyD
hY0yoFNoZpubUxyaa0GKD1+dEEc2hzesz8iBCapvNzc+x09n2DoHDLuLhg5pZwmIXfpi6jxG2oNX
1QpE1b/j/MvisqpQDaiK8PAk/5meNHgYN0BIDFh6OFCyLtlXNRUr1rSm+YHaoQ5GnOfeZl9CkcCd
L+5P9Dx7dbQhhfuqbWyjLIiPb5Kj3JViNAnKv2JlV/J4LcFVo+R4soPBBdYs4TzgJwwdjbSqlU+P
xxHT1c79Us2aKyzcg+XebaCuwQrGP1CAeY9kZoL9MWG0x8H0cVrb7lf8NgrcMr39dnMVZudq2rKM
AF7Ijc78jd+lhUecVbByoy4r2ByG9RnWG7H2cpoUfff9j8NoQckiSwqZjMoD82HXp08+pacszQvm
mfcVgfiS7ZjITpot2Bu17NRazEBM62PZVHbBCMr3VYIeLSu7IpkmWs671nyaycwG+1eZIC3UR96w
ypJSpg/8viZugKDPwMp5v6RtrHaLqsoAxtnlfIzakKP60rNksywMPA70lWS4LLJgUzVWcPDAUTiz
w/7ahKyFW1olowFVjICsC/Ol10Kv5ZrJWNefmw7VOQWZQ3yN8l/s2rpfA0o3N4G0n2ou8cTP1q3V
Jn2hQ+Cr5K2y1yk0qw+BzDgmmK0acoxrkCLKAb7juH1j+gNVeh0IJsO3gVxLFycy8I0adfTun7tz
tkpcS+AwWnrHUhHm4An4iPVjW/NRTvfZSdYQ62k2RizoaGzFNM1V5YcWvtT48s+DNYZ8LavlZoLA
CnztAek7kr6frCDyX2DY3hzX9EGEPqiD5aS6NPDPS3j1nzFFWiIz/B9Bd31X0r1RcynOg/GXD9Gn
5tFNnvCf76Swi64HHi5h7TsDhtuu0ksD6FSeNSYlFBFcE1CnE9bV7ErPaSopShLejNMK6RBq0CuA
AtD4d6asH+XMW7lTUraLlZFa5HYbw+2vXzl/jErgwtmlpHHhuITy09EqcgVl5LpYgBygqamqANRA
Khj4fsXxsPjaToiw4k7VWcWcotG4/AfqWjyCnIqhVM6T3wGNNjdX/3sTKELpm8gSAFoQS/8VjGNb
2bdImwTm+JwJL4FCfJj2giUWrCtDZp2Ixu3m/yWuivSJOcGLOr8N3+TZ7zU/bQXt2CL5bFdBaA1/
EW33KmC9sIqudbwEzAjOWe9Ux5Doag/yQc7LEIXsqiHVeWb6aRps2/Uka1tB833lxN6307Kr8tvd
+Cx3nrBG8In+OLfm9zp9eHwzqL87mKC6BOI33KrOTiZpjtgvx0C06cFzFZG7TMhYkqF5P33Dlrpn
LsMhvvCf7l9RIyS0Cira0lwRhSxmGb72US9jAOB/TKP6hvIF9uQ5bUBPUybbjefqlE1UoME2QOtV
V66DaQgjfk82wi5G8+hCg7TaxYUN21YJRjmtXLHprJ6LBRZUGOzE/hIkumUzm+yI8/67XNYGsWF7
A8rHxJE86ZNKId/vQ84G8AS/YlxKEYvszMGo+OTDan+yPEzFYmT7If3PqgB3/VGAa7iQDLaAGIhj
fOI6ol97LGOvglNxwf8Dw39q0jKgMtsVPYkKywZlWlRzjDI7QEQeLhlXc+b+1kNrPmk0XqAWbjRz
oOa+MeibO7mUFLzYgq9SRvjmls9fNTSUvGDXXq6g1nSK7JjaZIw492OLtF1LKfkyqZcdjmlHQRem
KroZOXiQCUw3E3ao/nNtrzMnNoDZ6pldzw/yc+ju9nt5/7H83YWh24n6EwpvDpu5xRnP15f77Ti1
qgHOrqrF4CKYmRux43Vask3g8g+vhAs5X/h+wZNzEGhtxmoUfxHvrnEVoR8/ufyrDkrsuFCxVMWA
uu+43Ty8psiwvOhUigiEAKLUWP/wEUhBz/7mCSe4zSaNDghZfc/5S8BTBnUu4gcU90Hwl/Eqqfnl
dPBGHQCkSoBFsAn9czy0Ad/Vq5P2HjvBT6k4Kj6x/vVOecZXNurrgl9YlJY2oZ6pKajbwJhUvgir
nPRjLGPbsErmPljaYLUhTlMzKMd4x1mdsghjCa4R5fPO061GK3R5ADjcspRpThsWe8TBHywodSwR
xyg49vr7uWkK21BFleDsORX3Oo5clQo971/yRlYx2/sNvAJLaiF1xsiiv+ndAWQcUx6aEBGuwko2
voBukR6OWUAaGIMU/Pt35x4l1+9E/0dp7v5k/uswKqGFx3bM0E+fAD8Esny4y4C8xTe/fGXRNPmx
fbXf1QBj294EfOi1SEQiyHdJ/a6rXv2E4iQU5DML4mRHQt6gbUyPf2xfZ/08WGfyYI48xH3raImg
FelVuAzrTh7Zsyq7BDqOPMjMSW21zboAF2TXCnFEr5Ksppt/SQx69xYJ/3DHXtDfyh7lyI1qJLLJ
3nGfH5VTwYze378AGpzwgNipgc4kjBCxzPsxgPkacEGm/zX80KmmsAnzydCz7oldRxS3hS6E/Duy
7SS1evtyxtGbQSWiHQQ2iID4QWFDGTvOX5XL5uSeNtR7btJXcpPoIc9yIQ1kRVsyj+E2QruuzP5I
XJyd35kSp3Aa2XA6pANbZInrroHA2ikbUTH7PpLr03DWLFaUrcuLpOtQAEtZ/92TdDx4azd/gmw4
cwS7IkFQBt1YS46zTDh7cCoVUXxF7cyBTVyKtuZiPcxxQ5F37O54Br6ceyBGhGcypPpzrv1x7Si4
R2KYQm3nEhC5PCVT9vOGQ8HCe0QaH46zYz33QZ8QB4OXj8GvLl9Fvap6hjVSCdmSYr9G/Lk0bNbK
xZKomb87i8VniD/tE/e3E2Xv2G45AXX5XG56idAY+P8Z+4gmXeLCNu2UGWseIskdlw4/W8ZSw4P9
+2c44MFORiAKSXrI817OLrpk+RgjzezU+r6UM32D4xkHNVGNIfz81QHZJ+9hlgYf/LckQ+shuylc
N4fprpbKk2Grx0iF6GCu5k6+aKBQhp6fY4IQglfTlDeYKrNGkgCGnuDkbIqXnbtfbPxe/chSuibQ
PAq/fV5aX4ZzkIdC5Oo0vFlu++zkZiY1K+Zx0iutb1lWshMFRc2f9FRvhIjgb40IRw2ckR/gAFco
LgiJ61Cd2BJqQov8P0SOXNz5u0mqBvLHzZYd/ma1ZMa4A1y2Df7tpZmqj6mkaOTRAfzykRQpc573
YwKLLWhkKvWTb60FE1jSKEbIIPnSQ6PzVz1ac55HOl4HWLbGaHn58zl2YLWh1ZcNTiljdXIRgkY0
c38BS3e0jA16JtoBOL36CtYuLre+Gowia9sQn/fiP0WWKIirPCu6bsj8cJhzvbV1XwEI3jjyhEWY
Ldk7cbbqQ23qtdrZKrFVDcYw7QrJi2EID/fENdiVDZIYxoFMU1YFZwbw77PdYvdoVWVzo3ST6opE
NRoCmmaHS7wBK14dFFt/wfn/iSP2/vPD1siT5MrZh+tsF3EueTRz+RVu0uMmG51xkqzywwO3ySOS
7B/KJHiwhfcRvmueYDt5z6ak/odbJ0ZqniY/t/pi+EJN6hc8SR3qRvOvuR5hShUQV6YJCAxCHhmb
nAMG6Lz9P3/U5YP9NPDLKReOoDEW4BN8rAoEYTFroVUX3+dxDlgfWXsphooXkT2Rblicc7UYxgcz
IlCWKK+GI0dqbweLCFTH9/X+C+5yWEFUn4b8C25x3f7+c6H63LSevppwh0HxAkXteWnWuG3+IrRs
gfnXhQqMoPQjRzoV5Pp/tNBNiXoq/gWCQRUBZoJrvrXppOVjHjaGKhAd9S/Hry60bRlBIY3ZHexj
aNYlHvxYCQ/7LAiwWvWEE7nQWsXHZGmzGPUxHTZAyLln3E7e7BrlQpvNVMXh61TzMT4qmX5OiF2Q
FcLx1nheEa+mZQwffUrAmrdMRu9iuK/E1M0+RC2ZHVBJhT00knqD5u4LpKPnbaxkQges1h0HRLz/
dTe1PS8iJdOXlY2pRt0AAcQ4sJqJX31PUd3XwPSmdxmHsCTmOoiVFIpIGA2iNV3an59kHeeoF59r
0bKYuu8GECwfm7N5tAo4qNUOrWVwBgZKpteMxTyW/Au7ojCMcdafBfU5FZGq2AvyVRAqQwl5nB4l
L/aZqib60DgECxY2V995MTp9XisrYcVisFu202L6rrMkw5dX//aNa7s5x/Sg2McZcKXjomtuWRAN
3PZKrFsWzpzT4VMysmFqC6EMYoxlTj8cPqSWnlT5TK20LKMm+Foxide8VtLUPLCc6wEslx6PDDPt
4pA7djRFdyZ1wb+dDAqnwel7SJGSE7x4IJbRNVNbRkrGtFpo8pi+8Qc/PgSZXTWJff5qk++cpmZ3
lbqbB/cGQIUlIBBeCuwK5363ILQ7dYbUGiJ8saS6KDooXPsiS5Dd33tsK0vwpipG6tX+lC+O6BCL
L/b2+Jl04IIU5fmJ4LaUly4CwJPTPRAAGwqBpKKsvSuijwtQZ6F1XHcCAw7fIQ9FPkflIb9XPsVE
HxMEaJ4FmsXeffan+UJ5+wOQLSOcWKj8wkswT24AJgcxcIph/V2EpAHZcGKn2E4PoeQEyul6/tZj
Ji304Jirt8QHc0OOEbF9KcSMQtuPIyJv09yjUPJZKjbCC7A6gL9J5nmop9I1t0K0ne65/XQoB4AV
/GCyA/DbqzimeYIyh2qROa+kqttI1E+w0pB5hOa9oosl2A9VZQ3bz/rwnb8c5fYHiGvm/uyr6Ui+
kk8oNyKfRqUhL3xrLidwqt8hFH9wgdeomm/1cfECxLg1RZQEx63CewxPrKF3FjyxIWl3NDBuPjbL
qYF8xlxdtbGKbOMkjIv75riOqZFljzEVEaH+Qg91OD8mnFcKIE9/fXHAN5NxjL3hgMVOo3LhBDaH
51pVreOliSlIoiRqOPJ3Mgom8/WxNiw4P2R+V8wJ61mt6sZYbN3PGvQa/E+ohiFfcwaaov/jmnUL
O+mJdhXMn3vJN6WMRQWcU60wlX4Vs5JtGDy9E6LWAYcrdvannbIXzK1P0Cc26zYNyvEsMydvXWi1
bLuQHLeaGbSbGE+ykrdCpicJPdkrauTn0/61K4+G8efZhPgWgI220s9jYqgePWDxJjqQI1F2Kh/y
oyo/IYXRa/8bUOfONDUFANsT3TOtGvFhPPfre9mrYvsaH4TQ89fXJPUifVdNeJtrsB5me97Nv8wa
oblnxbfHjgIiwVrjED7Wk6QNhls18dI8dPeM29AOcbdcs0neHEXVWjMQu95EZvVYdjtp3KnFvj7J
tn+v73dEKHKH4iTdeaoq/8N3tJbEwBoNhB2iORHAU6mwQ1Y4J1bbvqlaZDXLCn6RxRE9mzDWYRHm
t3rGRTPko+HxGYLk8u/LnKElunSyx4gqaGCjlb//FIX2trnBLp5xNHmc/+h24KYqN4Er/mZeCVcc
J480V8uNLJH+30IUw5QKDA98nC+KE8TiBNOOHkO0DvGWTT8/K5C5+Mg7L5fLau+cdJKNI2AojUw5
dIDdbbUC94uNX9gsVkz0NBPeoiaI9Dt91hgoEfLemeyFveKjQbiYznscXVnqsFsP3ptIoRSpWHI+
TZ6pVaVgwcUw5l3f64ne7H1WPNhKkEVlbSUp+YEEhPDxy8phkTbrFib1o55MzRt3uJiuKWrRAnLj
zXiWp6UJDVeQjUmIFvX5jA25pytxwA8L1xSGVgRcGh8apN9nIHkqDtDjinQdQLbIKT4NnkWTP/N/
pKTm/2guKBftE1sgANFADrkrS6jGJV1jb8fzmWktFzaxHZGFId7MTPAmIUQ/k1zHI+cB8cl65fsC
f/i+fbfOqlO6z7I+jfkraQLc6n3+F3henOtT400G3YR2OZLN66/hr/wuJuW5bLsBVlI0z9urrTQY
UzkR1tnYT0vOBtLuktUW7mIwdCB3DfZYSCYKmDNSFZ0YGeB9pXO970tKBrswDIWTc4aiEIB6GAzr
FR50x4R1ItMftTS3tV2t1mGMe2ZEPNMg0fI4Rz/SdIudMgIKwTQzFDQU1vGwnPHPdqb7pzr6ZNs0
EhpwG/5X2Xp99lthlaL42PYvXkDxqGuEyfedXYa6ambnqM++oRg8qeFulQL7Da6e7areexrwKYnG
axSVLAmvgN9Igdtq8PF9DQRJ5P11Vp/Ts2DgJj9GRHd2EhFIsglUO5JkZLI8xR9zyYRULAbIJJNp
OI2ds3/PFMWdqj2zcyCfLtru6XWKjVN6VKyzFdDmtGGIXXtaEVfZehDJF46LsAr/R7vnUOKrgMRD
tU9lv+lefWw6ghdECLP03jljmaheZXjLVh/RyIeniqSavcxnoNNPp0z62BywNCAm5m8b9GYOhqoE
QXF57d3/QlsQ70w+6KLB9Kbtw7L/+V+PsZAZs0ZgIE9NdOufLkOVoK2kiKzRcuK6/CGhu/QySceV
U1uvlP+CfeLyncpTzrHTBeD3JqnctKd3rc2XsI99yC4fYysKTAplHdQpSIIbr2sTH+HEyVUhO46A
sE6rtwrxTHWPT2WjgO8kM2/xbspKtFjWiHAlAUd7PEoOA1tKrSf+pI3RFq8pKFUGm0/efpUV00vz
4psm+cBkxqBSDorC2wChxBuVZ44jbGVuuMANy3FWrTLQu2Wjtdp+2tEhGcwvc/eZJxFtB9PtxBvz
iDyXzh8HNzfqyBEOyJRS45x9sYcOftw4wpdhSRDJXjFyEXNsOXjTulVLaCJBRHmrhJWFYKuurpd9
zJEQhKHxfjSSgRIk3MhrI5/ovED/7gWZLc8ecYh9iGgr8k7FbFxMEFB9+8teLsgWvgcA4qK89NA5
nnpLjLhJLnQMMd7usIstuddOXp+1R2U72lqFJCrXmbcIycfD+YZOpjIoNeD4Wp3cSdfLgxQW6ab5
eP4pjH4MAYgrVu2bCHtvxd7g9Y3B4I5WGGIJ2lt/y8SkO3qBNc2l2zjhY1iH4oeHLIkJ7Tt9N9Jk
oPmgWxZAWQ1WcJho7XdWgqm/2Yky5kmXX6XHvGudrU+aMjYicMpjcLrbv1rXyCISDfKKJdcaYkrz
R7SKvJxI44hgqsUBplIvIFEkSlRAhsBMVmf8IfOKvc5e+7b++eKo4bMFci/SUU2Y9GBy8wHrotYu
c20QuJRTRGXfv/vMJnZS/aydm+1RxFNeG3u95cr3LiOtwLh6BLr01UNd4W36htc1vR6o/6tJSGtO
WT+t8lW69ElGFsVc8VRkEzOnql4SLXIaAr+MZfcOXlkR6Vys3XZAT7aeXgBu0Ek0DPhhBo9LyT7q
2BR0fN16hVWTbG5Kjxkft3E3zNVYnNO/BohhiTt1SuqN5WZk8tB95vo1hdtcEpkqF9xguRTTu5VV
ypWhc8HVwqN39Fqwko67K184SrooAUW/aB9wtadj/DuTC+qbguHJRi0b2nNm5haMEicgu2KvcK1H
Hkc1GF8EN9M+oxQQhRts/6YvKLmWRokEnyxkM2vv1fDceWfegS1GA7TX1Kp/MTauW7BNRZi/jTrp
Mr+LDLSwA0U6dehMSfKCQueH4lGlCg9J6qyVgKDiL+BHNH6WFL/G/EkZWZ1OoExSMCZa0Fhp3np6
EigNW+TNS1TVSwhSeFD4g9a7VEO492XLWgpjjq1GBbzySk8BpTBwquVZ9LH2U92TPLFcJ7gMHO04
S3lUu5KWzf5QD5KwnotKnp818CqiwEDKi0wB2k8o5kkGg266yoQQs5kIB88j6LcHjOV9bUNLfk+N
Xpuy2gH4Cp1Uc+ntbxGoRq2y7Kzz6LdGAeCW5gz2nLp7eUVi++5ta8CBXX7hzgBOo98mKKac4Wrk
bs8BZrWquLr65HHWIf4X7e3gS92Mc1mtVb8iq7hw9OOMUf77Qd2tGh3GhR9Q1REOhvp0LsyjRjBx
kM0drivxcGix7EMnIP18pue/TxGM3oo7DXGO/Oz58OAurm5LHmyvUNDTXdkkLhx0+Ru7fawhvuTU
VsJq8QK/PPumHZVCjor7S++QbR2dt6u8F2GtLnYdgFILHx5eHHLp+EJEoAigYHU75nzAkuXCE/O1
/sCwnQhHLJLYN0NohaLIbDCnrPefnEcCHEw726TTrcSgSLr86plB33tZxqhcdCb/EbU7C2K9xZ/A
sruxuMSiARxrWc3viFYDeimZHz4y5qC2yMbVscx9FGtRAzGyoGDT/7BphO/Lu6VLfg/jOAFlkWRO
kqwvuW56Npk7/yPdCUs7eRqc/nPMZCGMKhpjerHHyb4lC4Lu4HzERaIWWExx/h4gCAcHvdeEXQEL
upMa8+vgUqg/qpWRdJdARVFrVQoQ2pk0aqr8TMKG0sEM+1b0SJxSASvSQA2JeRNeYqjzxOhvCPV8
ilUkbva62M848nIj2w6OMllrbwc6m2Zw/YBKxcEhSpFSu94lm7i+SiMmaRqTXwI6z2FKVLczmt0a
lHdwYzIV34Hi3OMuRTrPx4AdzHTr/3H8MK1QUiT/56KckCx6jbVtPQIfZPoFLFffK9g3pWhcKuZG
X2WrYOB0LpvdXc1E0RC0NyMbxLOmVxfNr2SimBMzzX0JUNJEGFcawUTIdsRUkW0BE/l3QjYmELj0
EjPy9JRFRqXihC7sFEWdbzMj2rWXRaDxszup5665Sa7TS5N3Tl2mUB37LT/aiEq0LaWvmxThgX6a
HIujbVbcigOzW26CDMTlajwUIcR6u+3Phhex+LHEMahb/OwmXZUymn4PfmDlJzQA0+L/E64IiN1X
HGKmVappO//89vkTh6j9EYxEdUHc5WSdl7Nns96+UFzu687K1UO7kdIszFBpGs66VGBCaK723kDX
F2KJQBxbjLZYmF0vTgL7gT50vgDuvfHuv1FgNuQfKYZlTltYUo+6iLTi8mOmN0+JJvoCFLiXztRA
bTgdegrPsW8Oz74vqypP+Quyw8zM7VDGHRYxTvMAAIte1ieQfaDU0sepjHV35TovCmiL/XGUMzLC
DCHZu2CF05LXfWrvDGk6zCQTjOc0/kyNWaRickb/orRmQ8uXar83aZPcA9jrcj5B/JH/Gkfh84jD
iTk9FEloqWrXpslGWoHN+VBlMgZgewdvplhGOI5yVO1M7nSHFMzz0HXkgjTZxxt+hyTkyLGRDSfN
PVB0XNjDqYuenD+ftJz+Pm3dlVRkC/DufsHUT1P38sZkMDV6Oquz5fWV+/do8pD+f0t9ZWEflGqK
2+D/o9iwhjP4ANApcVeTgAy8A0roLNRDw9umFjvyXLJQvhtMpg+3nVY8ifmzp8V2Tfn+uRJJh7XV
7o9pQV/anDNyCKNB1co+yZPVmrcBRKL+wKixZ8gUoM91NVvZzyzFSyp5Zs194aPXjjB5XCFcUahq
Qpj9WRmTfhDPQQEod4u8oYI0gPBFElPZuwMdCD5xydtc6abiWtjskbdG0qVB35HjussVFPRCgVtq
lxvPsjiLVMxecj5yPOAvPCH9lUKeKs51VtfmCSmsmHvOKoEMBj1Cgyjl/hTXdY4L68pOYvI3X4O3
73a4gZIpVSwKYhxtPrC864RDV9i4lc7qBicXz53YLG2jYWfGiMPxC5j93CChQuGZd2QnbIkdj/zm
aaNtHdOmr4PQdTQVgAeisFtdDF3R5K/qYhnRi6aO4NmLB8aEPpL9/9IAdSBUidZJvGpXFLik3Tdb
yOT467WrO9EsFtu5psJPAhXh8+HrgmXoADqjagXJ6LintdjmCfO3iERCyfFCzAQE5HHgUOQ6/9Rl
JzHIla9xxEsT9VVv5O8mjjIvtV5gePMm7vW15b36bgFtoFw6yPgLwlotYIwr8WLc6Ek0BhEFPvvh
wanPg8qCF1Tr7W9R+48flkZ4Jmm2wnvRmpE+3mS1IP5tLAnsmdUJ0RLugXR7DDYWTLkUsLwsHJrz
nzSYaURQ3THdh/n8IC88uFDMukEfuj1xE2g0tbzhAY5Wim9TZxfKGhwkCXY0M8hJo7HpC3DguMh7
9P0yov5Cj/2ldgnS81AmzL2kd3bkoJIc6muJSplI5tXbNP2/nG4fqe1ZSNoi8q8sk3VJPelOVyPY
E4gJGIKlfnZN5NvWunr1YckPNMnNVg3tihHXd06kx5/P6uevUusevLQQVWvJoMFGAGdTL4j8cQF+
8WSzp6uIBdZVlwR1jrsmE4wpg5GfzQ8X/EXJxx9JH36ci0KF7G+8Ss779me6BH8M+S+DI3boquaJ
GJI7xHfL//xsWzW7otVcpK4ZJcs5pX5WmEgtLabgWF3QsS6CUUZIo0qd45FtvXGI/lu7kx+tSRXE
cn+WkefK711IX1iOEq4m3ti2qhcetmpi8T65M++evJWvAT5yW/evK/1k7TPr6BUmmeUNWfmvZK1O
h2fKCSNpLLu3fn3qodHLLtTEwHS73D/kIw3LCDVnnPwEQmUfg3q6CNc5OMsVJbyjLacbQXOFM1N/
nTQoVGktsOs8Mt0ZfCiuA5NtLMgV2MJ3Y8Fu1+TADpbGF5LFo9DCdXEGLxE97JqzyeSnHlcU7SDU
jdIm1kFMsN6HSF28EOVamvFWespSlqWIV728ksyszw8ALaWv8yDZc3AlXkiBJ9zVvDJiCNo4myNL
ybgRiyQP3cGXj5SJi0CPjLfHWW/G96ip4ERYxzvYqPvTsLJp2iXpHPzKluvlGJ3Wrb7qNt/+wKcY
KqWHPsWe7hkHfdHu9xLuxFY9RIx6S0KdTwQXng8wnxyQsVPfJ+VAQJYFH/H4y3kbHwtwXUT8Lcmx
gZbd4LSiBYLbgSWCazuTbYRxDzRYAiMKj2kQNQPWY/jdQrW5YpEyVichgaKWvYOZ/bnWY0NpaDIi
Jfxokhe50IkoAhsHRB9oEp2qfupTfoEwqqT3qTT+hRy4awpOATIMW9qSRn2k+E3eFw23fg0RJpXZ
3bL1grE2tLLXvNQL0kpkr0xg4aJuROOYgCwP+o8R5Cu8MBaws18c6roFgliTttcK9nEb/D3aWVZF
CwfEnDaIVThuRNc73vWEPcf9pc8UFsfhbprUE7lGddqq5XA5sDsfFKcl6HSiMg3v4AHf2OHw9Y+r
PYojAQwlQ2XVpeGbpPmozxTctuha8hjX1nG0wiVgX+z2bhilqgtfqwCndw1Yb8gBv+Esb8yisyKe
FpbeIz12CvBK3AVDzOICAOydvh4iJrksHazzxk8oHg19PCSc4XAF2N9XoG13KW+7XV8s7zJpERgV
e71QcWL5HxYbgfVI4x2Ssgjks82aVQk7LO2IQXAgamJtihw6fDjr8Flr9P2vS7GTMoCrche+Revl
f9rFc0xm9kmxqpyY5/sng2ROp/mwIpH6/qDXkY31W4tvQ+hqLPL+FNJx7fZT0Qg4P7xPJjoIzhjz
XNXvf0FGWRXX3Pu82QQUGc5UsEji+C4Mj2x3l9ou6M9jDAttQGfdnVL4ClZEVBy3iI6dXBV8wNZR
K9JqvJzQwoY2yJ8Ciewk88zfEs6CufZEZGfi0BMFT2lY21N9RtQHhd4SW+dGwxRh0WSbC3M9w+g8
lzEa9JGUm5wJuyoi+xDNI+M5W0ahKZBD1G/VtT4M9WuLt2lgxszLP02Mc7dH1ECYOWdfyg5lJf57
0AVMpuyexyTTuGz8rcsfW78g5DenE6h/dEM4wewuOAlPmhBKfU0fepcOHTtzl8H7fdMgrbor/GcV
H+lnXEyNTUK+02R0KCw4z89zsAhfPoehPyZylzy92rra2kEPMKppc//KOabNtNomMyr+gpIQvGqb
oMmo6SZywnpwXXc3LU8ncPQCxGpfgfWOCVcQdJoo0wTRjViudY0M1wmDUkysYFumrJ/6habnFewt
3XKX5D3I1eCDp1z8Nr3hlsMPqdZKNkfCrCqkVuOa/DSDSpixYIEXcQmH1f9E2n4ONzdwJASuvCnF
GZMv85pzhh1/ADb3ZpOp03+ssM9Tn/h49b/o+Laq33fJN/mmlw1Xrad/biH/LhZydPMd+u2F/GdR
xz/Td4uqSKJpbNtjJ1uTzqLOzO7Zdu4YnLHkO3aHS3PsaogB0asjGUzuD1AoCidEDpcHCOhx4LoU
6OtYFqQ86PJexp/FOah7UhoLsgmKTvDrsLxNG/nwa6b54efuJiRLoZP5SrqEmienYkxxZIPLedKV
vP+GFHB+5lTq7ncXYfS9Oofjt2uaClazoV72OCQgEingJaSmadbMTLB0gFVaufbEZ64ak4x2lRIk
O3xELDsj1jlS6I76xRXyjhEBSqXTLAgxCBXJjqR94v3/fB3TnraEG0nx3SAl69UGoFjVl5KYvgY3
T7wtR8HjBwag4MDvYqGMqJFMLmrVA4OphKgeib+iaHQKdp+E5RU/n8x/D//GOy0hV2yzJG7J2ADy
EBMSn/C9x4XXZtIGgcd4FTbcnmV7tTJWnigXWSPEp1wNxWdKzWsTx7gHlp4JFqFLvkbaQgsGHQ55
WhAOCcA1QnDrh5PuD+GAEO+Onom2VVjp21jL+2N7k9YyyRFyAbvTnV/0eb8Zwp7Jr6pGjA7ZjGdt
JEcFtimYHFk9gkmrDh5r1vZXwSQB1HcBniTkqu8mpICxVnZOWlJoXDfHSivEA3GEEdqnKf3htm72
7Y5HAlo9aIU/xXnZFWa/HciNdh5ENB6pQ+QSwfoUwLvY1XCd7OTqGcpP7uFSI+CeIISs99w4GU2F
fW35twjCvhtM3wKqU8yu2MCVkwapaU6yrNJSpDXA3E1lYLtt2Cjwutp9LSsQOpTNBt7Yx6vzMuHW
98wFgJRJVznyXfPcyIixCZlDYYCUNWvRSnqARGJYmK3ZaHhTnNwPO9wAuciSkpTgwZCzSCYZCibr
Qn0+ZT3LcvsNjTrlYpBQczf9y5OQFd3kIz1gM5Pwzu5AoXFu6D74bu9kqGcOajwUnSKO1IEPqhy+
R3mWLNJ7PQg1gI3daHlAPhwu5uM74J1OSbfPEWUACLYGViKW6awEdImhy2FB+WgPcDT2UquojRNx
DwHeF6NSEB4XUWdOjiROGdhm7pXNIsnY9W903+xjzPc1ADs0a1J2G4Q1FUPaQTzZ8iKbh6eP3Voz
SpajBXG7/Ve4VEw8Ny1vcdc586IL75qB+wVS0b4eKESGXW5Cj1TWBEN9fxzfP3uzih1FZtjaUIfa
vN/jBMU1z+TNPwZngC12UlaoTK7bLIt7NttKWDWj6V7ca1VIiE+lrXsK5Ln1DaPOLTnxWHND7oxk
EH27JuCfGsEmjRaJA5J8CnanG+fYG6KWAHbjS/MFH+ook1rmKRLrvjkCyphEBV0IHRUPBBP2bEZJ
iVxdLAKjC1dxUyQMVsWUaNXDy1MlSNJx/wPeO2aFHTEP6Ls8cPnA1Lw4obkvLWwPYGDX4WVKrA4a
gbYTdbUBwDYRHoLhzqdLFqBPr+QP7mVg0800nSkT90Ug2+2yVFnXPffuZHi4nhyNFj0AVaFXIfPk
bAiEhLXXumJr+cv3EXh+WOs68oUgopkhcoeVpTIboV5jSaoypW/Ufw/oNXEVpx5eyErQ3pI1ELCu
ofB5hlKcM/lEs6trbyELviFuU/nn9OdKY8BWkh1yemUa6nW0pb9Ie4i0/yX8+C82p1GX+137lPFR
CF3cdJbL7hwgPmVekQXFmz37uo5PyD5Ln0Lwga4MqXu2Cd6whJonUdfRHgF+EjdNEqnnIxWIVV7g
/Dku9NzJ4w47b5eqqsOAtfFJ+gS+LByQW1mq3D7axhmEtoZb52mI1eavtAOy4geuRJug/HzXnvqe
FdhxOLyHeAxcgYcwgtemk1Qrz/2OQ8hedOTNIh61n1IIw/8G2K7Jqaf4aI7jypeNKCRbtpTdvgq5
qK9ZqXoi+4G2NOMHvUcOEuixS3cuF1chTOQ/Bu8TahFUtqf64qxrz9T3E/fdsQw91qx1LQN/Xc2o
Ysw19jh5ZmNFhapP0tleqmUMLY/9/Y6Q6J2Tv4Hp928HVFST9MdgXPhuaese22I3xtLUzP50rgBO
XjLey4EJ/k+Qr3pcX8Cw7ObNU6vwVsSrfStDSy2KJg0cRxNIBSrQoqiFXS4UCGIg+9WhAXp0mk0w
4lkBwFiYLxk4MX79W/gUjIi91d/rYAV96OKqrFvRVs9ru6J2YQcDbddR99kCO8zmGuX2rxk1AzOa
4lQ9sENkXwhGzgsGTCLu0be5vzqt8WQ2rMfi/exahZtsXHYAozsBmjokROUOdFVuONx9LEhg3TtO
FKRb3dDhaKtYFZIefXnLYl8zKHJD/XlsjgT3wRzdEz7cnHKNWi5TRAFUpAeBwaI51UCS/AVBes2H
s0P2ABc5hjU0aCp0+RLmeAnT7nOyAgW0lVEJMCdNimBKSq2ghFd60NmST5J+wjdJ+JlzbMkWqn3V
nl8eOpdswZJe3g4tmXl4u9aKWAchW/F25wdCBCEmQ0aD9MFjW2zEdXgF2/uohMyXXUQG0AS462yA
hGnj0jLFpMKV0cOeplOUfHiZv4sO5d3tjo+U2dsSSri2DmmhfKgG3yAxjNuHpYjH4+5rxssiipO7
20578LRAIKuj7/MOMoVxbWkWG4fKvQjpKVCZKMnPJq2c0jSm1pRbxJUF/UmxR35mbG26is37zXFy
ZYA6TxQvtCJc45j9HQTiGehSO0DIft8HztIAQivXHMpWCJLrX7H6FPftFIMxzc2eoR/zMBp25eOx
euO2y/zf9r6CXdfs/mi0naPCHXsaY0nY3Yzrm0O1l/Q3cJyLKb3JXFU2ElGzELvr4iq0DS8pIlu8
q00zh7PYSWl943dZYfhTWuxVb2b734q/dnbns0bFxJM1hkqRvqA8TAD+VOQXwcL6xrIMnLrOZFfI
7ImHFujhpjoyarroHiaw2171Js3G1KKT/a31XbXqRKREBUwD95QKr9YGu+xSV9Gj113e5u1YGhg5
taVjqgdAIv5xtZipuMysh0Arjx1HB9nW886XJnK892NYzZ0xahoVa/oVJ5eEGfipoEOztG6240Mj
G3nzEu0y6XR17fLxuXSjXL5cZlNmuivShJ/go29fT40A3Ik/EwXQCyUPurYCmbZYRYPXVdfltqkI
YUpXCEmZvt3eFOawTYNmBm0cyf2Um7+xDpYJwbsaoWIjGVb2MfLWuNLDU+TT1ISVHxiOSqIRKofc
XcQqRnX2ETyJeTniHS7snevToGDJTrZcJTsOTdrPFPLYexU8NAVTF2m/22gDxNYdyKsBRxv7K1b4
6skpPFErY3WMHmOSthSLu5JhmvQW8Kmd/hhbaWVlSKHENeCjKKJzByYLivXjzGf7gK2Z6mr6e01o
BfPX3CLRh3IFoO4smQ6QSausXyCkvqmmN5M6cD7VoMWUgF07VxEgypXToA+U0NXNc1qykcOC0qoh
o+XbKfDOxWOUcKkEL7oJJlDRJKftgADEO+YuA1POnzXGjZS1bn1ibrq3I3zUsgxqAYJpX6dcftRG
DMLoANrBFyFfRE48BO+6OQRZSFzBkEE7/5RoorK59kfOLKfgfN9hMIJ3NIOa8BKWCS2t8Jw1ozKS
6zbx4zgb8dpK3y2wscNcVbRE9qO7JpLQ1iG0fKAfT30+WIGhlEESAbZAhY/ePU85bQfT186E+qmJ
b/0MFc79PAkhmUfH1Y6DfIT9E8kle7uVJzzQqH1ppVKYWfpeZpLau1GUns0zEHLMQ17CrGla1EWR
GB3r9h6zYWu0/pu7dJ3gLPYWHUYDZitOkbOrNP+ZgU4mGOQccmQXQ/q1jpGhIhDwtI5XdZ5PpU+V
XypDEYsgbAvQDS+3j5vCR99VagVUsS7SP8vXNkKrIVqmTXdMHdL2cFlyLOlYLDDu5I/UWa4ouGVT
NzbWg53lWaEgZ3X9x17FxupH8TDskR7jH1p7/4wpwDJGNaA2qa/i9C8soe3mSaWvGt05g6QdMD+H
EtHyBpHNUY5Fgj4Q0D/1ElB/tNzshuIrQH5W+XI7l63FoI6njxVqQzCn+84sOggAioJDR93q1Asv
0R/MqTWpKf2XBPiKNUoc5s/Ehpb72WZwu+8uRjDrjg1XBg/OmGUY8JUz315AM11ellMh7QiNg3on
xEhJyUITMiKqLLz4yYczT5w6U7LOrsykt3IR4GXd82E8q9xCW/YunUqCr6uS+7Q61mZxAQf0yMUo
eGvYHZaWxl+gChvBSDIkWioxH8nCael7YrYt7rfwK/+k5C9GTXpYulBL3768bFh3J9rYN5N2c0u/
dK4yvkcLGFXozoaD0GZArP+ZPO0gWvSbuLzTavBeG8FkiGpaJ64MQZTGvGZpR993g7rEXTVZwN+/
iL+Rw+rvCY/xHs20fEXCZWLvwhOfGTJhCZ8QuAcF7RqYdIFPscG+N4LAGtwfTuaU3jJSzhrB8Rvu
LE7ZBkMXt1cj/UoOzKBPQSzhUau3aPHswH27DK7pS8IELCRV6FjEBC2yL0J28YOBomhCWdgtpZNB
wZtALznvnn6Lo9cIBX1UBd2eZinMLAJhfpKjk16oJEuCsmPsU4aJObKiD32+vn0f47U8rnONgWJJ
gbVE2Uretqv9r1tEsNy1vAmdV1CScoZeaTN6FS/9bF6jGxMOCmED6OS8CGq72BRtUcWAjNZ+Qxiw
TTRZXw6giL2hjkECB/qR5ArPDQd5xS3jUMU8BeZdwJu9oELnhsekLR25wwc+xcKg0LmvmIr3xtih
GqxryibwojC7jxqeQUOLXFrte8CRXhyr+YRgjnyaoKh4mQtnslTS6cvFd0czQXKMDTjtqeWfDpSy
a1PPFZ0Iu3SVIYB8cAWQHb7QfCK8Qmkpd7xfQ2U6UloowQurLca/ji6Cr3VWY9xQdU7QZ7CqGlw7
VnHkaf0U6RwU1h7SwiSGuj102wRI54RJzUzyuXyRQ/7dB/uzm7mweDcL925a2feGNmOQnX1rRnBx
P3KTKRVNOy82mN82f6ZM4KKl3iNPtLwiC9FOTm+aVhzmkCDpBmP6fpBZWa0RV6M8X1kbMb56+5Hr
c0LN9mbSj6LSQQtaoSAdk944Tfs/RklBEWqcgXfZgAafu9Az0JtU1K8YIMB8DOoRsvo0VV8vzChs
7fiZodGSVY22ngLVACmsI6W+vA/szNRfGxwrJCq60eX8FNzZTagdx41GsSw71hcF8IfPfwvcmtju
TdICwceFltjKnTwtNafxyiinVNTNUwKxBd3MV6O76ydFD2ImfP7X9q1zM250wkymPMguGYDzyqSa
DsHCNv+ubCmAB12i2oVkJy86JRB4TOETf+VvBPyv2NBFhSH9WJqcpEgur9zmvfJiMja6xYIWsSIr
H9G9KnjyQRolJcIyu51Ya9TelZE8ynrK8GJlh0SKVgmykr4LH/FxX19XZNvTQ6rLffhO1hmPXaHt
ZYVzPYpsUj0y9k09upmTG4A1a7WjBPOWt0huvxMlxcMyTEuQolHI/P8pdddLPOSFXNYc7QkqYyd8
rslTV8KFVfy3gI2OllgfqRfNPriID6M4m7b22v5DW0SrK8vG41XkiyfkhFa/C7UWP6nzdl7qBy7g
As3Spgueq3igQtc8C54DcA7MgeZ5rtMv9BCcHBd3rU6vBJttljX88NjRKAVmIzMZ9cykCYXNFrtn
HJKCssn4bpA6hvutJqZ1f/vmLG3ll5y9UK6JXBq0TncAQlJno0dR66EeHX4NiTnVi25qYwFIFG7u
iUzX+MieGzGSz4n9bytNfiM+aKaqGOPYjVoLDB3ateS7IRQXNy6yDeP8QmY2exbCwmA1fPziUxiX
d4Mgcq13aiZhs8OMuH1HZ9iTLsFHm+ehX7qbDgmaBlaTGwsozFUuj3Bh4FW4QqEofpDyiu15lTqc
pqZtKDoMiqtU3rBHATvbbMZRUUBMFzKdyX9XdOtn9RuruAFr4ADuESSec3RsjopSF50D6k7JtRd3
b+dnK3uyAAbGvwH3ARnNLgW5BNmUa983452RMDX+qev29Npsk07FuQoPrlTH29pBqfYrL4YWZYjd
dmTql8y1xvj6lB9CKsG6MgyLKtjyQWW40hWG6gHymtgrTb5ikkVNyLQ5HBTKiEtXxWPFWuJEr86U
NC9kTWlHk4LDBO81OxBFUwfFjN3K68kwS/vDXbftuXfsT+2vJ6uV+rPUcwdOkZzKvk67zyqlmbkL
F58F5V42va5Du5DQKAnWyBCYzbJJAPGRN73jjjn6LeCBl3dlJsF6UIhCGodKbOhIH8clrKnolVUj
N+LN+TnYBnNjywyPgTpquGfaC8dXxSSJDzSltPHutQh3QlrQaLQMSDkk9q2kfE6Ntfq0Y6lnNgxy
vn0u9JFhYQhVnEUA39NFRhMsogpq5bnRqL4OR7TouLHRUDdoDbQKs6FS7vwEkYOXUAUw98Dp2moW
ICf29lkHT8OE1zg0V78wtH0dNwsNISMlz/XUexwbf2PUpuqgkM2LVidbJixi57Xto5tfuSl/iun/
OcdJbncP4FY5y9umY8+10KoBIir0sECnUu+CQCVSD9+FBk9mQml8Bnv6o3D9iv0LV3FFCoH7M4ZZ
eaCtKjoDW2+gqNKWmBBK8TKtDm8BwUmMXfmDG10X3ppSB/gOOgBtiiw/H3SsDbstqYQA0kMGN+y9
LF1oUDtzxT2q//J6VM2OKqS+3Hx63BqMDrcXji+nvWn+axQzxxM3Mj92ZY5YPvGgD8rMcSyy03GF
XlqfglfR2zIoktpan8jPjTAfd1QI77GuawMAXblD5zPiDUEKfemdy0dx53JoXjYll4PFVjPfRF6y
dhgi7j7Fv5zHwonyo9+6J0UjEcfXTl+ARIIAg8TaThuep2f3ZNDT7Te/LyrF2LqNmY/DAy30Lzs5
hQ1kD0FX0SHaFD4croxaqvIBtfuxdDgTlgQuXWVTxOG6dveAmBGixaom1/Nd9zuP4ALWJNW7GWaP
1bZHXC1MSU8KsL2Tf8kltgG2RimXZlgZsv97jXWXMNPaD/2hox6l3fA0psWOcPuWpkLm3qIiqc2J
uIZZPhVv48oOsvSqkMzFdWzA8A3niKgHCgDvgQTfnP9XPageAnWP7teSajkJq8ksIcL4d0o1/6Tv
Bp6WRNWJeCU3rMEN7uQ2K1zL1IbQ5g8is5Gkjh8d16SEiVNYfcv0o1aI003F3WxNm+EHR9tQfkaA
3JCpXtY2ZfcNz2tzr6OnchpO6gOsas+L3YqIBSXwugd/XHFWvjuwrJLiolRbPEi6F4adNSyM3TCZ
ufciUSoX2ih381+5U955J8Rtsscb08l/ZsTaqfK7xX+8/TrKpLyRxa8OuTWcCnpCL5p8VM4y3e8D
uF/AhrbBqutnvwBOvfZRz0aZvOYluR+mx3HQIfmR6M8Qcx3uIHGFWw5D9Zagf+Do5CTm+5PDXnRR
BQBbZJ2FgGsj3P2AHK5Lmvz3qlsfv6zkYqTJLu3YOue1lhXji0I95dQTRPRcbikl+HbuV+3LVQox
I6s8caJHb9sqTGjIxcVXMj5VilOfwxMbNoaQf5xJuRZV8QcntsB9HG1wxeWZTONRToIhIuT/jj4T
qaYOSiLOATSwtcxThrVj3G/TR86wg0ybPMR74WxyTtGbZ19/6leQx2XmAcupyXB8BAO1dyQvOKb+
4dFDpkVsPadzFvANKYFI1hS81jpBE4hRg0GMBVw0bbst0RUcXV6VWXPtjjy0oUxKLkQld2tLSJlj
VVqIl4S6vRWZwgNZjSCEtHzS0HKU7EazsUP7To221+zlmiOTphK8CLILFfAyLjsLH8kNfi1nXbIQ
TWitstUBB3n4hMp3gI/ZUhWIGOmFmKx/ry6nozHmq2T13EoKmG77OJnTQWJeONghO9r90gsbalyV
sic+vIgngvWFawv4fWE0hMsOg4lPtJHSbUlAeEwwATyPQrrzZKx0OSLmKzASuhtaeMJq9Sl0SWW1
i5PcWqbBHCfR5CF+fDvjnmQ9FOfjGQm5e8t7yGDnYO+tEZQi8GQ6LftxtzEgHwvUx8iO4Ufk5JbW
7xihF7WDaYmtmxnuI/2tVv5ZD9spevRXj5lzbNiSEW2AHu6zk+t1Y8qqvFhXClFEOeA0LR+u37/I
zrZr8+c+DilIcMDhB8KUcBa7RziKSqb4o+JLtqyHXkKBbHsex9G5Cn/DX78JdVX7cXwvEdlghJLf
PU2FT9t3QOWYUVGKY3hsxjrfaeXUzO5CrA7uU4QkDrVwy5oXe1WsH+66EOlycDB3a9PVXOsH1QIs
s3wRG+uBNIlTs+uZTfuyDPC/0kM+j4IoqLM90CqXghU2ijdBPCCUzffqI5dwBA0NTszdpHdTbSsz
dWOW7dDVLpBtzxhs6Hee6YpebAAmFEyfn5aLjZvOSpi7qLEFrrcAT5MiB7sQFUrAA2XR7pHwRqr3
6z6yxsajrH/u9BZ5vz6FfFA5+95IYZlTWv0czHEMTXnsewUpQ4b/S6M3QMjX5GZ8MHmOZJWx6OYQ
E7N4hqQvx5q929zkAiwafQjplojoZEi6+sZV5UjSAZVojkAbi9WMnQjzRLFAsDh5pi04jNcJ/EtF
wy5fmIFJ4M3DrIkKOl3I6NG3AfIgs8Ejwg0eFKyou5SfjD5IoftQKj+QljxuPgUYp8M8GA+6LaIm
p4s8VR9Sit62Sb9J3800KDWee9wNW+oycvq47+nGaYpP5V9nOP3CgOVq3EVYw2tUDVdleIwirv8T
PoTPuvr63W544VLRduivwLfQy2R6R7hFR2mswWn/3/Nu9tAW1+ks1L/2hE7VSK+VdQc6asXnUdJX
Zyz2/473WwGfxXh8BdRAeZdVV7ye9kErN7l6eZgnWXKb8KRW/SgilPMj0g13PmvVK3YSmF5xWnod
Nw6K4owm79f8mXrdL4xIInLKCXF1i/JCYbk+zfBlwQxp7VQ+wBmM0/R3iLmc5E2Ki15zsm7Wrm0h
YEyqFVa+RlWSkLHWtJOT1+ot9jccfSMrthpZ4ZkzwZyoM+4YNBwhOA6nFokTY+k1HAdQDTxT/iy3
tOiW93bLZkn5vMsD0B+q51hL5tWNZazmfS7NBNynhGb2jy2TsALxxkBpk+w8wIIvN5dioUAingVE
xVRNoLrXCZhrctkN2q8vsILiHQRC2s0qPMJSLw5PIBFcUJoDoBSY6tbtwbx9n5oQadfWviZDRMMI
EhYOGm4w046YtxVZWn8mKEG0pIES7FQ1nKyeR4NRHLMJK/2k9JN8vc3rYKp8ni4/8DPymOoGcyHR
sOfu4kY+y2jai936WF8EPPnEw4wRWQ/g8OYAI6EIKQVZsnnK93ltUPwHv2DqwPf7DTyslvfBFJwM
oiinNzPRZ/r20mXHyyzBJx+8QNN9rwvFeJipu3mMjTm0bTP8S30DTTByR1TCG3fnMeqYt+2Op+qP
W+fH2nFvMiNDMKpx3CnUJvrW/EF5721XF+LMOEp39ChWTeY/3KxAM0HQYVwge/0YQ3YDCDAZWOlW
ab+IxUAZPf+esGNeEv0ls8iqQrZdSWtO5xOedKTSkNIfZjhRgka4AmTqG7Z6NQ7+mXp+yWWG0Q+U
W1OfqfthU/bXUZD6OCD//CFnWGwUkZAUIDFLW5b8OlT68ekHSTkKcUDApQ/KHvep2arVwzMvbUTG
t+0c9tJ+xoS2+mqAMpoEf7ZVwMHAInqLHzVhmeo345sA/y53nF3VQtgFKI+0/7bVR9mmysQoJ3wh
OzeHyKLfRcZPVZE3C6MBeLt/FlcaXIn5bgpzLL2DS/fT8aww9H45LmWFHFgW4oAu6MEVjuV7O8CV
Tu5lCKBoyA/OSMIENQqNEx1JB9qRp0KvZTj1zLd159KvFqYLcugAzqakDE9whG5ahRLZv+n4NlE9
ywhqPm65y4Xu4oJPwoi0ZK8Ovjd9X97r9Prsbgt1kvlGyIR5L9rymfpqzYEM9pkJU227DijPZpnS
g0Tu50Nb8t/qWGXm0FD8xI3JJJcPdXL73mQ59Dpyi3OULKRnlimUpCE5NWi/wbNPTqRHUErUYpW+
RJ2T9JoWiek03tx0eBWRqnopkcbl3EV+JMCUopnDsq0fD1JTXh3iWv37kupDn6cDmMJqZUvjdGs7
L4sTScxRrXl/mTbxL31iyq05KYsX36qgbKP6w0Xx8OrweD52G4pfsluBbNr4Ko9lCt5Sr6PZ4t0t
E9uDfb9QlwAJ26rV3tlGhpQf2CuG6V1or4IFXCNM9f+IfrPc0XT2unCpEQQ2lrjJYEvudqHQ23Ru
ywoiRI4Ap1uKBqI0CicvLU3CM0pWTLRhtiFJ5zpbpL0MKzClKpLZQHfqZ5Gsw57NnWmGtLB8XORz
uEBGlkGG7cRA3pp0zykb6qwqI1OUhGjuP1YaDUQhnAcTRq8/o5osKLfWH4y3EMEXEdDjOMb5ckqh
NywOqN+L+3uKFh29FX7SJNbWiKhovKFxXslHTy4E8WoW57Vrut9JLpMcKN6R0xH6gaMxI8paZ2Q3
QZKqw5oa2Dkhow7kusBvhv0y8YXkohhcr+ryIlEkHOJnbplJzhtb4zaY8rYbtcX480A+MoIfsCo2
sLeVbQX8ob1MRsGWVihKZjIWR8L+9H3LUdLMq2dEDIeJN+kU/Ff8AW5S88ZpXE7XdyeAL/d8lccY
YSixtk1HV4p0mmAeZqBpQWPvIgXGJquDXhb46iqXaRKmtgyiu8qdiOzBISm7xa40TJ/43KlWEpCz
hWBvrcB5W3eG4zOhWucAFIkE+tT8FhuzEOXMWCnmMNcpEhQxgOPCTJfzlOgfulRfk3FPRfEGhoR/
EkhTyOQdtwYrlNhs269veaVzEf/sNYLtr885TqGMzxyO6GcjqNSjsVMDDLPEH3XNhewY/gdezGmq
n2HLT8qFXC34uM3webyKKfEfqVuc54GyaAr6c1gNEHbKCpb+U04D3jFamY6Xu4Dk2qiQR7k9KjL8
LH9OhKQWSfoeOF56jyDzmeRTHbGRdwkm9V3AdhX4IcaBTWoMCe8A4SSVVHFN9rejyfBfc/HD8fHW
NJzGUbduPEdQd7mA2pSE1q07Csnjo11XLLxVlFGA3O8+/UrCbAiOAdmI45BjhuL1Anfb2wNPz2JR
milZ/QATVnh7bNELqDtE7NIZ2I27g7J3B9cYB+D4daSe5g4693eRtYG2zac79G++XDpJN/jE4MuK
DxBD73ZTdpfSdI3qEoF9fq7B//L7kknClxsex6iRe2Ef7B9pRnWKz5dXPF0Vm8LLhC9c+WVgkE/3
E1Guku4tv22H8TUDu+QajFQyrljdnV8JFTNGDP+FMTiHCDClEXN9WhRXtg/7xDy6VBjXQ4tBJpjU
bXHRVF4YWZbRj9OHKhO0Lvw5+czLfRm2tcC9sIdkta9GJqKDB3cIKbGFX4hYhGGpH9WPZz8hnN2H
6G89AlRGnxr0owO6oq1apXGbWfmOCaWpZF4/2yAaHtTnNfIvoVS/WjuASacwl7IswRCnnatVWEMd
KpsO7qTEHWQOzgdLyKNZGFRB5CoU2FBV5AlL4PJr8fsn6GUZQuqwqXKFIlrTEUW0uPV2YL+zD72x
DSv+si5dYFF6B/sy5bSltxluphN4CBF58Qo2pITUDAIIJnGwoOsSWrBFLYk1GFekEj2Vs56mw2qx
J29F/S5JXUvGdlJb/60RTd/DKtAhej7Sg7GZJRFiNZRj2JzJClp9y1qD0Dhpb+TxcqKH5aP8UAaY
fx7DX5iKCvt95t9U+PEK7ND9K8N0L2d8o5+s4qdJiRfM7/aOFhQH6pjM/cRb+jKXUkhc++F3vHeN
yFRnOTyD0Et6zSoNMAzu5m9i6mtos3HhRWFzSKkt/06GvDJkTQ/cOMyuIxTDOq/VO0Uzc+I96uAm
FAwH9r4SrYqliJ6yOgfzgjx8hjuB50pdw0Tdig6XQyMBGJzwFiKemtdelQrAdrrPggRgskjV1+kq
A1Z2/0/uYPfmdyuErvAPP/9GT4OqCt1RHkiD01YTApUjub9fFvxWFDN+77VtgTQ7t3iVNSqDueJ+
9azhrsfAg5QhZabXAi84wEu+hE6zvZTV1I1bWIrTb/h/mQJAE4aWJ59zj9Ds/7xN3/mqPiQ8xMTq
FO+5sOnEfTuzQuTRJuFzH1TkpQ7jydW/L6oYdYfrs7xdwxNdYvALw8NeiZgJGJ6s9zz3Rc0qr17a
Iu02m+OeQOmiGF6svXAwFPgAgvts7UPGmq1HdIk3Hi2Z9RoISs7CpgwiZKG8XgQekv77rHk5LNLz
WVqws8qPM18dw0QHq2KTJlK/RB5qJOxjumcbpgbmj+K6m+1cXu8MJP7XXrbCFWkLDP3/dQjqT9al
0fZNr9A4XdBQmQDJ+BUOAZWnuuwg+RmFEBrWFpXNx1Kp6qF6jhTXq0aj8m3O2H6If9azOW5XqSaH
rcs9YS21/gKlJxk2ZXuMf8kNEf1Nmv/5dEOH7aka66k++r4iCnC1OqCkcKlr+RaQuYZQ0ceYTJA0
PsMK6z/zGN1KfvHSEKmK/uEzatrLhI6qpvNa1ZJ3uR9GZWGURii+m1klUlt80oKiPSHOYyCj8ZmI
s3rA4b2OaIoAnSsFAdSlS5VDqnEttLwuZq8mohIIm6FWQBkcW2H6ZyX0QLS3H6CoC0zORdYwHiCk
wTIhSpAy06ReVIN7+BlTwb1LC5EhYLy2IF0+hCvwcCnXr7zshE267p7Cnjt0aZCKzzWW3oGYNaEl
x9U84OLCQYB1AghGr9BtZSWHdSOQdn3G8MvfrBxnOHayR3uS1cE1vGn3boF7UcXktrkadpqODmOG
u/H+Kq7Yxpr4yvxSdpFCuYClaarg8bZi5k67EGSnTl0rVGPlfgcJNycqE5qVgB6fhAZADTlaqGkU
0JyzwXcB38vlDXXIkPqWe75WrVxS6D92jpwVCDyzWpLGWkCVltJ7Sqhpih0/E/aeRgAZvGn+0Nle
/5RbE2BgAYu7v3NPkpe2W777SCW8whjhkOr+c95lddrHkNV3qcawO1dCk4BqTwgcoO6BsUj7er6I
Nw3E/uKeWDtot7fDksseO1P0vxw+CV+u9qa14k66HSPBj2JzwR6vZQCcszGvZp3wCvmSblhqMZYP
klxY0za4O+ESMcte6wY8M+YRdKZUjKjTT+wWEqhR7dN8CnJh52XP5N2/vqrYD8+Fz16orhUNIyN5
ZWUrCZWeG+UE/PKMnteABqk/Jr8PTZiFUhuOnGqPZHqG/d541xxUGp44Q8R6vZJVZPLIbUNptmMA
mbaOxgozUvXnYN8HUarH4bjQhqLbYEm4BieE5m2cSok10/gCD/EooKroaQCjS+zNW1Qeo8hy4F4r
RxzAH+PI8lLw34Po3YtkN34bHeNfp59J+tXm/Akqudn++wFWZKFHH96Z19tLTbeppAzCUankBLgV
T6HXN2Fhuq8WPOD4cTDlgXJvc6Rmp9SvdMxhm+vGVudx1oN9I47pJK/1BuCQGxG7hhuf4RoQ+m33
0nLDkW1e5hQs+6ED6vLAOnn34cM9FMCneQZ6m0IL7p2nd9uWv+omlU9vYlo3hFfWL7NmikLjNoYK
7BjHnZteIveD/plTdcKQo/8g9o2XcPxZxWq2sQ7MTD7Km1Tafop8AQd9jzXMPeyQ6y9btGIP2Gun
5WThjxPJvwLFsU35A/+v02DPnL2Q+xbAMLCHlHaC7ZO3Bbd+Bdia6Rdz8vY0nPuafwYBIuNnJYTR
sYuu2/mA9XofVXvLcGM5IpxmAx++4IREqsSnNpRJqZ2XFvJ8rAfHs50D6IW6Zz0H+3RPRGniZqnV
NM1CyZqHJwv2Sd/456ANMsk6QZFpG7c2cofDH3+3USUlCIbIHJIuzUR1n4xeHbn417ZfBr82r5kH
RtlCCLViGIqqFOKfGKZLec2hCwEwQM0Ojb4i0T8v9SrumroSQUeMs0Qafw85PwWewVpbErWSiP9k
XuMnJSRSXW1fg7rx39VMEWKvB849lbtCHyuirhccUP65xK1VwMdeW70eF0JqBIaa+A7rCArAPq+Q
zes8NLsZABhqIqBZyj0BY4VY/XqiVTBRc8HJUsaZOllsavRGB0i8ow42beh+gXQCUmJWyD5el4Sz
537+twg22fiAukTtZ1vrq6NnGF2P9VS1FIvtFHRi8BGa8zzVL1NeL9g+PCpMHuSGioebrtXyh+jS
Ngtb+ozKHkESJOJ/JDCbQsx4A/e9oftfJnKcRAhSgI7X9FxaA4/0KB4tlPZ0rpWY2OeAoICVWB0G
lN4N0lLWjJ6wTnoZujjTiuoGLpBWrExp7mhXnopy4byF43XKXOhErqIrQjWSpZpjatzuELZBbDdn
rpoYFTzabUBCAN9yC6yX+K1DSTzFYMX0F54mNZwHiPbwfYrqpSjSBV8djhTBBWVVW1AFo3FMxnwn
3oBU8MItsoEyYizSOIWM5TA65bpOrafvSjd0HZDIYX+CyyjJ2JCCwN/g0bpsa/g3uOoxoaNTCmTT
skBDT/eOXvLQnlkZSnCN+jlk+XQmmOWdRXj8aSgYU3KPdl+Y712dbWcq2V85i2x5lV9E0G5HlQa4
1NHPQm4mJItoo0PnEFT0n/V/DWzqnLhcId/f0cmLUfhD4fqMFBN7ahw2C6dvcR2iQrkhiY8a/YOA
e7fQ8Ls8XIaAJxze45t0tN7ffBIddBqWkbm+9MQSimjBAO1tU4KSZJ7KwnCXDungeEMGP8aacUhK
Fj5GRaN7YSLxANnqmdzQiW8MGlZbxW+8RPb20+OCqbAb6LEwW85ZZ+oN+OW5wxUsj35y5sBkv22f
hS+hgUL+O4mlISGOztBoWst4GUMIi6Kq/04CSFFmuMSVJeqLEYk5BMwiARj2SQUBoie0FKgWu4sv
olVvfgFChjSOnzBIIv84/SWBfk0dfGVf176TWnqQzjSQ995+M7eb376uPGQNzXfUsB4LyjCvhnwv
ngRuHPz1VS1MlxAhhjs9Yo8DrnNwYc1SuBv4A+1fYof6Vc5spSqqSI2Gu5SdUPWbogJ/g2jjbOzd
8n7sHsVjInwwM62jICyfASWbvWMSbCRoWW34U/c/ep2MmDf44DeiBGkuzuHb/sY88JuN8BxCxzNf
7QnGLiShEglvtXdUFuVGeT6qPy3nmMmAsAgDhwwGz2uIhYcJVccYhfe4ZYL0+QRB9R2mG1Val5v6
w9rfULggRwtTNhMMECUwa6RrZRbY6F15ediocoS/Fs9q9xB+71YRK13uBpoqXggH1xnWbx1Hr+Ym
Jq6oZ3kC0K3kqAFQJLSeTxcxHS4AziNtg4NwK/tEq/jnestkZOqFZ6c6FO27SFTm8AGMefJQMJfO
p1AcK49VBEG1TkUCn1y1IsFGZyIm+qjuOITUnTMHG6n+nDa1rNwu9bHwRQsXsY5b5yQkotQuDF4R
p5wDPbiwuci5/Xh0T2Jc1yA/S9R2Jwvocu27xCvbl6HRDssGjyIsLjqeSThUEYq1zvZMzjBGTknh
E+wsDb5xYA0USwF4xbFTm8rYwXqLTxW3UipNw/itCBNCunhoEBNMwqv5IwgC4ol5C5M2M9pym++s
h+euKPquSASoL2kl5r8pZcogVtNPR/fPa3a8ph3mmQ97zQpW23u6vGzGNkP+rOoTPBUXwCtkwMUp
8Nuj4++SBKgKavWvvdgtE0VcU0y/4inCKxvYmiv4FWsoUqmvwvZmat3d9gSV9i6RwhOpmbu7lQWd
/Cq2ADf3HdFLcInHTlwD3IRMKM/UlIuN17N1KoyDMDVY/3FLY1UlQmmLuoGU9x40prdp+PIzAoDR
ObHviiqBb/bxxR4nUMc7jQsgRrjSWuwhVjU7HlbIKWFAh6IrC3hDVlI8q4V89XAhczb7ao2izV5u
/uXXT6ZbcNH5K8IjAfqFwikkQRY+Z6s0FhQL4oF154cxHxaQOorgkT7hE3mraUSAqpG5gPFflOmn
eptP4fa7pWdr9v8IB38pJXyY1orQsTReQeqf0yEhsnn0Pah1mWyF/KQmyiRunQ+ercYfRjmsccyy
grVM+F0ANoOXNvI6s1cEoLp4ceobMOd9wyK4w5Eq4LatCJEssOTwSuv55qFIY2UOuSNm8q5+4Jc9
4I21Nac3Z6/oQal7clM66vdQfKyZoyLccMg1Hc3kdN6SxnYTxWAgqUFleC8g6PgVZoBB03ub/JcR
U6dWfaJg9uQf3PkQJk5mqLp8P4/IM1ImVIcCPnRlg+nmnkFlja4JGmzFEfAFaC4FEHEtty9ZQoSj
4cLLYYW/6Im2/es39aLKbmL9MnDfYZEDqkS8c1uBwLiLmMbj6lyWjhj530eNn1cIi7aSJfmsd6L+
xzEIzMGr/DaCNMA/UgnLMeHdN2EcrFyPkH+0CiDKqbwAehgWaJGAHITkzAb2yqPsRrrd37Ie0MSf
3kZzYyyMzg+u0m6qycGRzchFn2ryIuKTAssPPkNIABRIAiwdfY2UcV0UAV3Cs87bJKlpEgj0S+Mm
1XKEsxOO6rE5ZOGRWKtSvwhHqLuJtPvb7uUmEKN9vo+PdPxJKCvGpC7eRz95whXb+TQfYd/RKDvc
QEKdOvS+ZOwyCwmZA2uoq3KcWmwnY2jU1U/MbSb/QVjMSW5ap5TfYDobWoL2QVStYSfuimvlQZQP
BtlLBeDxTeTF1HBO2/VD7GiPnca64nzJgTAp3VogXKVSe++IoXVfeTcJxJ/FT5NWMbEfZVdy0dvd
hfiJ3y38p283AlzWXIU9pJUca6jyA0DFhYqrq8N22AfPgvdVjegClvFG4nVrv/ws3cMhcKP1yt5Y
35tFBqAqGPRSqE+W9ArV0ID9sVLtvrXDyW+whQgYWU8vAUtf8OhMvrWKr78xgsuunyrdOgyDOxNL
S04AByNT43UWEvMWLcaqz7nkynA/UBQa+fLgD3xWtrXZW9Xcd7XjeMMWoSrRYnmCkqdl5LnNxwFf
z5FGyyx+BwpKpZ+Qs4cmVOGhfHnfvgx4VV/xYJM87XhrdZHGiP0i+9fAMWlEXNZH6wR/jTb2f+l2
heazwZhZ4FG+r8Nq/bhJPjjSttZYpKgZXDU6gMGvVTOtaak2nPrrbnyBLKygVMeLtKjh4FTAA5BH
DG0JoKS27+JoisVlCZhPsZ0I9qiLEAxgBa8e+saRIbaEnH1ZpDs5HvS09dfR9eP8NorOendfXTcE
LDEUggKDJCxKJtqLf542RYA/fAx3J8LytHS0h/6AFRXlomD7AnRbEBgTdJzJ9gz/OOWKF84TBwY8
vLWCh51feyyCrzZXn/ASETtypwhvoytbzUOPRChYTe5gIogGdcuuLvKdeB3cqqyr4IyKjnoEgr99
9pYUxjhyDVT0ncrHY7pqCWzHoCSCjkQhGvke9raUA8n0gzUUFPVHsryaXHOgIRe6W5V5LYShkmaM
cObdF20kyyF7D+LFco76gsD4SxwhbRhhGE/Kad33Dsxb0TXuuEgRPHMTLu4R3+BtljLqolmnbjIe
t7EIIFoxIDPkb4L6o2AzCEAQHl126gB7oY+PRrErmCnoqHgmMud8aabmS78a2fDhD4Hq0xUYIQYJ
DPmdLyqZ6rgWlmoBiQrps9y8OUkaMn1j/epEUstjJ49hdB9onpfgzlRWgvITJXTj7dwjsLwBTTS6
yNXHEgaGTVogBYeSkNLRPTAkCAXp9vjuwbqT16RtBO8BcgEcJSS6sTt25Oe6jR90dgY/Z+Pj9gcV
sVPqVRv3wmZkCa45te18t5BwnMA1EcHW6Q4mzManqnUcxNYvWBLHx3+kYvg47DoWdbehrQwu7sbN
H0aDG8dhPXxwJEldPQ/lXlGWk31Hr5ku2E28UKdugxI0qyXIdh3hnNJ++psIx5V91bqUtBa4rmIn
Cq5VVpC4tdYO0P9GwO3EmUK6zpSjEyo1d7Sj0pkvPg1xFcSP0kxtwRQE73YPbOXWQMPZvcrOkE90
+b27f52E7t3yGzznEteoqpkHp5ufNQKWePpL/rjcpR0DSJgoROUcd0huiydqtH05vKvY+UYZvivd
HAOdfT8LbJ5lqptJjBCYzCtXstlkYtB78bVgE++JSnPoqbSlJmjsN7wopNCabBwvo8GH5Uo5Dkfz
1icQrX2YZH33gyoGPRx8ZE3c4rXS6M3jfG0XdHsXTOl443pPw3gGRo93NIvpdGOlOLf0w3x3K71r
4m/t6J8VHUbuAi6I5PTXwh3D1V6fjnpAzVwMM3S36TGUMBYZAaDt8auMfAzMkL1C+PFny204b5zt
5e6D5yHP/eUTEXGO1MxnYXr7jBT6KJfQJpbWBjY/fsNYNHRDQ8PzbSWXqbIlp1V0bG6SKKA9caLD
OWawMd9b9i4S7docSkuTgBStQPvUlnv9imKmSJJgcJ0/BwrPRjC/pPD4jtuOf8z/oIJS+eGNy+4p
si1hdZjKIGNzQeHNmu9TxCq+KkhUFqbAlk6Quysg8HCQCs0YQYk8FWKU1pVF+wCxByeU1GlQzIWt
2VDmVwXQ2e9DoxNp+LR1jo1io+MHY24roSChE9thDGb47NlnRenWaJXlbsuec4AeBIdyxQWVDHYT
LAPyiFsXXOSUCs8CmfMOjrpA2fffjLLPH0elXQwrQN5GS5sCeXHuyZxR5gEbhHTqrUGkBFMG1oAJ
dWBjgaQHvpD0VWS3L7N5UAkMR128XsQ1K3Ai2dyovnHesF5zyA+tUum50ir4zausCBC5nga9tpU7
lDV6tEAKWlDa100TQWaC8JVBl+z6Hj/KMl/I+t43gGflFenWtKZVeZmww/dwhNPHdjqXeS8UV4wV
R8zebMh+oGKUlydFX8THnqZ11ykxTJn6zNmKOIj6wi5QgFw3314lQ4JvKlaYNb/Xy7hWKCTBCYJC
OZ8qPCR03x+Uz7GZzI6btMN4Bda+e0QKlM77MNAB3+iSDcLn9EYHbkm2g1s0ilNT01wn9U+24diw
4wTEsY3OaPqB+iYSl1sguenkBwR6lonJH+BSITB11uEZL8t1kd9p3Y6r5r6UQ/nDfr1P/1pLq1Ug
0hWQL09Xjl31w3FcAvIeGSO1nA0nGhSPHfOqw6lLmK7RuhfcHiutGlekL1/oefVIrrtRdQHpiyad
kJioqlfKOXkftdxuuKoG0HXvdEL+dZ76MO8Q7DzXL2OJ8Sj8TE2ipZQAd9HSJyuwgRN3O5RfJ/gf
K39jBKntIa/nORs6Y02YOF538OGPo/6/a2M85Rhm2mh/b0v9MRi/1Ty+/BP/ap5N5tWhEkgXmg9F
aT+zhTFz7JXd5H6Ki+v0kPOLaMPH0n2HsiiqCU0A2mgjl+7IxKhPBFr21yskLfPxElOl198dvc8Y
PEab1htlbFeEM4M8PqTR9w0HlS9AmHbm+DkuMShqiiqSqXqEbdKflPEn3tL7iSPemLgnSl+RWOO9
+PcanlTx/tUY5/Cd0yFdu7F/P2bTXLAQuh49DtVAVdQkKWhZRqHqC7FPo6f4yEXV8deXs2gggMxA
4kBCv9e4f3qcleIYGBe7aIO3/WwvGCFWDE+K6nliJOGKtINoKocMlE8Q9dsmscLCraRHs+eou4K8
cqavXdvwy2YQ/1E0rf/Mxl9qE3WFVBDuIzUN7qbTZWwMCpxfy/gg3l8ZFhkZnnSuelDyBV4wj9nO
9S8nByeCrPaz6URsfiALK65MKg+ChTFN/nAt8jqpd2LKKuMzCqNPOtLOA4cTbPKc0p00+mkJh9cH
3h0XAhXMNW9AhsttVjhuCgASNhL88+Yrzb0k9pl+vuO7oyNr8xf4I44MFCyYlNuxBypYZAiCtAyz
YKtwySkiE2rKwWA0CL0R+smFZT8ViBPjyPEO7b3yVCy9AixJ8ogZ7lQySeq7vBeFqbeycbw9modT
EbCDOZka1PYcjotJbFSQrbPq3h8wYdOmB5Bu5b2v5ohy3GsCCRxRkcFf83Zanri8WChL7QlMpbqx
NwFyu2wGWpqbwkchp2oEiY2POVPWuirDCoOcvQ1rhTFbjBJgSGp4yqhz4hU0hox+tdRkip/wXI2X
XsFZQuuXyUVtnBVwSrqX36boMv5QXl9HEJi/lk4Pum+mGM1DgqCA97yox928qcaeTaLOinQJx8x6
rk+u4fB+saJEsK+OvBKW2Cimn3jozLZtMWcfJDzVsGqsrI/7cUOUq6jIjZSe2NI78gP/i6zPMToV
ZBR2ASM/shp0Mp+fUpEl91mCsZ3kGuej+TRluvXKf7Z4whl4kvfIhWyXxPxb+kD1i2twtts01KLP
PnqdVFL6wS3KM2ZQVDFVN8P/xJXdFlARWya3IH9+h/9RjS+h4w7XGW4eTSXEW0a7tyQ7oyruFLtk
nbO/tMFcGnYVu0K+QzhDpLacUarVHAtWmjVR9aRt1IymEGAaw9mi/F1ZJmz2CgBFvBI0JfzaglD9
LHZBhQT+SkO4rDh3IOnqzLBPtMw9jDNpCJZQdYq3IDMUd6Jx1jvbimNWOQodA1T8Pw/OipOE7dX4
j/5Q7Cugjf9usVnKGBhQfX1z/UqkOdlb/dNNEs8bBuTt6JRE+IHsob9YkK+BcAfjVAGZDcZOUOmF
vEvJv3RREpyTTgwFGPgWagOTGSplp/nCyZYQWIvjGR5KuOHoi1OxT58NhuJJjpnbohae4Fo/m3IP
vbOi1OHFpOGUAPTtbDiApWnp2VyY64lnFc/gp/QUKyraebmmZ+Xzr0xF1KHQoyAcQps59ewU4ZU0
T3ZpekBveMJmH0cyY9cv9TCOIZOFZKgupGs7VMFQtRmT4G2DHxRmVlxqBX9h5Fl5nP66b4mEiEyX
zYA6UbS0mi1IwHo1k+UKhYuo+JCSN2D8ospwN2wW+7NxPKF4Org/wayjVONhYETmMtnAv0lvJEBT
sv8tF2ucXvVY2M+uZPLgEK4D/ZLS3hahnQ1DIvX1s3LeshFSE18AO7CoXNtML5EbPUljSNPVWTXe
wG/hjCOo7IFs27fhZWPZ7FT9Tbisf9KwH0HyZWRugoDG2voHP7F2NkXAVMni7CCTetaRwbW4om0/
Qr/NMXI8Fwjrhk0Elr4sht06miyiMfRdj6XBellBLhjQ3ErjxopQ+PD7/yXSDiDkqAb6eRetfHYX
2lRid8FH6DHtqpXnyIGwNJgUGR1gp4d/46QPLL6TUiOL4aUheg8qSlXHDIts96Y6JkEUaZXHF7nD
JRIKE8wyRfDDR9S+gPnsWQvUpcSafYpC5py4e2nCpyyQ7oDUhFqmwSD0vqIpZR0Wv8qoHSwsq85t
o/3E63cwLXegYAu3hHS4MGeyRdXpNiWhn5akAXkG0gkKAZ/VW/cH4+hgEHJS+EL0R0L8AXPgCzuh
xB4pBRWfiY3tMCcnA8DSzV2+qaUQg9CCbVIO7+H3mtYt/iaKEz6MPEiQkyMl9dZLOu2cOiStDAlA
+FS9ZXbTBINdiufLDFVGBtMJxtR35kier/HXqybE2a/ZG+bmPvaHYgvXVX7MGB2iXKtaSr6LF4H1
K0tkHgpcCPdBegvVcnYfbuj2YPSt+J3BSveqgUGFOHJEL0JfHgcSwLKGQoNJBaEOlioDv9XtvyCf
uhhWRmnh9byKei9PNtzKZDB2ra7HsFXPsme1uTaZhOD/JxafL1PeZedGxrsk5dsJVHHfQJ53Pa5N
kTADYCha51iJRbCQy949mssga6BY1j9IZ8TUwsyvKHxXSWT7hhIZMf1PaL0wf8DhK0qk3qjbhiVz
NDNUqu9ZdCAuQFTZWpMt9WnIXw6BzATin2StUugNdGW1zHHlH8bTePEiwQfL9/h56HASuJ5fyzZb
9dbDupfUQ/bnZieK+CTvKpNAet//WVVKC4Q3jXH53X3QpZk8i98ydoNFHrHknmEieGg8fLuGcjVs
ZY8YSJemzQaxKsFr+/qB+hZrhC1i65q3z7f/4CZqwO3FRLcdVLAYnwDZ4Qei/FCNZsn9Ca18T0ha
RdSYJF634dXWgJmmhB2iXe0oHPa8DDyA9xA6CYy7FRQFf/seoJx7EIa8VTFKnAtx1vswOHgVMpR5
az21kLqw44tt2PrOirWxWTvkmyhgm0L15NVnBof5SDO4VaBfpi3m/EtYfIB/M7tm6lT0DSSRFr0H
Z41/pmhCY8jkNJ7kM6wt4l2CDHZ9buitAZfHuzAFSjuzi1YbquhcNiUIyCsUU9oj49ISvPBvUupH
YEqjEHxj7a7TxL0hMznsZOC8iM9lhsheD7GJHwqvyv3v2f3qfO220/ss73NvBis3EbcGMZbmNoTQ
9D5nYlHw2FrEYVsVP2b/P7fVNq+Em1c6xcb7KMfYTTrATNteIq1B/vMewJk73v6FG5rS+d3Z6g9x
R9nop33tsit0Kef+rqvh5yPJ8bKu2Io421S3MJomLledntcatZrR5ku2AnFHgyN+cf26d/3nH4+/
T3Sa8jrXbE/SBieu7MOQ7dFTlU+f7vt1gA7XojtoSx/UZa7IGSRfk3PSbmwPD5aMkDhf2wtnlx+Q
JmGBvMZdS99f/WvOjM2W7lQoe6iEcgf+6QR2F2xBwuQ+9y4/7t22g3EjiWuWVchpizjlsfPEuIf6
Ys3nkeAwWdY5kEe02KTYCXV83MdZA47LQfXQ+iRA+DwyDC1wOlpGX6sHr8lLEwR3M5DRCJ0zEIsC
ERA0G7eT899hTbfb/6lEHmpMLX6xqSJEEsOg6jo8VJbHWYa18Kzm6i1Uu3JPgdVbw+j6NmJkIoGA
OQkOGi2S3XO7Hmbpiw3aezM8FxeWW+sXegBggy81LryBwZ1e3LGEEXvuI9fGgIK8PMNf6vBgd/2M
UDhT/ooU5qdsO+Cu3z0U4vGG/DZVhDfhjQ9Pyn9UqkSUOTXF/LnIMZ/qxecR+B+bDc4EoBfYnSFh
HhyFaqEbNWMOgBLqUqGdkbJVpDtzsaTkWtFD8XbuTpoLgsP6A1qHF4yJzkPh0KY1j4DR90VXkWx6
yypHznBpIj+3tfuT87CibxBYmcdHnfcBNrdlkCY86gWs9RY3rSccMOcE8DP3p+27O+TPueP4XkYr
1pKnMEUQAXQDhehiFJQsoiLCxUuJ5/KqAOm9HBXaYWlPnMfUSAX8PvSphHh6D1QENGFKSPWjaiuv
iJjHSFJjhV2s1rdEfLwaJT4Xwh1UoZR8ICxUCQ131aQV7UKbapbkYiWuGmtCWYOIPbENqSYV/IWz
8hCy/UF1qnycvmD/2OJ33W8YlUBBMs5cVd6rsAa9U/RCrpCpUr2CMfCR5dWEZ+BhK3rHslgdHh+n
2+t5uYw1ARP1IioA7umcF6UaVv3ofDo7vtvlJ2iAYTIgy/ggDJsmzMRQ+KkK+LXoSnr/UdB8nqix
eA+jLITD3mcPrtL1S0/A2E9ttdcXzWHB+U40as9tBG1WfSQlRn6CDCZ+xLDsNZWAmbGo8q0NKcJW
Ap2ISc7aZsEd1YAtc4TBF+xr+NpUIa/KFw+qydHtTk8OiHpabg74+eEg9U4H+CqI9SfvC6x7eGdZ
bSD9ElM5QVZikrDxgcCg2OrI8iIOPgBWD2jRWd4r4lPDghTYNry9HUl9wBw+3PlXEMdFPsgPIzet
+2o9vwfF3UmMXggsUR3LrkFKctJwtVYRmDDTBMRvWd7/k6di8ZI5X9JBJmfbyolLflfK0k+Ea+EV
VDE4OyIGRTPCI/lhLntueSc+Vs9Js3xTRdM6LePkBjMjbb0g4sehlKD3IuZQKBJ6+vFzWnYlLzXX
pIK+3LVVqtfTwSIYT9krfiudQteJ3YHIS5Cl1MyuGaOoGHRNQydYGIsbjas5ArIA2br5R+XDjpS1
7QHApQFoev1UH/PQx1CCcju0XspSoIk57X8VzsbA8I2/jnLA3Qm4NVRJrhb6KkSnOxqqHe9hYqKj
/Fj5d3LVgwTakcQ7TV39uj19eJQF0LcvvNoWZklOQ2jx0T3DqBt1NsdMsiIJgIz1PYiPyKcHHbL/
TYUhfGuraCvuUlZsSkyaqhkVDY4V6rfZYnZPI8nFpDZfYl0L01qMRShxjQ55gdu5okBt47WIIFsC
UOTMOetvlo5JxUZP7W6pJRCymeedN1sSmQiFAFc4jaurPem5wVUCNPEvwrLXYVQ7t3oUKZODZgfe
DoS3WRocB6+VVlUZ6+07y67bzqpU/86siW7iV7SYdU8BZFluVkBaPenuAGDW7iLP5UjjrW9/N/aU
CbOjxv/J75eqr+8REDJmKF0ZTXF5SqAdvISvhgbG4zSiYjuwdcd4dQD+gRO2cea2ETLawQ8QTNS3
B83eMbOEqmVrkheeJDjjL6ixctm6ZaDNyrV+WGKAcLSCbOZGjbTT2iwTSX21aW6EiNg/AUI9XANn
+dxR7HTOIL1nhGT4Me+gIrtBX/PGXOOQAMsOnN2bc+uGl3PIOjkD70ZvKj62YXOnuldbHUr+SuZ4
NOPs60Z8WS3IL5NaAtm8BaPwskMCwqUXRxhKgW2fFR0wrv3LjDZSN0ZvGeZIzWnoAKkQdkB8oAdH
BmMKkqdtrnOwS/Wzkd/vWvBRU2Kjti4sW3FmkLPSEsu80MkpzQLSkvMCG41XuHuIFGstpJ58Uzk5
rvkIjDXMnd8wuOgFtpbdphP+Wirou7++m158dnxfrnMihVlGmCaXzv8J0h1jCw6HbY83tQeGs7H9
3RRn4+Jfld6R7lrDLzXl4KtjHz6w15tb0jpTKZaipIG0ixiELi+W4pwBWzIXTJfBJ7abLyey7Tw3
TwXBsOVJEM2+wkX8io04zOvFtuvlONAfoeXrMkx1OlsLhobegZyXOkGLEifIan5h8IuQuv8umaIV
0jNc3LkBVeSWu19vC3E3F3C9LRg+iXrmTuIE/auUStoXKZyHOepypEPt2LCyqYJzSQwk6agF7OHJ
8CfKU56lI339O33gQdbcG4L8SEBbWBRqa1rSaFRzw9zgPHXA05dpY/BRDD+qg8DfoBaEWLqCHXy2
zdMOeVI9Z7wYH1/agCvIZZiMsn8gvgVmZVg9Wm+gMSX+4nKqTNahMSocf8CPYR/GV1CHfhj4zKcs
RLsMyv4UXRYGImwYkYqD4GHG2Cvb747sJAPvmmr+0tjS0ap73TTbkYQHnH9OtIQc3zhh2ixhWGGz
8p6GgD6tEHrk6nAJysItHStgsI96WotXdr0i72RI79oHqtRdUSpFOyCfaeQeZRRIckvMPxbgPpx7
05WkoNX332ChHMwwV3gQ8u5qSGZwa173BXvkjxwcy/uy8wAo0NUnsr72FBvOtjEVkx84e/IqtLT8
C7/gSC/fnKSW+rHSU8NbRIIswrqgAjXWib9GfAwlnygIT2ZndCJ2saLn9nmnqRS407lgy4YPhO1/
P3MsAV+rufkHRDfPTe+dc3B3llSRap+dihL0wsBXLOjxEDxTOLee2ZYr95SBgDC1tHeVDYiABzne
QfQXb+sQoBJaP13LwLcOz9kvwEbjNV6LMihSUHBFfDptypbBhEYBr6SSbanLfd2Zl8/HhNOIdIlZ
siZ7EBI/MFwSMGpw3J/DVHrq297yJiPp2xZHpEoxMNxQAoukQLQTpCaZx/m50TWk6IHOr8/AN6HA
jzPYLS9Wwzfrw8H9VYiOMcB50FBeWbYELcKQzppkiTdaBP74zPc89AaaKxUc9lOK7VyJKP4czFEA
2tmK9V3SSv5tJWjVyVsIDnc41OtSVLNydPQOt5dCEJNQsDsxNyS6mvHxZZxtwTDkgQW1SXayzgw/
itPzdyGVsQ39maqAlGKx1wLJuOAoCIusyicngrAtzERvJ3/7cREufNmbelQgP9xQyocoLTXs+dtl
0ibINeyte+HxVxWmWZ2wPLlTiMwPOr/Zez+CuG5Q6A4c+AlSjygoLqnHGS/ShrcdQT3kKVSv7A0+
f0VNyW66tN+zq7exWo8PuhzgIwhUZziEyV0gGCsVfkYHRU7zkRbhlI+tkVcIzy4Qczc5rcR4UUEW
NIJlir/yzii+uX7gOVYiV6Z2DUeP4R1F+JzM4LC2y0iagMlMfL4xJ3QQYKPWmAsM4VYrQuQRksOU
XR3sqU1aQXA48BelK7sXMep7rxslQdTMeYRFSGKjBGXeqGnxJtINrDd21MvHL8ZtF7obyT4mewHe
O/bquViBVzEyrynuM/Aylhl3o10EkR+ncQqLsaPZk8TwoxC+6CNh0+Z2ud2ry8SJ7T+D9bzHT85/
57/tnbeAxbmYTs/ifPvLdDu9wTmge3R1ZSZCySsTS/Iaq9rACWcdU5BTBVEFEZCdyzjDP99yNupr
+HTQhtnAB4qibEjiU5QJ8z6nYRKeJchPY46lftAcshXDSDjoN/evmictNUGGMhi9rRPz75UBv1xF
dWOxjFp36TkM8x8V/Z3YSX5pkE5VV1GR0rR7AeC07444Yo4Ihms0S1sY5hIqBV9mcKBBoLpOnBxF
zPQEeKjfNlAv5FYUZaWWeNdrsz9JzIRdsMbplqc2bXFh0wx8W9934cj9Us0qhyPle6TrvwywruQr
JgQ1xKMz4tkP7kHPyD1AwtGFoDl63jRUNUjG5CkX53lWbM42eJ6850SD+3wKJOG47Fzg2IBPHlPp
qMkfQyKZyAPUCvq1kF5+vetr93oKBgxjjRukbcsjW5waO5E9tC57xJ33SYnqP9otGeKE4VQ++3+h
XKa3iQmRaXDYb77HHrYXOOk60KlZX88+BxufNlUPqpY0vqaCFXunzOHUDqJuRCX4KM7K0qNs6me3
lK1Yh4AvW7UaLSPOSefSIcHgKCTigyAt7IrhorSJq/R6TTkTny/hMz+5+AZmR7oMfgpUudzmA2ph
vJ0XT7NYnJv0Rs4vZvfNMgQ01urWvKZRArlCNd9fMd5c0rp4DwFZfwCkmjsHiPsIwIAJvotOzpP5
ZEWHU1v0NCOr5wNqPsFK0cKug2tAREoXiGqVxw9WdtujL6oJt8Gy5jYaaiZD9S1K/ijiHiIbAwl1
RhCJFGvYFyVQ021MvvhuuTVhG3ZQtk4b5I6ve5QCp4ACQJrlvkvCb77reiZycvkwXz+aT6EHGAa/
tDWwfsND3JV35+YKv7mtRTh9+POvpHfJX1profh1H/w7aFwSbXQR9hWpqjkrQA+E7V3sRcedarzE
poqHMW48kZUdIKZr17drLyVzcIFFguD3f3//drwxZYT/ZXklviTDkw7P0m3CWGcfLwzqnmBZo2w/
900F33Uu9addIxtrLsJ6mGfE0aXwr5+fRgLRJsHKG/Dufjq7lanAs7m8bN45uID9gKEylWXRZqTe
WAO9YtRKExpLwWCyA+lwAF9vXWJVGkpHxkkkI/zdMw5XeVpHMchojvhPXcTGGQpP+nvBW4CyLA2A
OIl9wl7c3OKOEIEq6VwmWUOXiw+eLSRdfHjrRIEO9C6PVOcYEX9x81jpIvUfufJZGhpZhiAKU0Jd
qWRCLoz8QnvEn2mw3SV4fsplOVTdkADsWdjq/zaweub7M3v767yRuFJ5lyhyJyDtwx/ySvE6QxpX
LndRUxPjdcq3AvF6lZ6gogNxJ1xHsn0rOdkX0RohhNHEDLSatw1kbBn3kLQxswFUXQAjc7Rew+Ol
w3mfBanDtXGPXcW84trQvpFqfogYyiWN0+vRTdYtLI6WacpqApyvKIu40pThm6ROHEykP4pnNODH
37Ck22kpd0RGInP0wKXc6YJSLY7BegkcNfT6W08IkpQMr66kfXlnHu09M/IznRsdRdo5BOj9UGYC
BXnmym8ZMDA2WgfRCts3gr5SM7M+aelIrKBrpj9VrvWF8ILcBcsQAXwSlQD40Zka3BwPwkG6x6Oo
VslgsMG02+zdWO6K1Q8YAVhaizzuXnXegzy9d50LMwb7H5060hjv6/on4wgpHgvdLY5YNVP0flzC
QDTG19ooQtb17JZLkOQCo0vtxGT9G2l8dXKsmhZAGEmFvlXwQkj6rVBxWSvlXcTjOrw8bJUaJLFJ
abIo8pvcB270vZYYMI2fsXnm4EnXyOk3g+fa1SheH4O0vo45cIqsihO57Q14vxje3nMAEC6vC2t1
47fq5E7+3G1eSno41Ai6kvqSPHLxg98VrsFtS8NNC104jLuJkX2Zz/8sSOhRreS51qB/7WM6IWv0
w44WIJJTUsYHFfaCmAijfy/LOTrXdfCFY62mo8bpAX5N3YCfYqrf5JDYJqZXNmea6FK8OufNQpT1
ZkTyRsWQKOwJj8GJCJt+LO0OaTE+Gx5fW593pG80ZMNa6goE4siD0hPuT17+OCbtCORE4hqZLoTw
EdjRKdo1I8wpWNqfgiWooJa4ZCRviJYWdGFu21bCobVcjI/Op3qFfJgNNrdgbHDmf3AWseOfcrj4
QlQ2UUa3Ga6jOSPTzMGge0V8Z+/YQIheI96fxVc24mWVlkimwgl5U1JZfutyHz2E0JXBQlr+YIBr
OHu+oi2Ub4RtXMuT3IOzkJHJIYY9yRaF9AEw0xpkRUq9jbBYeh8jhoVnEphUcGlFIgMLieu0gVkq
zC4XO2k61NwDm5oMJzGOYWxIH+1ovjTAtQ2flE0KnnzcQGgXnqBBxR1YO9aKEWHF4AuZUK0Dq5rL
q40eVND2RLeQESvoIsRx5CP6jRRzxiJ/SvbP2X0+QEcNHJJJa6fAj0OwP058k8IX2Eqo6kBcBX8G
DMr/Y1WCaS6Hk2eP2L01jFJydTAf7YecV2WmSKc2SWksguYf6KQUTthjlxTD+erv+ud/I44sLoJS
xbIqxPMN0r+Lj1IV0buMGFW1lUNgBV/DqgCjQB4RRXm/ALRUOAthr8shq7dk9vltfy9RlZAtHhIs
wBJWeQhv8hRyafRALFtu4OdPKi5tP40ysixGuj+JqhPpPkVLF9aRLBUoev7DxwyMzMU6q6uCRWK4
++vpslbngfSPr+WCkZDowIDxULS+DRMXOlK9MqjasI5waT/c2c+vbKM3k7FsCNf3CII9cWqwWu1g
/RfQRZVso0OwGb8nEnaIj8a1SMkPPbOZiOmkgDJs9hxi+PMtmoqVdW3zZfofbhjpZaczSobbAjt8
GfBA18b07aix6kuvyNh5W0hHx0U9jzGTkgN0nmUTEbQoBCn3Iu83+raFRNc349NVhAp4FCH6bDFR
arFM0LKpmSIH0f69V9kFKa7jAjsy+B/pKLIntOxbnTnfnGZfoyeGmAV/GNbw8g67VjDeVT0R/qFt
n2GYvA4D7tRCf+RkQaroQ1GSycl7chngi6H2/3QTuxNn6TlLRh9aWcPFU5DIezsUY/EKjcJVufnu
83wv0BL4MwGLefPT0SQT4fNvjrr1K6f9JK4oHx7VTi7pkPgDIQiGbddcqWCFYSEv17J0V2T4aRg9
+u0fD20jKW/R02guI1yPQgpoJGepwyW/Dw6FWacwtlq1Jpd5j+GKtFPEeQk2Cpr84WUym052xOId
hc74lM4tykPlHL6+JhvrRkIRxVaOjgrwgjmRXWGBjj5CicFsC3sjYIGq4JGiFfC/J2+8lG5sd9ub
/bIpCA+eyVh3RolHX/lH5nNmGt8Qx3aborg5pAwTnx7FQOmM9AC1Lsm2U12cS6l6FRNeA5lxK6Gn
AoMCwuXq7IeRGUHVvuDs5OO5cp6oA2mrCtnuTGe9FchVRpHi2M1ULK0SK0leXSgTJJ1z2nw6GzpH
BkGUW/cqkt7xGPRensJC4mARiPPWV6MCFcCGuxz89eyb+XNxbiWKSEhr8aKqWbtNRjoRr/it8Xt/
wzwQlxVn6Nsi3vWatgLXVR0rXADTpBi8PrNmwvGdteqY5ilVPTjMim3pdMMss5OdIh1/DUn74VgB
v5J2iRELQfp5OcQdPQHiOS6yy92rSYTtNUdECV8D3FHdRARE/7Ls7RZmm25hXWXHqUbuu3K7sJgn
qt5VNME9qHx9mwFpsvzVu0vlhJ6tHb6HjZKB2z/fHXjR0VCFWlsRpczmXlcKB/0GZif2I+zSS5NJ
aOuZmy829G4tSTD7L/yUNVToviqdGqWCmsGMqxNcCb8/JVCd/iF61zVjurLlYanWN76MvUeyjnbz
ouAcrktqXDGP6Mv7DOtVkJNcdPpmy0GOr4e6394j1MvETMoGpW0nm8Rh/5S4KLxZauxQH0YYRY2f
I+QIkjPf3cXVC9zque/zE+g3e7EQawAedGdU0XbfAJOQsRz0ezholamSINg3YosVVCWRT37GhS0I
AP6a2DFM6mAfP4FksQYEkv5FCtzeY+Ny2nGbtCgfAu3Qb7Y8pygVaaXKcRjixSb3/+PPu1vxX5Ls
C3QIWAX00mKggFiaUpaD4eN6QdnOGOoDBJAtNbfvfzwrAKkzF2vBVtwEg4B+yFz6XtrScG7BHpI+
aNZlIZsaCINa3uPcq80koLtcUxnM+ubrza/wkrikxPND/Xb5jcMdixcDu8a/ZubUYdNPGLt/lyoR
0CZ+JDiNSALJh9gYdY5tQQUuoQZLMYRDaDIx5mRYo+P8KIC2suCSi5ISNVFgSgWS+lr4uu76EgKp
Aokl+dFA7FxE3HsH5YqHTOCihStMdJQyWMVId/cLQnUNZn5QLL0ZNt6g/tKbShZu1MLEsOuP4hvm
0tiemPIFgV1tbRqyd3iNGHZV1NNMEnOw5y1EnbkpWF6CIYDDyL8FVKeTSfKnKlRRvIC1JRfmjYmO
Nl/2TVpLpc0B23WgnHvlnomB6tk9Sq6i8UougYRlwQUvZO10zU2vL2f9oN/8IsxGQf32dbDdaNGu
AuSODARnxHE6YWSAIynVZdJdlxiyjME2lfLnE0e4uc9f9iagSbOc1pknLVnJxgc8uCWTGj0Op7G2
fxhiHpskCzvxaeh167vjX6HXIYuSIvDF8JXBU6xggrL6Q8EMvYScijLCzy21Uril0k7aCBPUDYAF
J+4TCI/VGOyjLUyF7hT2ZbXBR26Bywj36AAEfDA0GGNuKAQ5vyjK+qdUSFHuG6VDxk4AYfojZdCt
pnRmXwox/EkGYBflW9K45fj9LVW8mRY92Qf6C7Ryth3LDXL2x4k/fS+GwFqSkLzxyggEFVc9DSjv
Puyb7nPlm54VI4abwkJnZtXv2zouwOjz15dO2WBJ88Oq2T+l18gwHNg7zxNiQGbnu0tVvdDMsTQU
HeebdAsNtdPKTa4adBpA4r1A/sBfo3o29Wg0SOgMWoy/ue/ZHmNT+Su+Y7PDb5GkpGj/uPAjb1uV
C3c6YOLV8wMBYdEoiFqchlM02LRJ2dzEGtpGr+0DcmCIX/OLovtb+EjpCFXoAXC4VeGAzebiVxf/
kokxr6zjtPt5hLwLhSooXnd9G+zhcylJjibVYUDxnBo2uA0V3K1U/iyrnMHw5EQl3RHJcgb190mr
bt083y3vHkUNvkwEdlK8ifb0/gWZH5iSIWVgQgG8rO/P00xMu7BRj7I0misDPBa+oXRjhK1RSfEx
HDtZz+vl+AL1gBHNgrkaQGc+FkDuh6bqj7zg/vwGgiB1I8uAp8LXHVhAqKRgJk+NedhovqQLllSY
QC9ZmzeCRicLFS0YPIIiAN/OEOKgrmOxBjwMu7P9+x5IBfEfJNR3uAIWBkb6JHxU8JQl3rbwkW2x
sZdJzZI5EVh+2W42bkbTTNNmwrGLAwSSezey1r6Ntuf/YJ9HPyTaCutkQRR+sw48kgG+J3YU66eQ
+CB55AzfS8XOOmZxnbzCLdnaoK76I1xYP9MXi7BNXvOVPYbgP/ayYiDUqi+e860CRbx9A7RH+1r8
YxH8OZ8ep60Isr7i/SfraOFTtCANMDpPI8G0zCuU0Me1kGe8wvjTaEKWcdJI7yxObHkGeCSK9HQ2
QAFh6/fMJlovng29rKjiQUEYX/J/x5TchUAAOdLaENo/iuPjSWHet4brPi+2P6mlzmGGufGbTHKQ
qCspUaO7tB38mddJQ3+XrNpagOSx9ZHsvbGyUx57ong+LFUYQC3pDsrQQqxAX84JSuf3xQXQFsjm
4uajMr+Et2qySON6Dp87LEhfJsW7PM2tQScjty7XNzaw1JtKWZkPBXxmL1NnfX8HYcBvHtE47GsN
KPpebg0oQW+IxmDZWy8OgbQw4bkpfQEI54wY/kN7JBWpGHMu097HKGgPM/6o+cA5m4q1IOx/W2kH
kwPUBcGYIcRxNE1xYdiOtbz057QEErokjtVjQfw+iQsBv0ZSpwtP/OR00TQsv+wNgh+rg0Zmaecl
IuoXNBuUgpaWzN7xzLEXT29BqBD/AozoTy85wfaSc5kE2hLhvf4IJO+CoO4PMDhGQ1EQ3xMJ53zh
IhKKfkZpd44e4ueYaigwu8TEl7zvCwuS9BiLuT2na1Zjp78jPDTUq4Jnx35OaFLiN+S8tpG+LI8N
kUw8FFkWyHHRulhU6cpsWy5LYRu+YjvKoKq1ACHGyFnkXNBz4HEa2eF+bcqdgDNXc7YoRAhvRYiq
fFRAjqm2st6MAMs78vSwsRif0WcQFV1PuTxTlGryPJAnALTIvjk6KCv7SmHgU83ew2G0XiZy3qQV
CWYXxhw+7HeKVxVkcBjFy345kkLvIL30o/jpi5hriEmWc4sP03jPctfohou7w/IVmeXMloqa4yav
gnW8fbEnpJwOvYxF1tLPD6XHMpVKvmEIQnATqOWJT+e1frNWYKOBE9SmXQH4KSszd2x0adgEScvI
WD6bMKIMEpcb4y4PnPEIQF4WrlnrdOMwYPeKYnPZ0uPTUOswPl1FFPt0evi02eAaFQxIrZmobQ7m
DQgOyI0KFrfTn7wG3xGzoxuotFzjIjf658fxbW8zzz22F5wVts4a1jUHSlWpXqU8YZesDruvkBgN
ovEmTr6CHMEJBGRgeyCajo/CD5f3K1xnPuDKngUPvrMLG/S8wIaRR632/9H4a4gS2VoKurYn2eC5
UeY6434UqaZfKt+XA5TlnphL2QD/+JmBc1N5/96Ry1WwLSm7UhboZS9y03j7mcCeARPnEsUO84nZ
yJOwNZ2i2+JOJJBjmtu2U/U19JwyspXrdu5e7adxD9vd8bmYENb0FVFiOCq6PIKmpETjyhd3wlVS
FGWDnlDNgiFk0oTLfFlPix+CMhTLJl745tSUT+RuCbyRuzKGzGSDYex9TZy3HQkvJOtGfUzLctCU
CHNTQLogFxC6XxRozwYgHnKNYRdJgJhrEFh0l1pW28j75HaHft4dHbxxl+0JkEASUrYYroYYFWAW
mv6Dj8wWzITmNz4k0GPM8UYxksKVmu/7xWiaN0MAlLsQWliRFMRTzJ10LOJ/SsOeWhqucrmATYWn
XrhjYoSfvjJcmjkOLeMEMqenvOTKAM2DNhU2OcfLzNyU8ck+YLhE6EcyU1CImkn+YCM3QPLB0/Hx
HcUhvBMmZb0rM47tb5SU1L2hRhqxnxntrcj9dv2kKl2C3bS3DGLC4AupjjZHL3O9SQoN6sTjFNZs
W5O1ARISG6kvno0bayjmVIBo09h70VEi9Qn8vcpDgZTnKOo7er/PcL6WleLT7pxhBrQs6/tBeR4R
dP3+ffkGRZjjNanK4CxJR79Em43CgZ1BcAyVBPlF1i7ubJf5R5sZBLFj4jxGQEyUcv4uty9hKIfu
oZYk1ZAPxmBGuWV1rCjKaHON0MiwA/G5Pde+G1418WBZ4uoP6NmOoty6MoSe4oYMbWQ/lV5ue3H9
dUyof1FasKI8JylhCtRvJ5JePztI24OZHfwJoml95ocapRaWzyVIhh3Xh63Zb/e4hk4woE7Cd8B/
mwaqjPMJ5xoioGkk3uHNiC0iibCSUGezrIa42U+j41sNIboapqul+j6Lkxaf5ICpDKUlWSFAo/gq
/KClPwLLGPH+5uIvCheTz1uOcOfhiZBlsfmFd7caOJ3gxwwWpHAfLFEnq/BRd1FRvI5pZS13uWyL
q4+xq20GVMxXpkaP5WZ8G4H6OO9r3hIC897PDzdLiLu6Na6u7jvVjipsMDFX+LGbdSoeH/UNQTAt
jwarnKqUq8nlvPvbVjrQWHSshZnKsJJ3gjoKoGbGFiEy0pk0SLTALjtYN/slh8N+H9+mUSyO3ci8
6cbsG0AR0PLdVJ375eb9CpZVHOsTSdCHwtAXcJi/zuvw38EBkZCS7Np3HhKiKMxDXG1HtLe4LKjj
/DxWtsixHnBf7GkGDyns7y96SM7HHiua89PcvCdR6iWto7Qex176rgzeamozEPucORUmjEh4NOZ3
f1weevO4TKg0SzSV9t7uTd7fWgElVb/C0JdB3MrroscWKfWYbubrEynmmAJiDkB/vtqrTJWEQ34B
hHLudpXuHPCoPcdOBKaiyP4hDcH9Vge1qTK8L0EUcECyGLJl7tXmfVxtzrsNxGmp3hW2NHBBT0+D
QmWpRMztv1BApkH1Y0WDAst9NeZo8XRKcaDpyjKCx3c/yKtPPNg6e1qO/qsKOqxZspfvSKYf+3wq
84D9I7wHsUcnmuHJJdPFqFhzY83PxEtYpwUizc1GcNd0zp1ohk8VCfYz0jOJ6IJwlqEPZKtGwcz8
aT4P9+zOkOfYnSKSVSnASl16msnn1eGqx3iilHZcSn2BEcGDXKiLzNbxBEGdc2T5np1FiSBRIq9p
AhUqynb1Ulw7oJxB4ArHTPbnTyymcO3OdpsPwcD1DJ3iYlUszIX5Wi65rdW54otjTueKrAVkWp2Z
DsGJKqefhuAKrJc41GFUr89oPqg1IcIG6R0t1FC1Wpg4yqe3yWbti1e4eHZC9kakA8gUBX1dQi/1
wkETpunF3XwcapWxXtev/BMjSsU2lt4autqng+VB7+z49Yz+xWpROMCPUmt54FoxA0xJHrnivxOh
FJk30VeM+BqWqvdlAPiRluOhbkyrWKL+haw71PgjP5UY/I5iHAcD7XvjzHxcrLIxXRbi01oorM5Q
8Bqky/vD1Sa5HqqTRuL1qOzmHzL/Y5v/xArrKzV83tRTdx8dEFVd0m01Z4jRgZIuo20sil3jwuu/
fPrJOEgZpDs/C6nEjd/Er15yE9O77U1B55eJtiwgGudV9XmSPYrHtHM1A/B/v2OTNOzvnrK2V8IG
EBgLTGcguJitIXwHnYoHw7uTYfiHtXebSoO7CpdAQqXRVlUTOvihj3abzs9ONqA2WiSDroVK4e9k
yTR++OEuT1VEaIkEGJz6yebsvKEwTOuwUn7G++QtQn1kdeEZa7Png8FHmX5QN10TEkIda46xBmyI
VdJSA9s5KMJjlwHxq/AGFzQBBK6/oApYLaxdlYf/1KE9hVQ9K/ynY/vHg7PXAVL5eYmDiyuvTCNn
/KLuluONvJjf1zpNf1GuRL9lDsD1aLskkrD/sSeFlJg+GvrtSWHm4QVXLB69ZC4bzpU8H5aqRqty
pLA3MpmPuU06ujCv5mm9c4pVZjaroTA/Xz9O6rTgHYmwkcUDImi74EwHLXmGgf1cA3MgsxAe14cV
3hSEqX9k5x55B62isJX+jh9nhPzUGj9YVvWyCBVuF75J2a8lzkaKNKC3eST+HnxhStnLnSXgM3r8
qDr0tChb5MwBJODpzh95plR7zm2I9LkBW8FyGKYhYhicYo+oVJDEB8WDrRPsXeXRzVIygqj6AwYq
VuAhW7salyl3zvSPy+4G6sneHGetU1cRgQd7BaA2GegWkEVBpXaG9L7Gm8uSZrz6zB/Q9qC4tZ51
0T7sy7d0FyDauYKTX+owKoDb1/91Nk0oEcKaqqBVF+OJPsR9GIoHVK8Q714hvcSKMvmZw4d5xiA3
sze3TJBMJyZuKo5qRjVU9GMmjYgZxnPxqyApkPJboXql/QSxlwfc6yFg8TPT3EzACJJlyTGaeKqe
hu7iS2wEY6YZkfG6649NU4e+LnRrUbvLx2b4MZ+NxSiRiyj0TkbyMK3F9VpDIDOIDyfCo1+HNpWM
iFVEh3l5IOv0dyMQoHAWwk5ICHhEQp5qcD6iitF6WSXtnpIbkJjjd2QsIg+1Cq1t+2sSyj1cFePP
TroCw894baFO9+ddFF3gLMMOu2taXXThAMIsAUsTEsjBda343mvIbUyvRJcKb+N6If+qVYs0lnR7
M1+AK3Wpk8SSf/66B2QXg8nLdWrOgJQ2635BYLmbCTXpXUm7RfMc8bejzOMzyhj/sbzmpAh1jMLF
f6c9f/1HqiXFjXGfGIvw+4AFMyGIsNLjbGOkqGCz2ICjA7BJjMvjxIh3FJBuAZV/cPFBT+sI1HGE
ZreuyOdlmV9cqzZ2t2mntEiGNhw7op6aqScDy1MopPk3fYqZGyzBshqBflg0469gjsN69PdBIuMq
H4LpFFZDPLFwtW0Ic+pLsPzlWmiXxN+pr2QFEWG5lA00GOsEpZOLZpHLtI0NZBFQkVPOdwx5nP4H
JhmHOnRiE9y4qSD/wZIAXznhvEjnNyywmnyMsYsBCc0a7jeGltzkHUVGkJ8SXA1NDqE9NzEehK+h
I2zoLMtSXitrulZeLgAWRK05dDJYQGs9ISxd36rv4ZyNs2wIT430LlF8AAGswMjJMHDWSqFWNRut
Onu0AG8l8KxT4xU+RjSIdzE2PkQgGpo7ZdtRE5PJD9kRvw7Lox4+uSOwG7lEd1QE7vNoCOaHRrKJ
4Hiswq+iOqSbqFuw8fWFawh5uVvXV4K+GZlPnJTwbzr0Y/JN/0So65BzvOmrEINOhhme9UBRABm0
A+2ay0pq6fOfmW/pdVJ+YUcV3vEmrUCKu3rFZMlNtRyLKh7HA7DZhMzvVgp9Ian4nRAKO2tKveRd
6Q9KTf04lmJteGwl7jnf/b/deLNGg749OBHwANqjg8c+bnEDKVVNGnnXDB8J50E9eYajEkCnimbo
AzXatMHA4kGD63PyyPf9Dt2Z9AWL13xQOyIq3AipXNohEZyu8Hqrn9pCBc19njhlCvzS7UXKfLo+
voWjVFRBrSi0cgZzs+bgxnYYIjqoGEdME/nnBHpBcIIgzljh49QncNIt9QWW7KMUdDFfSkFwWpQK
St6Wv28AHeONgk1a+DT/Cw6SaZpjGuftXcNoCLftXSpcDVl4s2XkXPj51zsRKw6SnnLjdZMfw8Hb
HbmHM+5udP/Tm+cf/gdgWR67a7BI03lnD2aFTi2l5vFjfQQfB7Bk42XvgfJNrt3b0VrOth3NT+5q
5+Je6y4ivwK8ABUXcad9lk9DMHqHP1DSK9fzyuU3sE/ftPsZwhilF8ufcv/AJYpb29R+ODuj+ffw
rP6LuYVJQjKBUsPB1D8REXfCSRGnbxOOjw8kC4mS3bBnymANO9WURYo3PqIHRMEMsEP+GHTLX6V8
gLpwcYDftoxMGa9oCupEX/FxJw0iNeThLPaUlMCtY20eSAgqUkG+6VbZ9E3IcNZ6wb4kHiP/CD3n
dLJCvJsyui1uMjm14IX5TUqcscrHZLU7dCQQWXDy19AaDLNYA4To0AoskLxY60TlCK7j6lKoKgri
zkrFyc+ICxpT9G2gFHxzxh76HvnUxIc66oW16EBsbaB1fGmLR+NiKtpcS6FMYD5lkYbS1EwQJhca
blJWzkE2SLVbczE6iTIDrMvH0P5rJIyy3drvCTnmVgIKqbELVApHrGpqoydjxptZYMQBHYwjVKX0
4SSUrRVS1F4DKL6nGR95oAusucjfADx8BEZlgPUcr+dgcG24zxiY/cbxDSI13jhN0JGhuR81auMm
+ObnVOiZTVrlyCLMYGn2+zDq9fsjVamOc82rLnEFPNuXHH66DrLP6fqvumzy1f/grpAAXzbFozl2
oPzuXIGxpJA94v8lZmQ8X3k1BqcLzm6QvCG+x3iYiCUmToq6AG7yk/1pwnb4q5jeUNayUY2P21Vu
/ZVZTTSAc5qAVdTsD7LfqmLHfGGc3GhzgvxwopWuJ67nWf3Q9eSeD/0Z0LLUIzXhEZ7fJrgOB2m7
8VIIrWTQ0uErGTfmQgiT1rI/C0PIHmbSSv80RLS1J/iDhG8tcB98b9h0KQfjQjzaKp0gEQwAyzTl
zISE1lqgvw6HuajG/VQSwFYCYKjkzEAf73gIfJBq8OOoMyu8l2t0EWHvj74jTnCOLMWATYWW89So
raFtTwTcMPF6ZdZRME4jktjHgguDpgHaS60LU2Q2YccWl0dvDwBCk2SA8qt9gLE0B5s+KyqXTQZS
wQDXHmKn9FoKtTqSx+aBlaJ4bjI2J5EuhWcyDOBC9tT+G4rEmi40AyxsiULSzXcfOgROTKS6WcBB
AtdLsqHJlcLAEwum5Q2z63YMj5P6XQyqVf+UJ7ybqEcnDhNelQ8BSEfulhOyWzKcBBaf6yTVZMOo
QbALLwBneAsOynoj5lmIO/n5FeuDNAiFMy1rk+y3yu7eC5kzWWB8L3S5zylTP1SIgCOesvbMiZOv
S7+Q0Nd0SV92x17r2T4ZVuh9F9fA+b87dxiuZNe3yjUWzTEUPAUqc6r5FSEcitp1facv9QKqiRjP
7ZAa9K1UqCn68hYvw6yoBT3whKc3FGO6SwjSBkRqBTnJGBdyVBP11MfI6bcq52xFnh7tg4GUJ7TV
vike6gLN8kZfAOagZVhJieHyKE/fWesdRcAHWCiYpJRM9k2LWGqvoiA44QjclfndEmyvqrQO4X3f
5vlzdSWIGf1jevkFLaDfeWyxj/ItqQHkorvJsCf9Vah5EnxIAmUfrLewNa9+ujr7NSE0dszHRFDM
ehI7mQSkFczMthLSG0TGAc0FQEi54ck4AkAY4+0vS7nPSjP72f8XMBBZZJkzYzGfcMzaWHfHVxdo
xr8x2BtW5WlbwwGWl7xkso8BC1rDkzQJRUKlTcxf+thcM82jmMgmWNPzrDo/arnw1KfUPgL12rMy
1o72Z5kVQd2FPDegsD0YJMXt82xEsA25sjs0nKDG6qrJF9bb/xDKifBhh7Kd2G2EEfK44lrIJ8NI
aYwio2TnVJeDpOv/0h0M3UtHjGGok32HCd1lXLsPZOFYBqjdFLfriibjvDoLcDb797hmiMJhwjPM
5+UlZIInt8jMVy9/Xj+I6ruo6OKlw9SG5qoMDA2QDco09RtfbZgKWpRiowavxgLhrtXOIjktm31t
aqQPu5/GwBKP7TaJbjdvdsK+WbN6kb4/VPlbckKHDWnBO/Ng+sC5+pB3iB41gSV+2gOyRapFJ+0P
3yAYlY9lSlEQLQkdGJvcakzI2e7iLjDMAxYnmYWjbNlA0ZXATcCy4+deTrn8cgKf0OWSn+onayos
NQyhZiXZybzNjtwAEROlOLIysttjXeJXoCkB/tTixg0LJ/z/1j9QyyOVXdAqEvv9D5EuiALeg3Hi
xgH/vSXrFbVNMV2l9L+BOaCHia+hMkqtTJVDMfjvNIO/PHdVgi4P0Ujiqt84YgUvV0gg4qRVvx1Y
Gmn0mKt9QlFtx850vaoWsDF2xxSAGZPh83CA1EdWEcJZraJ9/2683TUntttxsK480qo8EyckrjvQ
QnvrAoGEHFwcTtKS1fxcN9NKMiNDOlwmRHfyLDJ8HNhK8DXfUm9F3xJO3G9n2iE+U3h7z05D8/2A
yAy/Gv3R6PDxF9a1FNwOy+5xVRAj7gJT1DeivNFk8X7KwUoofH/yAuU5GKrZM3KDvVJdf62e9DOB
Wrl6jfZRtn0yyjl/Qlujl3N5H6XiNBtR/l6kTl5DEbZBhBLWD/MFmVuOl6UN1xxMEF0Dbg6g94jg
QTax6ZOxhbA1utQ9tiNZSeKc43rSVPB9/U2wBN4gdPDLSdDWdsIXdNUCZRFRxaRGbDe2x2ulmV9o
4+WAyWDpD0vlrT8lorNlTUWabZlRMsg0GTZZIRIsJZGbVMq52Ol688fzb87/bXyYJ5MgAoBS9e/L
TtoZ4itxfy2RzEQhlRgvB3LXTnextiOKzlitmY8LASzrKDJ7YoO9vsMGkyeh7CJ5eoq/O9e1WvOS
IJBCjYh/efppSYOVoZ4ajQXkNvSwEexzGZPhhHJ/PZGtbpkQ7EsDDJosKruSpW90VQ6KOTRpu5iz
ZWMrt8pRwuM92mGY2fiaU+OkA3MpV4v5Omxybj0l5oyMe1/zU+4ta5/V16XrWRWAPjWntdMzA8XG
Vz04El/bnoimvA08m/5ciSyZdNC0rm5MMkJ9vPQ4OPyqOXgtP0H/gc8+L3vSshFQHUPqpZdnUJJX
oKS/ZFPi/bcnnVFaRx/G1lffU6jl/l3Mnxocq2eE1fSwuwGZ3ZkFyEq0TPkw8woqXw6ova7RDCNO
7Lsk0UjCxg9YQSDxnipWYTGrIKA5Uc9Htomq4a/FwpiTkay/9jMGVnsjmvDOvoP+9fAIZIOeB71b
tAq1W0oUXVhr3w00vvSs6kSI01S/UQqqAU3Nk2XoFgitFNxUrS52fA11cse8vBZv8ZysKFyyL+zL
dM7wAmO5aUa0KaFsP5YwN0G1MFuEdTiU5UqxpFwucmzbKlwvBfh8ICmCZjg94uA2vRp1EKLifP0r
6g2JZzFCR5fhEHD3wtuASdyNeTXcdz2CTTNRwePnPgghcmYErMyf0W5Y5H7FZZCSHvHqzbjBhT4f
a5NaYphS4+m57lkpL+yL2Qih9gumfmDhpI6I49o7/2k8A9j1R6IMnqd3QHeYB5u5OqhpFyyzNlti
4fgoK5PPz5L+/Yse6lcuSjpS2Yfyg+zJ6hOosWw+iGy1eEe5asJGlnMjnTbK4A3VN+7q1KEyIPtN
zGp3OuRPenmSxKmKDdoasY2VTQxwv6ivsNer62Gcdd6pmEABkLrjAUyaRh3Hdj4cT269sqrYlDdT
rBnLd5igucJpDUIXXn/UgtzWx6y+O2G6nYPsaw0FjUTG1tYTkPv2Y0yJNA9atz06+e6JK2CRcM/x
vgPU+/EM4TfZX3H0xMvAy2BLU0MmhwDAHxW+sy+kaw75SPM1wl1YR+CaCpfNijWXvi6veA7eL7+N
z15t7GEHa5z7oo0wOB/Pr7RQ0LNpCk3M7VxzTdFBwsrd6mKWX02vcZZJmqGBesgw6xAFL2Pn+9f+
2AqJoTkR63hZjf3r60IIhUWdiWUJxg96OOmbd9WC0mpoapdLoqGvjE78laUqWnlsEbXt6Bp1T0wg
vMe3M9EJ+B79tGfT5y+WM3niUP+PS36a7rXr+PddYuS02lXFfgEI7HNuV2r+9ztMxHWnXFAmGLdi
WzYZPgXPGYqu6OfRLPFgQv54raW3kIaKTNryDwjyebG6TNLEDST4qmOAZtqlPCxrtjhWaHPtjDqu
95XL988EDS/wtqliyNouxvPjL3Q6Pk3KtpvRSwCIPcfKSHZxcjQr5UJhT3oJrGQTQ7wFBv1rxmoW
cH19TPE4EDE2LcJzCOz0Ekb9+NpncODmalcV/71iwr31fDp+ZlB8Sy7YyE1u6/b1+J23XQfEcHVJ
wj86ACZc6a9EMBTwsnKOr1hGihFBSIhcC6p3dD4755MpJiVyqWBs22o5IJ8+XGbIc5D2LhI3R5Ox
hMLnVDuCTZF0k7/ocHe3VsqgT1Ov2eC8GS324F3EC9AU/8VSC180QG0OjOlHw/y3whfadzPXXBEK
6CKvHrcAflxeS9ODk0t0komqst4SbJDpwLxdK4qlkZA8TFz57iB0js4rNupC4ELyZRy5Zh4+P5hk
VHw63Oho/bK/Ce221tvpKeXBD90LFkbpMj2TVlyDCOVTHdPA4SG6E7Z3Tka0Gb3GdEVARE3rzm4I
6WhiTudyVUsdIV+MMoj741Xg0LZ53gPSYLu6CQzCV0I/JSU/78y/N3vLy7mLlSh51zDv2Rr6hmbt
xHwblqxmaMsFMmPeDYLDvM9vW3HgDqKz27919K5VCoU2udJ9HLQj4ZuYEfZ9AGnL5uWlV4Scad3m
eGbRlE6XBufR5jHhCxTS/JAZHy2I5JTOFXz6UBbXWgY7U1dszIJ/M8LNXwQsEeQMfIZ9dqKNtty3
DWCEAHR8UvH38SaoeKatqvXCC9AkdhOQmiRhJeP0/AFXyMBTNue/PGgyoRHclxMEFHpgoSjwSXYn
L+O2MwZZQoFxfHk9BTyTrA6aYrzoaAL0bvrN1ITG6OOpKyi+FulrEpWX6ly3l4JggN7AdGXKjpjz
cV0vwUYh/gvIzoEbLYqIeZxT1fCdwpd3ZPPP3rkke2FIfK2lEgtFj/Y3Oh8UitBNsYSsASzSUbYF
Iqk8Z5jckKnib121N8byoCnxHYhF4WmeIaE17CdShQ3yjlTAD+ctB7dPYBX0PjKfnkQJOCOKCfBL
N8MiRtZw0HQNT5oGOZeF6owprH1iAi8CkrDf2c1VPwnOuL6i4iADwvn+DnICvKEO5UttjzRxzfJE
TeAmNv5eAbq8cFU/Mrl7UxrRyN8E25LUbqP08qnbnrxZ5qInEfRm+2OhnH91D1Qwk9DAWJZDoLgO
mjB2CFDwymZzcn4pZEfa2VVm434wz2bRXp7LEJ7evNgNI0OaW5fdClnb6ZlJNmY9CaUxhXFjJVL6
sizPzJq2apo64gcaUigaD/i1XSwuLk3WrU9ZwpgFmdH+XjG7MVCd39g49CUveuEQ9vNr2bzhEG89
7yEJb2+9BVg9RP7z5Sgnj6b4jTaJA/1XDHucY4ilFIyrch3k8RiJfRA4o3ErqwPXL/FAzHP15A43
sABSnlElgo537poLghklLWmVEwKYc7VPgQJbhCvhHwMGyxApXJ1OMQfJevsp1Rebw3fz3AYzz9hj
tM/WJ6YCaUPpSd/hh0Z5YwgDL6J7JOeznuF1IILQaAGYGBEKC7fuviu+sqpsyqa/VBj7jNMM2qbu
+4UiVJXCZYt6rDo+c+8bYENaCS6sJ9YEfwQF0tr5iDlgrViCTEcjImLnzTRUW1Zm0SI52o0v/1Gc
vhIYpLO9mtxk4iCltf6WWQ/V2IFiRUOHm2nwooeqXFdZqagnOiaqfBnLNrWOxsOAsxH5GyvqH9L9
a3v+0SsjOIPhqXb7vGEAg1S9eUwsbOkdsymAkunwxobuX6SNNL2RQnNrbYpfPgCzoKcrSxH3XaKB
qXxBUA3i8dV1/AAOjVjwwPSu0whjAvPB93NYDT094DNMOskeu5K1GH/AccZveVnZQxw1uRuanDKD
m6a1kec8i+mk/OxzlbKcXr4pvzncXhS9f3gPUDqlvlcdnlCo9h6bOS0UgmiPraqZB4VMOqcxqCqQ
xNtvblbfehdbrQpWlRrmfqqIlFo7g0QRUAG+V/SXTJEjMwauwnChvGhC0lgrah5frrF9YFKfxqyj
KEr9y6IQR4FqKvatcS2xqOYrsYLijQ7GyhW83iZowXZKXXqh+WqgMzcPltEgRrNp0QLEZzk2objt
prOKZFT8RkOdnr3eyEOeJMWH3VuV9UQGOPhlYp9H3B3xkzVhyI09+GnxYwHuAkoTsxAQuzrNbW0J
ECbGgHsm26E9FVjYPg3pSbGCuL6LTpCYMLPDOTa5ejnTskYOLraCj3RV67K888Dsu2XpHQXj4EF5
8dyLJl+Cs/OA9Qb19ucLwa0MEEXq9R7FvlESwWM7iE2cPyprpHHMpoDNX00eAhocYyiCmpB4PLeX
UkTd5ug7UVA0C4/zausMaBFbbfKeH0LuZkiBaH2xNjquoPrUm2uNH2Oi49hdWj2+g62JzE1pODv+
FIBpP+p755dEtHI8sN4Ck4J4jM+FYnU76BZw4aiEvMI5OOewxbwOnF9lo8I9ngKp22miePRCIFzk
bWHOTrDwgNQ/TpibcpNCP31rBzPN9W0hK5qSzLyd1zZDa14OO9cJdp7QG01XUeSVK2uXJ2RSDvjC
wZ0clNc1Ke5hmmNtlduGSAkbI4TdLdIxFPG3y+BM6bfarSbKY7B7vi/D0Z1Skg91aOUlSUDGbrzw
ISzdSDYThY7aEcBW0LLvApNT7jdwBRmIEG9jVBpLGpDKjGqd+2bDTPWwRZUXQnQ7lRBARUke/+h2
hQ8cjZDlSq/Z0KTd+gXcgmAK/dNbF2c1Tqz+U84jvyjF4YE0y4db5wAYWchSLtT7qWub5OeGYeKk
0t1VjoXAdz2pbtb3lhQ9/QNxdNE9Qe84dZe/f38MEENupQSN04KTXbC/zanBcPpLgCv6FYLOYoKc
oDoAIoS/+ZF7HzTTC8wQ9LhfWKemLZuYRd4wbyQDioQeXwuMfuxDy51GbyJUZ7jv559YrNvydbm0
xATJrzFtHmAl6+dFeNRRsm85iZQAkcAeozSbaz7BS7hgw24oH4KK3DKnz5SODkYbsCAxPRciSJSm
XYc1sAynXfSnJQeMx26UCMSM/LoM3uKKE5GTCo3rId9M8J5cEJO7ru0v8x3VDEq+w9qLbqHORaJ/
a68j3ejMO+bL3abgpfBdLV1zBLu7c4+n2gLMOhO6lxcISHg7zXp6jDyw6Xa4/Xd3driiMWYSfm5L
sppHgoqVOJBLLLm+jJorLKKhNKoBrjVuvnp/IPx6fldGZSpY00+7+5PPI1+ItUwOFSi/i7IACtQI
ekkKfJWzTjFS0HlFhnXzLKZL2sL2qcjA0HnF7d5UQDq3loC+AafYcGNBMnHve7b8savPdxEsqLzx
Td0X3xQo7u7psFEpkLj3mBI7ACr43LWNsSRPZ6xls2HpTQWLNM12BEQ/AscvnwYD8K5omUzprHp2
Wdzq6kYVKIlNjaHsgYir289YsrQYObmfRflERgynHx9TpDC9YxCOw1EVUpCMR2SLTvlSpX7Idr22
tiE9g7YavQe0+hytjw3+oXN6oLSMl/OhgKDtQiw75dng/r8S39zd12sm/gGclwqxekFIXNVaJK2I
3j4cj3ME0WXAbSVVGhxJkqbtzJpAbflB9j7wD5gHZ7I5yrExvzn1O0QSsXverhrqav6tn1D6VrAL
30Qj+ZRpFWaNto2sFirM6JqKwW0kR1LGDG1G+uMKb+phOZFE98cWlFAwAsK6P+W6C+tG/muF7axt
F1Ap8n2x3Rs7KnNvN6K8vkgA7ZC8rILK6hvuE1sZyl7kdY4dI5njn1h6+efGHN7yna0FzYtflzCA
/8vpIcU4jG38afmYDK6M1+2wPbIOh9V1/1JnRrNJD7oG2AfNMlV9oDCh7+Vgqz6AXR0uMKWX+19p
6OYxxP4mLPl9ErtWphFa78KvsOB/Hj8f2KABb0NnpQfr339SLc5AlUOFnD53Lg6OvmRrfvdzr+ZF
a6ewjLvIvcsDU5HYcFgz9c3CcBesn6aJhvNcq2z2MpaUKIs+iWvY5utfZSBweuGmF1VLsuEmUBf+
K3Lw0GxFlVMt0khbtKiKv9BPzWctIu0k2w5ZsuIp/TCw1fEw1b8L8cT3VT/t4L0XS5eCfmx0JQ+v
c/naKcc3ZbylG3X1ZCralV0SlJUXy0xXVvNVGLoRjZrjiuTEvJQodGlFVtrZo+9zxNhDuWWgV9zQ
uOPhAWTZnNw5IB15q1LWjGmcMOKh+TqvJ09NDJFIgQDkJt5Y42cdv/Dy00V47FG8yDrAGQieYSU+
eQBKNYZxXvQYXZzE/9uMT3L30a22jUECUi/rgG4l0xI2hL68WAmtsE7V7zk7h/ePvepdm72Fmr7l
lEtBe7eqdU7APijtAoPm1/MNbIXigcM+zep1RFazYz43noy23ifyl8NXQsahpCTr4s/nBRDpGK3m
i7fs8/bwSeJYC4+CAkS4+2ZyHqR6rIU4rMDpe3TadEenB8bmxHGUEKXRjauxaY10/Nq1bXzTqnDL
GROhTtgePqFEJFEEltAw23tmD0zK8gK2MEASd5UC9XtHy4dwsV1mDQtP2vma03B6qvJBNfTpLYAv
l21yvykKtiQ9bSvmCAhE1oicQ4DMigsTciFzVmlQ+xxFamlj40n5ozfEGmRN3QkrqupR01M6/uD5
D70fG24cuyiP44IPKzFCyvLoes6Dhnd0PLp+SASaFJQ32oxsXfWm3x4ubRqsgv6qeYiysJiqLPCf
4ApocvcpK1QujrJzvfDJNb9Al1fEWRE1vuQixqlUXxdMbjx+uP4BdNlcmih8/OibzYPCEoTfbSBs
7txUBMy4JwHLyGy4ZvH7y1WlNxoaE/qG3ue4SpK2ykqpSo0opDMxO2RAKT5ng+dEQYLhY7vKinnn
ECVK1EU8IA8TiD1mG2dlru6l3B+q2AigBPuYNuqBPakmzYZBIjj/WDsrVDA9FiYxoNY/MZ+Ojlka
9WOMuwNGFgj040R5bFlqH3W1vtuY9FTRPPuo4LjTAOzqR/JwOxSpStTEMIepDvL2EdMXeKFVmJdS
c6BYkuL34XKNQnXhZvp2ry6VCiYv3sjRDaElHjxK4v8AcHS++LhNzZVb/3xKWpIW5Qugr8xS2tZi
IssVTI7CmzY9byLkjRuaoeywfkIVKe0citCpdax3SaVokmlvDhLcd5oMB/q2cTvO+zn9LOc5UJj0
EnFji8fC0GDoP4TsRq9iyJy1/2cubDrzyN1FzaJQZz1Ao9A4mjxOT6YlBrUt6LoXIlVTZVi4QGnV
5jxBP6bctODWzzr6Wr4dn+IOoOed4hZi2XWtp/TQvxJJfyaaafP55snu9SJw9sSuP0w6E4e7i7mf
hZ8e6m9nArrjDgf0dy6w4O+JSQ6N/D7bdUClBnF75m89EfJk82kpnbDm9RyPDRS+IAlsY3MNYxI6
HXgQTRjE4kWloOfIa27BkPTOobmkPR1WEmvaz38Y5iQezvhnSFTO0dp9IKBydOqZLxhA9ATh2eAR
dlQG6MljEmDvZWOxoO+/xrJyxushkQ6j6QkAVx1BIkqNGMx6y0N2hf58xDK66ff5oy0g1jk3mRos
PqsYG1QwD96xB/f4GKwLVyIZ3YSH763CyGwstKTDhnsxh5OlWW6PPypQ9tqrcjc3klsK9/nDcXmo
zMhyaFhP17w0B7EWPVTJA+V/gf+HoGagxo6Z/iFks/eEYp0Vrg/pPPrjtYkve7ULlb8s6KoFTcxT
+h2MTvbHEnuN73D7LA9DODdoJ03+lScGH9Ljmmuy+RJL/yctgGpysR2778pDjozsPO2JAqHe9D8w
8LDyMktjks3ifSkA3RXGktx+N16gwH4Di6BvedrawJdzdmhKqNzwIFkoZWBFxapyGr3BF9A83Bl6
KRzB4+k2ZHssNI7A40G9Y09R/rLtZdMoek2q5sae5xSyj01jTQGvJjF0/p/7uZQMohZBmqODnkkt
DrYaQ1jW5tpWOJE7BpNoEsParN+wjk9J5HiSlJIZbBE+R/c595VVoAgP1gRdMHz0WlRVG24hM8a8
nKSfawOpjnWk9+gPE7lqDi6LEqe6mdjDvaTCJfY5tyby0qum+I6erX4yhnQq1uN5+aR4l/If+Qxd
fmqoMJduhqKDxE2g5+5pcKI8TLhFtOpsZw3nJFsH5BH7OsZk6Rw7eeQEAYMDhNLZvQubtsO7MN5s
baZCccdRjIDOyF4mbENjIZ5zzgXqjLfl5ZjRTudPmxA3+og0q/fnQTYFcIkSk3jBq2D5NWpVzTkp
aCPTsqhFZk65Gobez+Jlv9MJA8uUHoFPPSECkdPDZq6263cdjxSUUzI7hcq8jox40OIdNkhGF/M8
9aSNebbmfXgdsYBszwQU6qyscduVInJq06lzbyxQWnjNelA5JiQleLM7CYU7lUD7SmzUDapGy1wk
j77CyVvjLRaNhKSwT2wfMSGW5tZRYv6lmmqEs+L8Us324nXpXkYoOmZ0aTk5bOoEFFe3USfme/Ir
etoV1AKh+HI86qC/A90kgP2sJtbdrAgHfgx+Q4kKuyMdR3lWlAqGdLoqiU3Ng2Hvt2t/nyWEbn2v
X158snfSepheK/VSH9IOlr1RgJsDu6g7jfheJ7nH7TfEpRFM9OVNnUl0q1KfApZ8/7EClKUGMh/l
UkoQOSzggYwO9sifTtJ4jxwotDRtNkgW0jY8PEOEeiaTUKoS9Vb9BmRT9uCAlv5QpVxUihIdVQbv
WL86fFewthzIb9zsFER0/A5VUqTK/iikcVQ3cYhWIM6997PveFHC7prylHVfecWeywXS9UoIDf6Y
SlY5RG5MQ4bsctukXjdoKj3go8AuAnskTE6anT+scsgEUHczjdvwZ29699rRckQgKSlxHID4p8Xt
Ywg9kEwp1C0Ar6VltsSb6qe5bhnPqeLcd5wgbsQIHVWcXIvwm4lV4F1/QjEoTOUCtTfZ2tWEgXNx
QVHUlY0rOMNuanTTY0rviNO45LZSLJEmcVMsuwcEI66QJjf4ZBEL+HIhDwIwaUQHM5GsEi64HbS9
li5Hdob+aPRagQmkfnIBHOrCN13J8omyL8dx3wo2/ScI3YWSPgZYWZeA/vpraB1TT/+K4IHR1XAX
d0/XwwxRpWfMyejXj9FVA/MDJg+rDQbypfnweNMMdRx9jI41vza9yIsJN0T7d2neWp5OHmgpSS4i
KJ6bApWUTZXKm7D84dlMCORXSD7WWslaUJfUn9+eOtJYNY2qtJAgtWnR2t9AEf3HnMqAMToP/dZR
gWUASJK+YQuYG8mNG2JQDXGUR+bm+NkVn3qPnxYIlqDeLEilUtw3Sa2gnf71mJZpxcoWn2So9QlB
fmEzHMOEFsI9SltExi4AdLuPskf3cuZmpfUwX8olAuF6O9/YAZHPzcMEzcdWbK9dTrsRzyiA+8AX
ifTvuXK5IpukXD56mH5DAu1s2oGPvOhufNUJS0bnc1rzjjO1eA2LHfajahCkZdGMQmAtgqPlEjMq
wRV5v8OyUhlqwntlA4IVuER9u/sbmvGCKvVwwItlMTW1AwdJEAzJM/CVxr1iMDN+H3hVVa4MtmY0
gC0EgGYAB0obXTcqLniRSSX790Rrwcl/Rp1y2IUgq2itZUO0krDasAJIDTDLjea5VKkHReyvLzqx
nPuaLddqK8WyNVfNFhl1LxKUaOYyTDXPyHxsSSrezh59CpK9khpGpuavXy7dX2yjwcGyvunhxzIG
e1fiL4QPKs/5fiYUEcNXsMWDYF0yODUZTU9R+WYqiH9LNkdWJjJrAlyD7jIYuw/oKs3ceoq6zKsm
Sa5Hm1HE8EpC8szkyxtzzUoIKwwJOMo9B96ALGL9QTGj9064V6VMsBxTDnB7CgY4+BEbY+/uGQ6H
K7dvcBa0B/+8mb2ST7k3zEUTGXH3Mv55abH1hwgvLIovAAKJhgqy49dxWkwqgCNmm1AsUKqrqD/o
RlqkXmCvpeHoAKyeOqdn4qEEGy5UiIbcRtQbsjKCTH4e5kC1J1Y/YmP1fb4VtRREyb34KXruwyAy
8e2kDvoeRJ3Jo90g+tWL7Wh9Ztv2gcptWWC4+NpO1S7ZhlMczp1x6/z30OvmbN1ZyLv2/cn1rhl4
DwSwj8KwdIrDYBheBvkK8sGqp9AUsCYAceu3Ja9ksL+l6hOcd6XHb4ho6dkKr2JvzRKWubgbdfpU
ZCERl+lgHsbEObqSy6jZPrL0TzojEA33nIrX67Bm7TWVf+9Y5fx32QF4hcAqgi3lg1VoSLfjF/+P
WLDQIzAF/+y+2wsq8GGqTMT7g+uKjHsUmNobNZcDpbeeLbZzJcm1obz054bMg/18febTL469eE+N
8azb5HAkj3Y5JflNTXuopoA0JLNk76HCZ2w2noJ5KwS8n/YEvImkv3OA93/5O60icX6f/IFLl1FB
SdeX5Hu1v2Sf2Vg98kb3lRSJTiWpC9Enr63UQubR2WQ/r6HgQLo2p0g0dAWWYerVty18DdksNYpf
CDlRY9xyr6T9cKrdFfcTR17WHU/bnn11EmraQ6xOkrFrwj0rLP228wPjydv7OdW5tusJ3Ss1ISqd
x97I9h17EJ5rywWQrwk1Y4XeaZAXkk4BTw1Y0TVAKHzmbp/seojz68WaXmqSqnFowBQ1/OQu8TAz
fhou1K4B9YClNiy3KB20JOpoiMf9u/2YMer18bLoL0JEWHZ/V0P9SpeQG3bM+56mbMAbQP1TGtcY
Qhcl1zDJd6o6kzWSgu3FA4zSmzBCQ6cV+7AboDAdxXf2/em233J9LiMcokpVU44xSv8kB6mkx4uG
UpJwoIE/jKNmJ/5XQGlopxJyCS0ynFOi8FOsSQH+sEpB7LTX3RK72f6DDQ/dE7KDTxu6wz9Bim6G
irfPAR/PHZvXol9IVNDDYpJXqDhFSAA1zDrCVikiFgawFv5esUMGlnkAqHXk7xD629wCa+EWEyWy
E/iVSHO/iDJnUS/sEsIjfrdON89qGRz1SMSk+zFaG7R6Wigw0cus2Q8z8VuEjEwHtRzzm5MyE2jC
KfVsaoNwXnmLuHg30gYaFbWuEzwyPfDJjMbb1HlbMDx8L7U7ZhSiVkizi+2yLXGtMvDKYq+Y5DAz
4HJp9+i9MWgT1Mb3UIVRCHLPXcAVVzmCv3DwarqFgvGlE9Yi1g4PaRdTJldgqQEdYSTPLZ34iPFQ
UxXw3GzTbIaV1c6G2YreNB2gucjDfQevt4PMfqLAOi2FcUnP3veut42+Hxk9aacSX/OcbY/LG/x0
Cyjc2sxN4mFGPWfbsfu92rKskG34uKIaQfrCCzfT6BAWVX68l7j1HEyODdeJLIItdBhCypJIErMm
wG5PwC4oQdjKrG6sIte/1pVsyNIv+Fikg2ZneqX8g/Uk2WTuF/oWsO1xolU2UQTrQdXuUAYNVdzq
zx6MCJpoWsQOL7QrgxEnmp6NzIUOB80kLdM0M7PBOCmWyBNi2DJ2MQmw855eNtGnevBvBRS/iuS7
qM2u1r+avZNx2O5faOKYdo/Vjx5RC5Of1droJzCpdhUMrh086uguPG119cWqPCJzSMOexogEMy0x
av438/PchH3pOc0f8v9LJM7MYrI9WC/UJHMxH53X6I/GgJF3pUFNPRJ5c7Nq2UcaZFSJnmj5ezTE
48FE29cLFgoYQfl/xrcCKnVCp3Gdamha3CRk3txdmOG2pEgzG497o1BMz4+GqNJvFZXj3axiGAX0
LoPMU18yQWR6unKctTcHlZCuVDHT6gNO0lNj5o87WRwHeHa7KHk+RlJGl8X1sgyha4f5IT6g89U1
cearxhBUS3WFLuQVoGrGpYNH94xWvHTONlujNwkWXkgDNY3q+4SaDXaGsMVoatI/Wq/ynSz8ME8I
mTrLQWV3FTb2+SCj/BWZ17ayd8GJg150amh2iClsCg0iDHs6/G83ohVZMXs+JuB3fNXUQCvaoVmK
zo73d+aLZO1wgHOBwDVrDufmgKygtbroQESZfrFGqoGVGjlOYQO0YipaxTuhXPLo8ahbJ42QSl+F
0Q/qtupgS0bS5fkeKlXiCd81CgKFUlt34tadhwC9uO9qFjm0hgXfmeCY0eQySOd5z8VXymBRax+j
SUkpCBP/6UtZeiZ8H6eIA4dhft23KWFjbDbxDUaz7gz12pUJjZ73JGhymu8zP75//D2bK2KG6kuk
eC6TVdHU8DENXhlxINZIjcJ4+li9vkZ00WV9j1IdtdJqs/HYjFKKV5Avok3EMtj6nJ7ftI/ju5h+
l/NDCMsmOn7YTQuV3rROHpYNQonWswG6x/77518VF9NftvrUZ4H/sG/o2dC0mSohhRVvrnpGuIqH
YojWs3MVMThCyTfjmco3hVmJ1ZmhcQ2b0//eNJIpBjsbXvZ6Kn6fK/OEWPYwozaw43IGU31Vaw4m
zqGdJkcWIfSSzOy97P5pI9AspPBXi5Anv5kS0Ppa956mSTedO1EGHKRIBo0m7wnET06EAcK43jGv
dh0l8BAvzxRK5CmyGxV5hd+fhLYw+J9PyVLuAfWw52X+U8XlaeRJdMKiswHN2ekUWTevqsiWTlOs
F87JLwLznXlog/KkxBveF/QGpyjafciukDUbdSnLN1F/ztx8G/DNBM5q1uCzmY0xLpzk8kxIXfTP
d6Z+xgNs7jFgcdRbBEy/1XeaXnJMmzLdFgM7SH88yeW++u2jJclBb7TEb3dZ1CnN5noO30f8R3ve
6KoQHtqV6Y1xMDkGcQ79SXlscX3mWc7VPIVlkFwtZHlECEWA4cAtebh+3XIvvi1sIYl6DdVogDBS
aZ6HYpiP+2LUU0yBE1XA8QP9QVGModutPC2bNK2OTt5NPFBcyeWaw9m5ZPiTR17PnLtFVykp1g1b
vVQPbCOVKbbphih7EW6eq86gYasi6+u5eCEjnH/Iq/4yrnLx3JPWlz373IZ3lL6Idtmy44rBoriv
/M/pmZoQVqH0SQllaaYsh23H6MnZ4SA/BWwZTHsxakFiYwv8m/XqTq5N/CyX2zWaPMVYjdivk555
CIcePzZGzHBECwC3SBado/GAo65aA8otJRecs52PPvD15os3m8rvYMMjMgUIkuviwIEZJndHmcAP
rZwzFviQ+VlLmgv6QS7SkraBPJzwGTTjECK54s8TiDEKVj1aP7QNvZgm8Dec0qfS6+53tzyj3bQS
4xokgLYZ9030pMT4NTQBjcQ2rQs21sjRER92MSd1ST7kxFA7LxcTtwhOZwpuzWKMK23BYi8z6lQp
Y90+wG0qJ670PBF98gbKc752XRfudRmemqApdZi2c85wbtC0ET2tBy5EdXNkVZ3O3pQyW12bHm1x
Tj1cPCvnf4P2MiCy0IOuFDkWSkR5u2/Cl45Jrru2BnGybOqSzdBUbPUyWdrwHKK+4/TkfVkXQjyS
1Kr9PpEPp4IWgEGH/tDYybHg6MTCNgf1Z9nSZuYWfl7Gwxtm2dLr7wwevpynZ4vdipye9rkA/Y9s
zGblH0o6gXOiLgdz1f9ur0/bvcPcrfs+FAgnb2nrKoJoYlEJCqF6wCNuCL0IG97YQbkdtJUU0l88
BRQpUTaS3wbq7Ahb9Q4NHsvZ8V851k/Bn/I5T0lPZnkmFlhZdJff600lMWmkR4d6pwbvK4OZ91WP
NI7GNzFUkvEmQPzEV8uvytShtMXTSOoyfi9D0fk7/DcLo88J856qVlHcxbQpY3rtPxlbV29g5C9K
LMQ0D4rcRvoPFm8D/O5FIC6aG5wV3xjtOZO2UTP7+waN05gP4V83SLhdyn7PWdHvAI+0oAEXKtIy
pu2O8yP+smLkon5jsSid1w/pyMV4fAiQumqUqhXviZwKiwiElj6WmdU03QEN7ApHN8z4lt99/Atz
oX24j7U2qeFRRS0VakS5WiaQ9UDlsIJfR8E2v0emB+31/08RVC3uFE76OGeD6Md0pxS6B5lhFPbd
Ppw+owsd62rhpXGAxYlT03LNfA4YSdi7bRSTZGVeckDpppRcnLn2xHm7Ls0cXMie4Bln95cm2ZhL
wATZnbXCFuEZrufcMbwbCgfmW8gpggQPODq2L1sDu7KsEmtUt6/5STcVePvOCgA4omxolM1pAkMQ
okPa8K38QXz38+IiWeVWLfcX82Pxi1i15XSOAJK6lgQsvwfsWW8ljOEusH7EiewrbTOtEOe4aHti
3x7Evn9i7bHm7182863MIOtcugHzMOR9Vl66DYFcCmuR9Fomh+QP1KQTpnTfZzSh3wTHtjyIixyV
tG1aUwoU0POu0t5DRgtakOa4uv8+MCWjwSHGFf0eV4NMwOC3idzMlJ4Kv15+ZDl7x4YrUyfhpy+u
3y97R469GE2EL5tBxMIOqXzljfjaFdj6+nfzNKKYspZXMyVzdSFciTeHcFEYeo6nLVqEurYzQfLr
baOVU8qFmjSX7+Xi4fA2poULCrOQgMCVu3bHdyGTzSmvm7OoRzLgKdCrcEUCwc+ZE2PtMm1+gU0c
O0BWLOaa/JHzXAd3ixE3QNbmj1yB+7j5yeYP+t0pswAx1EAM+jVH/sPtwVUxb3WPyvqucEC7E2cw
Jwf06EgwR1JoJzALHiGk9I65IgIQsXnW3k7vBVMjgnYfE2JvRkps8vwK/C/geA7NwVed7pBW/gGu
2JniMcfapHtlGO8GrPZyfBasBI3K6nnK9CKDeA3HkVtCBa+IHonQwvTI2aWMdGtFHrruUeGj0yoQ
Z9nWoXff1DNtqLLUMdlZi8EJUWQkb/VwFKhkKPzsmA97Jvj1gFjK4i1Mn+Jtw9yLYSY2dGGZ5Qwg
J6fZuMcJC8GkmYB94I6FC7zDpaVOTmO5TxMv1gCtogZxVjG5SBnC3+mwXrJ9l86KNeu1mSrBdb6m
6pBv/fYilz4kT1NzZHF3CR3nVWP4D4tKP8d2blLbOq2BtZmjiQusSGstsRCYq/MSXTzRFExoGBo9
NrEzoze8lBJFP1awYpl5wEjzArH6flTHWTrqUYOhINuGYEoHm6hpY0OItp4b84zf3k/2Qf+Ueeo2
6PgasGkca3/okPJAa6auYwT+PNG5sQNtFp4uCL3nyYZ89svawpU4FhFcgjWoGhYPPKGK4Xf1jkK4
IsaKH8zZ8ji/NLlMWRclq//FJhWpxRFUR3IRYcCqcG08qtny428IGcFIw6ORf1ST8kG3RmDkhmAb
X9OROQC9ef80pPZpRNFNebbdrKxVC9ukc0ClOCH9CQrJh8INjxGidXxakdKESUzz2K23NHh5dkfY
0fQ5xjQT+wjEtZ5MrrnpbEC3ArwalDJ/kBmXsGGIyIMZw70hfQll1/AgoNuIdlzaXfKDgkD7IpZb
GrkSWSy/nl576hdPNUs5D5XPehB1CIX8k22vzYxAufMuGTU7Plau7u2+n1iU9d9gq9IKBZdP18w8
0vJxqmbd6B73A5NN3jq0tOfiktE8Q3eUvPZVcfTBnIUcu/tg5iIuyGzjWNaeBGh3z+cyJKjVUN+C
zES9MUnswzdXFaT2w2ipW7u2j6NARtB2qAtshg9R7Q/W6qUvux3AOxNh4iK6+AmooOQCeAKwDef9
CrAFWw39ZTG4b5Jeq66ZF45R0y99wq6h70Fr1xNg4o+4sODcIUllRjZCUp2hk9SnHnGvYphQrGfy
QR1hBQ3/rndV9axkZ00qTzjCB3/TW4dwjJbmUPowUgq6H3zcADuRCCwhBq6GsT1KfFPqGAE2d3lV
Fik7D8XB9GMfwWQsDZpvkkP7zL36O8cMiQH9RGadt+PFWdtaMQ+0S+7/oIXsgc3pu4k7AjvRqneO
mWcF7LSmd5BMsAKmsNtuIx4yW6TGRwKcNnC78cXb54l5Rhi6khq70aw/2fwgZRWDMh8nRfksDsYa
LoKxTU64OIJdavKFNaEwILUx6G9f79SjKufLblgcNYmq0zbwSzk13EIi0oNK/N5NZiniZjKi0OFE
s+3dAC0sfbMBszpxz9PfiGtPBMV7vEBrIgCnTGd0gvMz9HbpvoyDJ30OwEe/xeFAJkGm5TdaQIuE
mOoBuOluDnm+HnNN0Vq/iSYzHjMxPJWtmJUGnUJTnXNrO122l5eS3v5+S1lStlx5GA8/mY/usEzI
7+3EfIjoSAfVQdDJcpRrxUmMc/fPvpF87AABjuCZmtkp+24ICDGeWQ1Ja0hyDPz431tP/Oi5TuRD
jH1wmDkzpJisF85d7TZq5A9T/8kAKaZ1SK01RUa/BGZhGXti2lUm58XjnJ3/0HuAEpTBzMRjTFpu
q/1hU+RM3FooKnaYFi+ShWG/RWDaNCZp83XdtF71WLaNjl5jZNASczhDt1EAbCTWJU2azCYuum8g
BZub38FqdkxjECZqs8Pv7U2rTCdbTUQSs6MFj0zD/UpMsOzXckoJHtbFMZd95Gy9EqG3lxbCzOL+
b/4t0ZkinooQJ1rXc8Yeo484m/Kgpvfil6iFg7vRQkqyzW42Z8I1CbFyO4AeFs5jiL/XhYbroeJ0
f8Q9g4BSX+zEdf+BTeRMmuKoXSv0wWtr8qJepbzq+0kaGsi4y7VQEP0bCVaEnbyD3Zan/hkS2/Nb
JNMKpkAT5s82atjghGOEFHZaGBzoM0qyEkwcFrJAQ4IKw27gh6QywVn0BS05wyY9wOjbj1b9KlZS
A28WMiHuryeVrbwf9g7yTMjGOX+4QGgU9UTPG9F6rEoNkkkVwyEYLFENkXRVQfsNLBJU28Ja9UOZ
iUXIxbsKlAACEKZNn5qZ0QWGO8Dc5iVMmICPELV3bzyCNOsmvrFu+WCqZG1h9eZtrh2RLDi0/RQb
SzVE+dgsCqK1DJ0HhbNlxXuwI8tNTwcbFEZQauyJZI8DsCSNLzyNqdLHZ5jmEVRPBuVYLRPW7JEx
Q3VFjE09D9NxYQcKx2vwlnIASjhX7PxICDegAg7Y+SOEnJx3+Mc16zhIsg43qmdczkQMFNLrYEcZ
pIaIjY0+B48TK9g6IV9hmjzA3fll6ZewT2fLuXQz6JtyYZ+5guYWQEsI1kPy18E09zIHxnafuCIZ
N3BMQ6DaILx1JzXJ8rDttizO2BSNSHYValzHAPLUiSBqp3wigjIRGEOgDR0AVhSz6UAepdjMLTBX
qk0tU7+/XGSsbU+fpo+Jm0Fc6mh/HF8z6TSjg/ZQvKMWgKWgbj8rjxRvFh58DBOfSuzuFhr/Qo/i
Zptcui863NVGFPtjltaJcxu6/pc6fqBsKbgGAygyLWXNXnFrYsNI/AjFVBH9+wT0bPptj4cSyNXa
6XnunFQoZVudskBQ1pjMW5bTX4TouqLoczjL34Cg6BWoCOCiPlviZI9n/sQePd6kqxjltRQ+MSIz
WeEzAjjERXyFp4I1vOvqVis/mqSfGR+6yyvjq7cpEABcPrhjfcJ2sT+5WLXfT6U6AgFVRBXS5Ifg
qcb7+Wq18dDpX262PBG8K828/I31rxZ/HxCOVIHVcP6Nv0GuHwFLPgqEXNOWRiPbxW/zBSzRW7UY
azOQw9+l4YENmG+ULBjDU1+3dNRmz0r/XKlRjJgIqjil1cfwK1IsdjHYUQxMUFefgSqxHbN7ZApB
G2U/MaBKcUgMxhF16wuhG0SwsaVFSNotWw4ZYtgkIx8aaSCs4+IBoLyj/mMCNhnBDkwqT9PAdWvI
9ZYPkMrqoFUSrDZ9B9zVlVMBspbJCmFe0OXUzFL59oVtJ6FydiBij/WQ5V5zvUvCxIi4DBhN1th4
CNuTfHp/j+PThmIhUw9H+Hggn+DGQh+1wyxzQ9Tbzr3s2DuZBfluFreV8utuyQjKJDoxf9tooeP3
woE+k8YbCXYLcyGKpmsE5WrdXxwNInRNjUIoYSiX3S9/WVTeoe+FH30fecA2IMXTQ+UIxdEAPsRv
87qFeMBnYy3w6+sZ+ZDZI2iIqXqVokPnXP6iZgYS5La12RQU2MW/VbsavUiHvQn0riLXoYxuUMFK
Clz/6e5wuigCyEUrw3OupxNPn+fuQDmZZQyD+ZNFSOnthfWQh+VWsNTCIMvmzh1VlYeT5inTDL5M
F6YrWtIcEkIxRAPjkbfU7QIHOe1d1n9xzM0oWPYlE4jmPMp91EsYi0gV1wLVHFcdUo6rXlrbock7
bsT3nH/tPS+kPb4GugNXasIDdmv1SwK4KyddUpwN76ajFdudvoSvSD5Vvc1DWDZY5PPAPRj9iGag
NUC+roqdeOm5YcynVWjSnBDUQU8A4aCNkx25bRdtSE3q8CpoH3slDinwKT6pxBW7xm+ARQyUQjf6
TC7w4WCf5Mfql9QdNxQlJqLxDXGFbLe8O74S68TP4ZzM08I/J9w6qL6is/3kDcOva5z503OgP+v0
FElvknUyXRDYyw+xYterCs9VucDKFzqz+v2saH/V3gCTQDgZSqa9Fh5supjjQ+1LnzQFjgtF97Jd
t2lE1AqiU9kNOt/n6dM/d1Oz6LF9ftJRy5TV/RsFME2oagKom+sZIO5m+1Ymcn5MDI1BMQq6PHU1
c3iQWzjHX0QHPJT+TmCVDqe9s8xZnvJ0GF7cbBhuJSmxq/tM9NCxpsgakXIcM8VkekE3qnq1rKJ3
PIObhnizyfRkLgX30wAguaZpxKoDyE/1Gsq7f4OguhdRPoCsfPaPM3dowfy+LxfLN7DGO7RrXvbO
36H0velBoXCricEvYuz47UowwaqOpo0yGOTK1Kg29UYrfKPP0FxdXqhdxRqiwGA46MLJ8fJ5kA61
Eh98bBTECfjUdUGfrzORSQNRunELrhlIVwqmN3aDq0bqTsz8KG2+pAiBwFGc0KQRII5Sel7fEjTy
kcdZVsf+oWupc4gt3T0JMzXvhVNDqKNPMjiWhjdPjABs4d8SRPokvcJH+BF8y7NBcLQCjVK+j0sE
23rIeTaEl/OuqzSUH9JdNHIiwQp4XKMI8+LqzboZfOMTNyYLCSPjvcMheN3R2zkh/z4cGQy4cyeG
qSP6iLZOig0zZzpMnHUkqAa/r2vlaB9O9Lgdgv3TL7mpmz81vxr7hcGencOKePORKPTZWd/IZF1f
qImoty4cBsXFbEDdXQVrB+G07LvUJGXcyoZyqtvYsROHZkUVjG6s9amRDz+KRIPL4dAg1Z4gGNPT
qoFUEGABtWnk3uHNf2Knsno5q3qh7iap4JDx4vc36K+gr8OuY6DlyZFUw7dKCe1MlkjhN7Hhi75T
QKyBdz/EH4D5RKRyU0DlzJ1GFOtv1/zHCMceuhiRMbgnS1dJrxc17PEuJd+LVsFqp6zZD3XPDeKi
vEHQ7eBfRQtRLl9068xKMqryGsItGyzlOQmNgfxsdtAJ6ciUnKZHctS7SvSx3cU8lfYqfNKpgltV
dP8aI/rd3ddGfrP2vhXiKDa+GKXNvXYMPnMpPpbwL+v127p4mbiUaWe236epNqz2KSS5VkqsLtmj
3wt23hjUdW68FByL5HPIwICUV1Wao3QULhACOnYVZMx9P6hUKpeVEEL5U2F0Wzeo4oc48MdnkqmI
xogKDLXjF/1YijHIJ3Qp5GtAYgym3SEZIKlV499N1PwN2zUk/RaRzGhBt6vIc0MkGaY42a4RqoXu
zpdP1M95Nu9j6JunBL5nR+C0tZJqxksBEBICVisiQY9Y1FuMbWZD8BTNKUcvIcB+fPU2rs9wzQZT
l0MG6nYiSXk40tnbDI0/glvBs0sxBAY3bcJ4SFkaU++PckUOZdNN+blgOdDeJMWwu6l2gRTBdYv6
XJJWfRZtrA92H83T2rAYvlYLg+tzGduubuiGlrv20s1d5YXUKJFDSOZJuqnXWU2bKhygMjGj/Fz8
z0Z/L7jMJ0ov/Yax35/nwdEbGPa7ob2H2xF5mX9VDVDykZYnvqAXjaWX3jsXFoGvEdvLPqc4lIc5
LUG0wNy3m4wh45yFDO1dC5mPwNhabDWbBFBO0WkIsrKPR9UcwCdj7j3pYKZ2RLUadThJ4GojuTbf
pWQxFiWqC2WopKUp2T9mie1evHMdIwHrkqHjx6GvidSivV8caXPf9lxxPQtYRjbqItoknqfLm/MR
jMYeqJqVOOelYl4ag73vE98riIzcDQNvF9dk9lQJNx3KbCQ2ctgjUh7QCQ2aeT85Dk6azxxqA6cA
DD3jiLWgKabbZgpf3M4s4r2GPChLewx8VwGvgo4fEFjgBqju9rX2aOPkd/2zYoVdj0HBwGbuhF9A
T4syVBRsa2uXvewfL1FnsKZBXkl5tIleGKKlCzdahgCJSen2+Y7HSlMP5AJypDJ1rWTYV8V9WNnX
ZIXjt8VWm+pU7f/6qZj1KHvRKQkpF+zTYPB8LICesJT5xSkTJtyHpM5yvMv7Ert/7qXZ6zAS8Rwd
ndpUWDptrbQPGfyataSBC8GVoRgljzIMXZYj44qgYN4SjoRsG244ozFeEq6hrc5gAS8NnduW4fQw
imwc7jKZ/hxOBBtjEsTTYGq5EO+fU2tD9bOGPUrfTMUpIzNPVuPtw2CP3khU9iseJv8OIfowjRaF
j3HCz3Z0/ihvA5OphGODV5Gs/Tya48cSnTojiF5j+sSxf6NEtVNC3KvN2vMmFlfnurZYt78SU3rw
zHO1xqaQq7QGdCPAQ34APvyHpHWsW4AAXweXKg+39dTGWu0hs9pWmO4fkOL2kOogh/ThQgrplfGh
8daxDXtFg4jUueSaQ6oriQ9v0l+nAHfPSo5N9UhmtJamx4qZbP/wpuiNfe7FwSonNoU6UAk7ONqW
ZCfxdTkKwJVuJRG4RY4HH8Miy35MSvE9Za4fWvXxcZlIiO1f7XFaKdYD3nm3M0qIg9f90fAqU9Mp
F6I7cQDO7vTacltPnRSTXYw6DgnOBkUFUdmSGm0d94FVx3ts/dm4ws4KoNKhyMpy/OKrio1LZLIE
ODeZHqGr5SGzjm9apPXq7DkNKf1zqSmfSOn6nkixxlO+jWH7zZpnN+xd/HHMvyTW1IC2KI1A0TDu
kycQcfIke0NVKB6iJFDjMhKIw9vUay1XaW+Jje7QsOQPPeJ3YcU1LdxiogywNJiOczOaUat02/GV
zT8zTbUOwhccG4b34ggRxSabdt/dqUq0+9o1TN6pKyO0CdMfathhKVShQXtnGyeik+BXKsyZF0Bx
tQMCtGez0Eq6o59nsZUfM7bQLv2D5A+YYnmCpqbVmElNhsLkjsi/YkhN8B38CkYHx+8HR6IarROW
Dl/DzLtvgBK71l1Usgt6lqtA8Iz1+AKp5kHS+qexrEpGUGgrqglpY4Uzi+c5uA76TrrizTokZRhU
x/U/ZzszEJ9wKfqJJbExlWtuhmMnnuW5obXk9MQi0TGWTKSNKaV9bEuTeAumbbizZNFWeDEE5KI+
I1S/9P/VK4WhwnvtS/ETnY+z7LhDNqDkMFu74fXqmm3LDSmDGCazyChRSF6ZAwf+lWwKLEytvVFv
qrpieV6j5EDb8+p5wPycbScArvyL+DbxOB9yXiItl1WlO1G4iycn+pxCqonsOIarzHR/ptxZzRAa
k2sauGF9TPw2JiKsYYsA7g6SsiXFJorm8YI1GZIszSINn+k9TT/C4VHeeqjU1DvROA8LL2wrBSlB
57iehwwhB831cs5pquvEj7lki1M1v5DpOQBR1ThIu8D2azHP5N5iMDfL0+KMvNG4JnIwmrAft0wA
/kps8mVOAmvcoATzGI2CIgOs3fGLvdo5WF/ecgF0SBQ9Vo9fIfbRqEbPNSxKu/txA+epHFDyQmMl
xkJO4vlbGSVqx/0nMkIHYqNYgatouZZ0/Nf3NJnUy1rBnAOWuWrwho7XGHC3VVICsCDVoXKsahYV
BhWP6gNgBqpzsdv+3WUcPngyhfotYVUWz3eDkarERAxtnG/8gCrpWPs8gDPBGE1MeC9/uOLH0QAG
dZz2rGbUMi+afzbMpYvgUYeuYWd1vBnDmBFUBQNckaCpas1GiBxfSV8k0uFgHt2csNlouj8Uf42v
G+ILRZ79oLRXkZmbpB1ui7ROlYHbEPkNnMswq/JkdMbFAteTxu6CsTqGsjk+yxdl19XDT2nYMD4R
O58BmoZeOz8QPqNtVPpOaBtyswd/wjf/E5yyM+rXNaONCnlVoKAljhshaSqwz7tTJ+3rJsN/B6yn
LMCTr8I2MTOhnul7U1VP9QIEW/z2N7og50rNQ/PhHnszql+kf+ryoPffuFFq4m/ruHJ2MdQ3Qs8B
d8422Wkfc2L2kOvmnMRWozMITxejxCOJBgxn2h9FZhnHf+BYbqd23OHzWDxHbLwngoNQAkTiPT2l
43yew0rCMvytJypgZIwgU159LQNfs2+cP8Bu0WdWtD+bMsucHDYDqpqrwjZChJiW/gmzf/wraHYe
kVb5jAO2mFiSzWalf6ZjdZS8Cne32CQZ5TXqKYLmtfXSr0XQJAUJxVwHxbDXVUbpqznO4IxuXkEb
nDIXvMHMbQgEom5FCy7NhSFgRehVxNbc0GADt6s5q6rvgh2URMVjgo2TutqojpcmX4pt/vU5pAjW
DyVUfVzmyWsEo4229c/EXjI8j5m//pe/bEyFr6dBNsXSuyIwZhiGynG6M1vUzdD+j4nQPWoxQ/Se
0ok/6GQEgA28CNS7+ol7WBuqxX7R0gt90kAf/qWSd5BKQPPFdk683z8e3cGRi5e6gZydloKvdKoK
4D1soN78RCU3CcAcZY6duBVcdiS6OaHEkCZN3cJHDFACQESYBXsfxWKTuhfrc6z3iS7LjHjsAkYF
6oQ54n/NNqh38jujWKzrDiCDuV/gI28f8M29rfjca4NZNkj9SbasZo3vlT6jYM/bzpoUpYPW5nSp
cfFAFAtub0qSufs8RCXA5xFQrGEcnN4MKSTQRF7bJaGHXFh/oGt6N5zCdFjz/sPGftXCl1wfS3GX
drvubDGz6djjF4PpqrB0geFFeb8Mv3vs+5AcggCyJ/YyJggiYerdTdaEJlRTLmNuyAGg+CpM9DaO
+h22HOFCnlIDWVVWYtyoVJa6if+Bd8SMRJqjWee+My/PrzJ9/8KDTFrIowCke5nDxsREpQBwGKtC
VcX/yfx0tm/+4Kd48Hv4U0T798f93HunyBMxl2eF9FW6T5pXIWwAkD87uwolbFTX2FWT172jTqqZ
dgM2J74ay02HvDl1T6ziICLhsMXVKzjX5nOr7wUzSVGOO6Hqk4wERIV71L++zZSSYUnF2wALLXe2
FLD4UWw8Ef6AieVwYawC4MRlELmfqxTf6gl0cji60WvgQ19dRwP+lh83Kyji0+2cjPScbyhm7Pzk
0WpB89ameIRqKeMAn/+NX+K5kTzaiMYhoJ0CN3ZgZIV2ojGsF7rKDd1Y2C/86YK6r6TCR/az5kXA
IuMzi2wovQiB9353jNaNUPd9ajCEC+QiryOa86os+0wBTUXhT4k93BwgslJGOvyCRseWlom3SGd5
rnmIU82cNwF4babW+DWhae+HmeWnpn+UtpFrAdeALBj3EVPkzrhjq1H2HffTzSWUnNatnNoBocpB
IK9hsYNPGMJh7AOPVjnoLuIYoxBxUoxiRnJYRvzd9G5gCrp03+AgMoPDbyTqvRV6WbmkUsskvB5u
UqMwYYDvtv1ren3VxNdAl/yfSnmLFstuyXfzur0w8xQBCueqD3MlyjDyY4DYNpet6hcoWh1tonZb
Jx9X9TpzeUZQeptNH+keIZhSxABy5nX/+fXmuywnyqviiXwoEoQpVnO/3iDiimYDj2blqIs+RjTN
X7zDnq5ENxdRY98vDSyAef93dkD/ygi3txkCFYsZmElfNsvkPBnjEr23KqNyVH/C2jfmlfIJBsWI
2u/kIi7x5WOMziHFjI/05BGgvPUgvB3Tt9cAAgLGOV+adK+ppursE5s7VctkcZ6wFElcDeJ3URQi
p9uGQ61S4e6V7nfThn4qIbg66k5AfMoT1eGELzJzNY+JkzwULWH2F/E5qbSivrE/ZJCojDyRe3HU
aoxL5Tgq3brRJ/giPW4w+p7ppeXJyX0FSTI3KerLV1jTDakAo0yDGFHkCGgMoEY7g02sP5DP/jsr
dhbbTPGiTv39iLZTnbw+6wjBTqsYhh2zKwygXSFS/U3mNhRUDq/vJAB9HMFUmGAUHpJHMiVtI1aO
3CYeQ94KLXmhCnM2JnrBqqB0w2IFBHhdvnmEYYmw5izL78Tuv2CqOjSmsV22Uqve/I7WQlMQjpDm
Uo03T/lTFTxmZwze7ukSRl9DVBGn5M9/l/8zVD1MRDZkjFSfeAjWn8GaBIaIkszJc+sIGA1729T9
J92el5KhG9Ik/5PRzvThEmI31UD/V2zuaH9j5uKuA3j4ZBTIEsszw6CoUMM2jQZ5dH7iqa/YoE5q
uZpO7uqE6SQhFFGncmZh6OjdOQFESC/Ze7w9zm2/9vYvM3DRcNyMdDSSaevlcdyceI1/jTWxw48x
3RK11osIsaf/bfepMKWLw9nOajXrPP/ArE8jhKI79dq1tlXhVWyCdJYkfzr7fQTs6zjbSZnP/lT9
9HyxvWVgfksrHOo5U0iiaICLhIV2BknDgr+mK7RSzadUdZEyWdEwDcu/s0ifA7BQjJgMytJLp9pg
uMSzKCDb4Gl13IQmZZ2erNeT2cv8a7n7VUV0L4QYd+oOWaU1+o4jutNCer0SstokKENSgEVu4LNS
08fOMpatLYcMruRruDsAZguHdWy4YzzDouq6b+7x/wRLaxR8DJWcp0Ng1tvjb1hTikxfaUGzxw7J
Dn2FefVQiWlSmUJXqMw+Gp9DjiIWxnHjB1aag1U3lP5GgvgEjhl/Tnjj/MwoG9KJCaqxvaLz7CgG
XjJCw6j4al2/Lip009yZXmwO6aAfSHwolvYuT9yAjRcgdETBUUbhRbZFp0nHIXc8Spm1GNxD7Wo1
iOLV7VuCh16r/LmiZfmqRbVV6jynQcegq5yWqETOYMEE0EgUHbgk+rvSFJGMc8lT3PXXVHYwcvQo
zkBe2zBbHqdfqCDf+54zlEVKjmE8pil7DIZUmCs/sRIbwoGjEBC3FtrCRXeN3udLxhNTGGOnbVoM
2L+5n1zJ6ATLtsMZrKNC9ZAFUwlUlHN9b1dNvJFSUTxwWT5xjXTk8ppQMLpTz33YP5QPQk50T5kZ
JkFpFMnhrhBVyQey0NrSLV3vZ1AimOVsLteQXAlMOEfrd1TKmlW4949mMbcOzapkO+La2qJg6Zu9
rYfwcbrWqxMCUL3PTz/xFmEsvd7GvuHaPBwN592L1MprtSWRQkti9zOjOwXkZuwvMJSDqL+eIRtA
hFoepWMtzUktsB0lwV1wwD35QhMZ/heAMUw60M2dzDqaTK4bdcw4JFiMO5INwHwhsmrNc05CX8Ex
UNhl9nQU5e8qspxD+L1bZNWeNAclOTq6BFbDuw3xqrVmL88Y6SvLBGgg015lL6R4/XWmwvVUs+Yt
MKuJr+TlKA9HA/774JX7vrHAiE73A0JmE9EuC/k9EMGxfegXxDh/EA0DKNY6i/xVu3sZhKD1KANs
nvAxWsxOCgfARGCoMAUolhlSpMNIwAw0Im9m6oYnSSPKvaxkkI3DjC7tr9xk7EHYYh1WV42y+gqA
PP6SlBPNH3CsrBmHnQLsNxOvFFjCPM7o/3vQ1YCYq+W4/uhA08LaU4TD9cLnrlotn3Oqyt4wadv8
TLprJ2AXqXp/N7SOG1JOUXXUGExXJjRSMg+ZvCQXZelZ8XlN8Zwaeq6aB2UBAYloDLuKl9Z7tyL5
XkZqW5O9Z70zJqC9ubleQI5m52QrcgDs57HL2XgBH0KG/2b9XfTwJa4lDTG4rxmYLhmyS+cU8UIp
fdYgsw+pPTWjw8m+0P+y8f77fZcAIf7CHA2Dh8OVvS2OskZDAVkPrRIIiowjhCcSzM60mCWHHn1K
JYKW4INrTM5r800RBiss5tQHNMbnwBNPZhpNo62BCik4wT0aI9VCVHN4D8jWgrl656mXjPM/n1ZX
VTuzztT8XGyLzxFdwLcdS/Y+ZkOEu5SpWXJFX7afVnF24yo6x5p96mbMrLsPe2esHCjaoUpXr4Ua
p9oG7S4RMldY9vXM5k4hQ+D8PKkRUkEdtZ77tarckmSs0DgUpFw8gzrhjinPFCMyDDTHLIMD1zt8
qKdCRc3h3d/EsWi13B87neKbPNO6nPHrZzSVYmQCJmEaPMPjQ/+ACNmz722vvjwFjKLhIs3mt5nk
V3D3okj5QZTDz/wmq0EVfbrLUu+osMnxjoh4YPjc7C+lEgTrfQN5lKCoXf4pgzPvqVO99WtTtfgr
tZ7r537npwXcS31pnPYFJmk+Kq/l11jPBFc8/t4z0dTDSkPtymorZ9PPGWD5X4Do+N6h29dIjMB8
wdsNPSjvdCua0OKP+WgAw5ZwUe9kW9GaYYBqliku7Z3bPp3bjI/pvTSo3vUeYTFuYk+Da5m0uhEi
42vTymSNeX8AJRvQXBQmT0e83eRAog86mqspd5pX29V7g+kQcqLP5mRDa4viBCJoTsqFlspx58JY
AKSubl8qV6yRVfQ63YgAHeJZ7Cyv+qQp6pl7PYMcPuYQRFGiwfLi92EBkN1xaNntREMIP9F+6Zya
JTxF9qG6LloLa7YfLLKcKMaVWvrqLlCJ4KouzS36HaUK4eU0Kago4A0LygVlQV5tkgb3MsK0y5sx
wOmmtBSDB/f77OqgCI7pPZOuaqy6KZTU74uuVQLdsikq4B2aw0Wbq6UF6j7BgyaGoiAmV5ZCv9gd
wHmWaMXcTZzFgV7whGHDzn3mqmBcJuIfjz6GDyAryW6GftEvgn/pmaBBEuKQJhJJU43ZzDxiJEBq
NipP67AjjbObutB5AdFJjlbEOE3XChWgdg4Ay319zrAxF7lSK1QFRRvhCLok8K0ovvqcdLhwT0Ba
i19QHqEcRq6JoQaG7X+nIUox+xmble2S4tYho7AifP8xYA7/pDK9HrciOJ8xTXKkQMrtD+x0hv6z
Zs5y6Rn+wmPwrz4dLiRE1LrUmbkc5GYj8rzXQM20zzaJR5wurLxfEZC+FehVAUiDR6LrjKem1+/c
BVzBJ0lRgcrQNiLSDmze1u2LPM1GAfDXUJ4MdNzv7ewfD1nICzrERDcv4l1+YZ9ZLuB3vcaMk+BJ
LP4WO/a/tGojks3rx22kBxK/A1rf/j2vUWi7ThZzMDZGrMHmL9Yq66EyHTMxWVjs+9d5YmD8P1t+
PyRwq8aPPeKyl80mlwucu8V1bUVKrPA0esMzcF6IlYOMJUp9zpWRTRxTgh3BVjYyp2zMaT2eByjA
AVViNT8MFl2zKuArWGTQo40AntNii8dXGnBO+y47mcWv/uL4eBB8P/aRXF6l5xtm2SphGKHXPMXz
dZt+bO95WN1PX8JgrYTfq+z5o9L5kTvcYy4PUugYCdfrcKJOs5xSqTwhSUh7hOGFkHC364/evt66
KPei4K28J/t+HE/02vDehQgBNmwXNYDNV03nJBLlJhaQNyiIMxyLa169ul0zFUc8+/Cj4Rj3ow1v
wvftT8uiWpnD4jIX6F0S+jvoOlGFWdIcGhGlUjFG182gPrgpNF1VbpLBEL24hSGP6vAwildmhEfO
66wrOgAyczqt1Xh9HMflEuBBdcxcPyFkRkOTw/1nVHbSp+VmPCycUDv1FeZQiVWDs7EI9ArnGUoG
d53s7M8VOUc5mCtznFM7fBTc+yAj16f2opT2yJxPncxWd5N03KMl7GxvJhuUhFNSUwKc2lfmKQgv
hE8mB1lY2b7BxYWhKnIX2NbxkM5TN/fLV1Mc1ukhnRlH3Vg2YAFPY0PpiWLVgecZP3u/RlnsioKi
VAlj6eb0yQB2iDv4jhkHxN9JGFcB59ngv+c3nOHwILZfapOGaEaJlKvugvWzmJVbUF2HCOhSuW6u
VV0QWMYYAPwNdGovrA+Sr4jFH6KDVRZn5BevM+fC6XwUIuAwLrz4VBBCseYvwObK1LcYjuA7axu0
2bgfr0m65W7azQbHL2TT4LUHc/KacaDDICSHQInDezhyAuVUr6RV4vrASDfxyFViHaN4aN3K8Nsg
M36CEYBf7NiWtcx+ETlh2QJupLlBSUsGO5UOASz68mSoMpaXK7Kbv3pZbj12X9r7f3+2HsiHNrwV
PbhIi47+/al9KU7+yagy3tM/DT2cTfxYQKb0648d49mAcmIVRp++V5hI54wVZXgfAE+T7v8EbLcP
N/VTjacCTj44wKhze/bQZMdKPTK+uf57CcLJLRhbbM1r/8Y+jlXqwt97wUzsbXC2ivfentEUAXL/
RetYGJ9saS31Kv+Wb1DZOkIL31i3ONp+Nt7ZrBGOm42KwFaGlo3uY+s1kmDFsuMQPltzhMa9iVps
Z+hKO+ZdsOeuHVjCnh7MRoO3yW/f8odVS6X0+mdol0fBU6IznN0V/xNwUULH39TFOhGXFFfpos9s
HwkQi2C6+W1L1vj7HLciZsJwK/095OYz5oJ82+oZh/zLrXwAsMiooOTrBPycH4TEgqjINU0LTh9s
ZfE1qRu5GZj1RlJ9GxCmijqZF59jxlsc9HhD/xCm6D3sRpKNR9JUg/1tSbatiIgAAepQFyxMyf0H
UFB4ZSLa5WpynKy4So9PLKh9xP3wEfrzlDMoIhNhMPqqPtSpbDGzawBw4gk/MvNoqBCrttWwmKSe
taenftouSCSfC6RsPLHDtdgsmCuUT0lIQHjFAZog8hv6snKg08/T9AlR8k9du/HHigvONAUxk6Zm
AazvKxlphAyFoHsvhVDYvNLbkCkdMg4Izg7aWG1/2vEE9eaJkE53V8tX4U2DFvamZppQpjkGmST4
G4wL+93qH9TTdjB7IKozLolNEMJVAKbj51EC259WUbzGf1MMdJMm5v3mnKjLyFibt1vN/is+KC7H
67CutZBnDJTQF5Hlfd7fs3KYFZjnOBGIO+HdxYtUEc+CxrcsBwFQ499kf6RWpaSl9y+94PDt0DE1
NeyEMUIiRsVfhmADoRc+LrMrwnmQRfkL+1DPqFOyxoqz/QqILmBAiuKYyuhPrE/aR6VExSBjX3Jj
4yHtU4kbWNEyR3nupebubfNi0ls3Y1MwggfTepSZE5+pFqfQYMZUMB63oNqXZFiq2wDQ9V6Uk1gS
/DW0rzTGp1ZaqhHF47dR171mV/DgzT5G2Kh0OFP3lQDgtTkFtE9mSf76OMysrohOWGuWkIAl9nfK
r8SjP+brNt1mCvOKjpOqbsQCMQFbnnsA/WhQi8oCNEyvLVCx3qRHHbN4TxcH00D2YDjitTfbPgdj
yvS9r2VqFut/0yIw8wyFRDlriGljtIbbAShhFo5qss7fe+AQqQtELu0Y1damlfPKqxh67p92tM9j
389xC+KKeXmvQiakwlkvBocliaDiwfk8WE75BefGe7PvdybmLsO4WWDAFPFLaMGJp8phjcv5w5y0
LgCPcySvUd0bZuSfvGwuAy7TSvwKXMr17x+y/wU4bx7Grl/GqxJPk8vqvHw3ebptsT/L0fP+o4DF
7oQVWD1LYplgViWW9aI5y+NZ+pL78vg7d7qejOWHYCv1EaQY7TvL0ggeHwUr4tt4FlFHeLbRVpuD
WFT4PcL85gAqSlvBUgaEFF1o1hceLjSkym+zW9qMDGcZtWiz+jqyySWvBagHYlYxf3bp5b6uBx6c
w8yT2rM/qcYNRlpzL8q9gvh+AuGFOtJZPbgoJSvOGlc62hGt9Fhq2WHWF0YHYuNWihzF9SEsgEtO
MIIKJA4IaAijblx5pzBY/ofa/N9CLZEnBXX2a7T8S+XsYiwwZ4W9AsdYBvwhvqOWDNHyj0gUUxVF
Gi2UEfEThMf4n0pQsd+tGRBuU2R/pp9IFPqfc3G8RWWaRTauvc4Cu4YzkPnOZA+tgBG4qECQOq5L
bJ7WxdpB8+8/XzFoRNkSN9YbCnqIx0H8wLA1okQ1BeKKAnq7eydW5S4M6uhEQj7tocj/PEwrm/6d
EpjE7JqqwsKwMIX4r5aLgdlnHAzKIsli+ipcJg8L3/hPSw2nLNrd+I2QZFPGi5fm8Y+uQCXqnq6y
v9c35LrjdokM8ALQ+ha+0m9B2Hph8x8I6jlk9XylrIG4Jw61VDqzSM81sh1nBbj3JvEW8QEU3tlc
7bM13pDM3EZs4V44QwNGfgUB1Rdanr2MhbQ/Cv+vlQeFlAceF9ubjGxcPzjH6LS2lXICvS9nFFLZ
UYw6+3O9z+ZvYx9HrUsMDtNMx+HR7qd7Jmn+1jp7+qcNz99Pi14ALc+nWabOKBZb6wKci4Hdf8kW
XLk6kZe9aHek+bpjwMTjeRnPGW/ERQBooGOIecuD9hT5c3kPghu1MfxK+QfsX8UYbXhUjb7VpQhO
JjFI8T+HjsBb317KrVDAx74grDr7xG2PIMbHgX77roVt8EDoM3hpxqJr7nhnpFWDoLBwSjhcQNVf
hV9x3KemrP8LyJhmvn+FWtwI6XKGy/TRcug0Jn4UcRIafNuhyughmsPa01t5VgIljmCSZPHl/Baj
8afmVKPHw7f2NwIGzSaREsXoIaFfFglodOYhaqQCtQPsOiwzD4Scm0YG5YJ0CdJgFdEjKEgKZ+gN
bjBD0bXKELRaz3+6kQ/aZsRQzmdsHRjDGX4c5tUAakCZcU0iYFbeDkVPm1QeW/uVda8RUIN6EMfh
xpCgJG342ztcG5i+cEX9l1lFUhfDWE2qlxsP4Ink++xk3FaI73iTdEmAdP5Or5auTnZ7dAWttr+U
6Q+oQ5zWr31nmPsnV7BZAw6TUOmFRYeUHMc5OQOhrrFvy0RXq7MYUM0DA5p7Hqsphq5YaeCflp1a
0RztNYTJ9itq5QLal0YJqFrd/csMaR+FZTiaKUWCHTjW682pzH3NGf4nH5ebjlgamvEel4JnQbI/
Ksq0VFnuD1mqvinNQXRXOz4XGTkIRhzIm4IqrQi0fvgZXIiG7Oh6cbTxZVyU7Cm8A6LY8FNrzlaw
g249TJf98tEUkIL+VInmwO5ARrKp5iRLMhvRsGMGV3Isu8PFXJNPdqHff4HoA/GUd9d+V0Wkd6CM
DLITuDbnkxHQJBlxwA26XGSH0KzYo332YheKBZWOwm69cMImLtFOxVIAZct7xWAU2CpZmA+G5BbZ
Qv6FmmglXdhivDz8yYq6Sd5ZLAytnk9uVNHKxMpPhHSp+57/Gtb8CKQRAFrVXIAaD3ngOEkeQ3g/
QEG4wmxz50MtWeNicY5K29NXdF7SQUBeRm0AOikEyPXlEzHV5/WltP146J8XZFHxq5pJ4C5EQJO/
WAFGufDIkmT4R47mrkkRIZmSJqfx2PHblCMS648D1Qhb3HkYOak1xEAKB5Etvgza8SCnbyDlfHqm
HXJUxr/QcJFenWLRLqL/LzR0aIQ2KdmgZ7AsrnfjoXkuB4bUL3iPaYoQrxs6n+2Y7WhEu8fbAqTP
YeU/Id/WNDzo1TBPjNYmP+cTFtUKO81zDh93eKy5Y1um/r2365+RipdWdtiZFexkBp96UmlCEX7o
8+YhNMsQZvk1b812u6+RfkYx2JTsGzMM3cxVD0PfamObWSL+2PY7QqaaXOq4G0Up6U000TikhfRF
FN0lteb72JDmXyGywpLu1uaiCyILOfZhNUuAtbvi2xvENtfsgH111huRV8QvrwLqgZ/t4tnhqvr9
Imc6W18hodjCq4km1YpHLpTQKUseAwYDnLznCoU+V78Ckinx/KRK2hXwqYwUR1e26Xs7vcC1PrDV
NZf1Y6NHS4tS1PxJPbTfOO6N6WopJlcdhB3omZIlF7lrpMJZ1tCQK+LYAay/yhncO1xBEKP7C9Gz
VZkPyfFHWOpuvxMGo/gyQ5O5Le2jRnQCKcjTXqj0IG1DjxyeVV5u+buUuE8cSGJ3zFcAz6bGtyNE
5W7tdvA5+jnSt6wO0/58ZDdMrj+veavdGNJ5ZTnoud4fuoXxoLsN6kkqRMxHspYscUJsj3i+f1dc
mbFnuLA2FoRkMjO5hiVc74eCLgny0iISrEKqUx4xmutMRPdCHzBOvj6av9eCFIP7NdWHNK69S6N0
6nJ1gDUqtuLWIeUTqhNNKU4nN/x7teew01kKIvfZxuskvJwFQuLGGPo7NTGJT2U8vg3+Ef1/FLS6
PZLAPbtle59w0P98vUnpggE0aO2ZIu9bc4XJvrm6GeE8WlJPn/I+RVg6/8iDUPIaulNl/OFTGZmI
gstoBCC7VQEZFuflp+6QsY6MRUIeck7vH1RZM7jr1vnIa8X4R/amkP+z6TcPXIA6IzTq/1SssyjU
Omox0OrU9NDEpl9INKkBSDDkfNdbXnyFzJ5zbVWZDwPykxZRCJbEpHQUGDRco/J3O+cY1njVWFBM
xo+B79f9Qd28Hj4CbHmFvEVWNVyo8Fh0FyuC8o7jveBoLjPWSGnZSKRJN04FW8LFs1iHLRM/Bsiw
ergfni5NSvljFTKdSnGtDVxbAQ02Htq0Dwkr3VZtfktuYG/YErgWCkNkq7oQJNLIlF+/g9c7f4fH
IJQ1AJTVG1ZBl4RfARBpSq8/4nPiCYbCLxmblnLksKfHh9BpTe4f/q/kexmArBJ7AVMEbHJmG3Kr
XXY9IYeeJlLWPwZ1d3JJijZPwNlsWc5PF6LxpuzPtcFVUqRlqRPJSNUUCcM7S/R4LhoRU/Zv3j+a
YaDmJx7Dn/Tyvc0UwFww9r9ziieKDRRpBpCWymkhvgKM5kHomlBwf/A1FwhMR6cmaBtlXH0mQCFi
dzrN4GlbMZMpXfUHO0LFz3DPfxULqliAvC0yV6gixeL/BvZf6IEuEWY2veX5+y0cMnRTXS0gotgl
K6F6deROMTU22iQa2vBA3kXKSke1RcWdSgCKqjLFpwx9RaCIOk/HXvRI6z6R5odvDep1u+TO9e1N
SatkNFAuIaHT3DjA1VVq4TG00TKpeAhShcXicaY/hGG87awTaUbSCUH7cCXEC6P8nvKKX5jxzX/2
N62fwAz1Yzw/k2tWWFv2O/fWSKvemasHvmO+cQfyPqcGlu9RsyrtoXbfGKSSGOW//wQL3bWs6/B4
PRMarcETrDZnwjvkD/MgXwEvt5PqbUTsfKbXkbb8qiRqJIROIDj2X3lQ3sek68RJHL8PO5+Qn8D7
Es7A2BGqX8nZfj74NTnReZnR3BD20iYhK3c214uFUe3ndicb2D4lndP8Vuj2g69ZJQCVmoZFoTf4
HqYyA6QPirtaUUt6NGUTDzwpD5oFdoYRvG+bAvfepJN+8Z3gTNS+849UC5osy4crHbCv00PiJfBK
4r+DpPlW5lndSLY9vbSzf2UaDbOdOTLuexfJH/TqGYpO+WImVQs9WoVEuHlSZDSSCbjl0OIhZGIz
S5C8J6DGcqQYt738FIUukVikpcfQgqnuKY8sOxTxfsngkqGTWR4TyQYovFUPOmA6iYQlhBb43GAe
IUEqRudbwOhNI9Q/FsENt6wBhl4nkCSd8nKqmM1TUsVEB1RGU2WzAP5PCkek+mcj5ILeHJ1Daj0Q
Eq6fkphxG+g4JHX2E7y6QOkXAJaKOy/kJMkrQ5xO0VZfZw58qkVnxIk1eV3QTuUF1LIadS7AO0cb
Soi4xCTbOsWMqrpHJFTwxe01w8a5NAXxzpw54gq+yUYiofzxpU/U2ZU9xYpnMVCkjZozuBQypjhs
XSD9kYr2/wo03tWNB5niQSnPTMhwtZbyuaNunQ44O8RXK5925GrQYunB2KNMMJNMIFI/YJkHHxjR
eHBqAwiB2ffqGRQiBJgrIv6UcaWsLFQk7jtDYoqlYzNMm13voj8VnokWPYT+XpYbwUpXYkstYc0F
Ipt9bMFF4mbcysVzipJ2EefGHuddrlRD7t6a3XYbNweAb8QyKOdJnCz6K6CMlXrGD/s6ExfsM962
WTOT1E342c87BYG+bENOnCxDdR+JByxvOXkubA9OytH/4QhVpryGOYTzVFOgKO8dI3A+lhvSbzZa
6bD0bTfA9ZIklzyDURIsLuFhrj4LIGTYEFYGxB5+e9+NGCsekVpakzCs9tphNHbEpXvPfp6LWOpg
Q9aBESFmINgyGUJevALdKtLoZUKRjE1mG50+U3k+L/HV61v9VN3JtvimqE8Z2A1vJg1P6IKXoGCc
E5t5DsXPX8jpvaUV8v11eh+bq6xLxMxaRAU0klawqbRHRB+tXVh2jQ7VOM9zCoc4D01neXUkOU+/
HkzQ9fQI+AEVRk+vbQ9mv8wUwj6wQbDATfW6ir7R7CrL9P9TjRFn8hG9R0ExogmGsANWpUqmCHq4
712WU+hza25q4iFs1vW+D/UggvVD7kCmeL8NtFoL09UCVQBYz9u3oGT1hZ+2rh9K7R2dqIIYh1KB
EUftYSShQMxDnWzkIrFP+BiO5iw5PYwixa06fiFoQk/88eu7TFtV9CyqFM2zc1zi9TOMoQ0OubJs
kFyNuaE7hlwxtiCySMVh1wgpwEQmNRASe9BYr9O4s7SLxOVq0Vq9btxQ6gEhWYMFO+XD9pFN4aqU
X5lFo7tU7W+RxBse+Mk6kbwLkQgNNw1kyMbKj5VBKZqOHVHxS+QFhWw6CI1CVGrGVxgyqUVOWa46
E0EsIkoA7txeYeqTlIDlqcPbXO5Mts7Rfh0GvpNpBTjN6V3JHDHOTMJJu6Y8nh7/RxOxScqLljC1
uFs8znGowsSVzwbvgCmD93SICEtn/ygoyzCV08Tsm6N8X7r0C+d+GrPMutSbn4CdJwArMnhZhkfW
9WwEjVqwRc81cVAlFywZ04MSFb0m6PCnhkfeFUGXgXDxMZdoq4Ww2ltJhU4puLvOKnxx4kzuhb2u
ejWiP0niy2C0LDdxKKAX8tc/kACSmIl5JG9wCjMEgizdqrTmnuep94rJZUuWlkRl9yt1KX7pA/BY
8V/4FjHWfHc7LrGRzPQ0Q/7nqrpeewCeMYEdapZJvAVqZULpjVa4ikCG3inuln8eelugJm3ywUjU
FQm3lVN5aXS3kU5ipN4P/UkgrB8bawPSEG878IAxtiehmNLDMs0T+TF8zoHndRLd31/H1kkDz6ci
Bn7Fpmp+wfWSUiUEor8Xv/l1+pswo+0HCtDRinRKr9+46ny/YlNKHbX8XDGg1oYll41PyrFnAdM8
flU9/7K6CLACuafb+SOVVvm7bzpTd7isGFQCghgBdnYRWmMt76wTTDn/Z8MRBVcCuCw97kfA2dDA
gKvkBSYyNE1egYnt5VqmYwcQ86Q0PHwL+Ph0GPMqwCArkGc5UfeSCeCZlv63BTCA247ITy/Hbabm
OPrhgNL72Ddj+it2ra4SsY6shrdkssUhGWKKX1K6KeSLxAb/eZjmhVQ45egPlBIL61iWvo1X+ctW
160nCF4Accrwm84SyGzRTaLt9npzeflspoz6Iw+Dl4y9mSpj+NOHlMWbL9ku4dPf07A6pyUHEztT
D17P8PVEYGD3yWe9YRpJ19O0PmVGNWjsZx+fJ32DRSPNq8XfjKZnFVwY/Ec9AN5joImO+3Y/RVuX
9pB541Ijd7qTVBTQNo3SPN0HmKMiNuh+v20NiEAjSebLlnISkid5pqA9t+QrJ8BTRKVieEasm/7K
ihZp1GbkO4pbeSANdxq8obYKDcNozoQ3IKsZzw3SCUf/yH7CnGrMx1f0pZrF+Bg1MhtxAoG9uAfY
jJj0zVqs2HFa4XuTmFhpeSmFHjgN6bJ1fNAdQA+UeHlY6RHZp/B8XcFVw7XSwkig9yLF1fx05Kco
oD1qjtO5PQSgEWUvL8zpjmf5KSlFhBMtMawzJBoXtsW8WbPOTuXR/qwCKm9F4g0pmL3ubkSJM8Wh
uxTb7KhbpZcl3zIcBhFq20YITWPwvm0c/a4BX+w0l5yn0qs86KNhbs4kD+f4wCWtNImT1qMLpiUI
fSkA7zU4HNuIXDDMcz1o8NozF6f+N6I8kk6babOnw77oJvVpBNeZp2ocab7GCM9QPFq0X4eFxrE8
UpBWtKRU/jOP42Cek9k+D5Q5H+q/IPRWiR/AWQdHVj8oLRMLzjh9RoTxgMdG8hDQxojKLy2L9Uj9
VWrxVWuwxWYozR89YvVIEzLN2K5jomCgNYuXj2peBo+w4cAPh+q0KtUKjWoYywyFDPCuZbTTEATv
Qh/YcKjd3ie82k86OZhcIlvVr7QMw2AzlONxe/Ch3vAmXiTKixm3FHCaAuUBYxKjyynTpKQeCZ0t
2jGEDp9GWV7h/B48bFlsUBVHWzHKsC7n9YvKTfn9tfE2oAHC8LKRvyca/0QyXx45jSbc9qw3Bauo
2HDB33f1Zts84aaOnJQgn4VIJiOW3ruUCz+uHh9g4jUKMWxRKFNifiD0Xuk9GmLOQD5shkqvr2/E
kBOqLjRHnnLnNNCBR55vmvCdCEqUdw1NA3KmatKmzvMB1NjvnRdflOTsBLz5cQuYOcpkB9uc+9zm
6Iz1Ew2qpURd0RA2ty45DV9g7EEpqgtJDDBH5FW/j2kct0A1dZXRF9evoJ7TN+xPTOscO2LcOKmc
CIP5fhlBZJKq0VM9Oj/OdVY3qf0aBj3dS1Ye40j0ojC/MscEMVPWxFvETriqIZficmR3DBCKBRIs
lgqgp+zrczs/cDSJvbHqCViSIOH4zb0XXNxrEaSx02UkDWva0azox40aVo5sqToIXZtH7I+QFgAs
ZQDn98msRqsKWW3j2RWOnRi/2s5O4ICjW4HrLOsWvshAubSImvs3B3p91h8bt7g/IlZlDyBj1rYT
APzOP0iOr09tiu+/HpSlnaRFMyuymwhrFkANjmOj57HrbnZRAQr2XFGagH6XzSUtrU+Lh6YkPVWG
lvPa0Cz4TN0Qqmr4ZnJ8XZCsFuY7e+ycxjKIgQhsk0UUZR70Y3rslCNXspiCwK/nFvxxXTyRhCMG
9gFr+IHamquFnYt3oIAvv2hXLDMCIq3HUpQYmL2N5Mka4O3RP2R4YzOVXVgChUy0pVPkfYDPxQk0
v4c1RDAtQ1tWAihkC0wwnkcFPafUCvv3yVwL/biA9NsDbJeDjGt9FFWzkylHa4cJNEi6ggoHIBzY
aESOAXmrjPkEyGfgaF+4IvBzz9/ohhKwXVn5S2TEY5cPJZowHyLBuaMYhxvbodGxtvY+BrEnCuoZ
inzZ6QuHMePs57OPCYvAHQ9YXgZezj9fvhjNJiMpxJdUderj+ChWzqVtk8CXmBfExbfToQ/4Ycb9
fxvzK2GlybC9BKl76USW+WCwfTSqR1btyPDy2HSpo+A4U87Gjl3q8H1qZ9jdRq07HHbhVlqQdM4L
WQ8Y8a+IyHasbwGjaVdhcDgcFBNzSEwNE2pL2GC65CmVnbg90eK2m2p5kE+VIHsK22EDvmMtKzDm
ITP340WJJchIaKY8IPRsG3MMHllWyWPgVWZLdjH2xjz743uEA4in0c4p0G6EYCv2bfgV1lEoJnEv
moBElQco8eQ7rb9LA4Ys3zC5mPn6FdDSxuxBpmajX93VcKHShj8AVuVLo0f3Tuz6qouZSVr8Bfls
zudWEYE5FeDSmPNKTFASxIynPchor964l1z0Hok4eC5f9Y87xb5oGZeYLLmaLLYzUsPADpw97EYr
w1JioBFM5twNx6iMF2z32kSCS5oVsAamW0u9xtpMlZ3FFtpCDi8p8duYmjx9G6jUUP/tTBF86OVD
DQW/jMPiGy46NCRbmY2NUfSjVpdTxng3xa7gzYWEsBUYrr9MeUPUkz/8hmNAxvd1NqeFYJn7br3N
DQKxIDofDIaO5sdHG6tTqCYq4rvPTfxQOvEC59QkbfqK7tz0Njau5AFxOvNRlvGA8XE7gP5+hEh7
Ngfceq+3w/FmaQhJCXtY4/nh0PHXk/QIez0Rt517OWeWhWR2UZRtcV7ZCtOIMj1YERopN3jYr0ay
OgKjXLam580Kz5STV+WzKfJP28AOEqjneQpcTjZZJmoYFi8cLshshFZTmZ0mAvd09M8tO0arISl3
vQXAoCpWkx339RE5q2z8VtrwoQqjLIgEELsw91yQMi699nPIMhBlqrTCJItp7JpC2mNIxPHsuepM
Ksh8SvlDktE8/19YctgdoK/qP2G27L4rMQ/ep99qCm62zE6KbD0fGCcIKEgb4cGiu8NpxskbtBdG
CIdlxWKvxj/za2QqF830ZN4UyxS7FrWOshCfUt8m/9Csqwgh99S/qJsIaCCxRiZWAF3Dmhpttn0Y
m1MGDWsgkUP3+RoTQn9P6r2um1aJgWdcJb0F+fDJ0INHC9UcMFGyReqG4vBkJyl5qxfHhAqDtub/
nz8ZmhEF31gdnCttBeZVWPswlR9UtUn09dRTGGTk+aBvrvqdhxwya4dK4ecgVDDtbPhcFX1mC1eJ
hitY6NyjnyWW13ibUIaJyEb8JquxEwY0lfwok/bWzkfLZVJ7xGNaH0QtdadBQub6ZL3bl7jUJ3Pa
qJZJ2dT7iu6SBMuuGCTpBd5HiPrS3kMR8xPYIfa+9wl6HrZcHBUC2vpPExYH+tf8bxSLaNyAdHzU
dZZfjSWL60Qfn5J7ubMnDdBol88AwdVcrZjoWl1x9oDTQXU70oX+1a/rpAUhQrb2V4BTs6cwd0SJ
wn9ny+Kj08HxKCtETWXn1H8EO4hgh+7OntYqOQDLRITJvrKwQFZnEjAk4JOX7+Z6nTHoP/qcE8O3
b3b71cIbP+JzMPI5953jlQMUTlF4dLnrK6JgXVddLuDnfgBW4IuXITzYCukEQ2y5Q5HS6fIlQ8vb
Ze3Fbe5X7jxV3TYC8428IKIXHShmpYGU62Ee0ta1FLqnB8w3SzqNpGpy3lOLjafrEpMcDDeGBGUO
oab0g88WYJip4QPq78Hz7paMT9V5nJZittL9hoOqgPuQ6L2JFxa2CyNWWMKz/5YbILPBzQvUoRLH
Oegne6l+efQsl+3nXqsYUZMBwgHFDyklnzoxE9dowc6VBC3NH/9Rk1XiWdu5LS1WO6/f4zk0s3iN
fyuE7EvGtc6aQfTymwjIyE3nuxM42m/60Poyi8g4YRwCivyY9T1wYeKZRbtuDWW7/0cIWB+BMOFX
kFyu5c6SWA22NIvhkQfkeHEI5Doj/ZGwlQZNGITjLL5W+4fcdMsvmijt94LK8zQU7Nl4M4hGMmfk
AmnA7R8KBKZXGqLtCiFjaFgvumZrTyca1yG1KlQ3jsBm6LZomOuKwbbJweMofJJGW97guZ/eVIf4
eQOEut6BnOaHPWZIf1XxgtZOvrd1Pcl8gqnH+M8OjD4VAh4UQ49uygjAVOgFpoXKNQRCB7BG8icp
SGrFMN3kU+pIW54cN+V4YvfoDPWi6NVa7oeF4nwLCK9DdDyk1gSM5r+5qyDIs17Autd8YbCjJMNi
xF4J0+VrzVOnzhev9GST36TSLvNLTaBqrDIQRfw0dkS7Njh/pd1dNsslYjEmjOtWDHWwqu4aMuR5
RUPwjnvrzvHotnvIfLiFHlpzw52dAIwD9AMIlD+/NvyBgjSoSNxS/VGyO1rIINEjD/uTFGcSzNYu
+kJVf1mfuBk0VwtD5xt6Mfnb2u2VZDLPSZTovU9ddl0iyOYATPw57A3Im+m5AiiyHCffmvzQ7gVD
XJNvfo7sGGCEwggo5wWwZZwmMLE6r7ibsPWVFPzZ/MGeYAnYNng31UAHBvma82T76yHELjJdxNCP
rxieuPYlVgSWZIaixF9IORBlF4O8599F2XCqF8ACZu8jwcTsg2tPuCw1zTgyUv9hBlewXE+M+8t7
khURzZ7WsD3aZnzXm7iIa/qgHqcTN6TgrI/6YVnQqpQI6Zr148K2yAVPnlpZu+PkWZiYpWphkeBZ
hIJzb55w1xBkGT+Z+JAinjL8iO47tB/AvBKtM7r9dm7dX2KL6bLG16puOQYs4z4kZaReW9QK3MDn
tapf00/IFDvG5n4+Rs/dvdY3+AaPQ4pbIgzhm1wZ4nfqSulN++7UrDHeXk3xeD0DHGI9SIOkteKs
eQ2iYgK1TLZZ9XKgtB1wDwJk67wx3Mokl2gSyUt/MKKa/AwezZAZO+vc9aGfutQyx103N/VDlGCe
CTul+IfwxxhnylurnvHRMVXd7mpmx58y/O/kyEMnnMrVoxlpZ7sIVRUtvolHWLEfU2tqCJETFTfi
0T773yf0bdDSVewLGEjZ5UCoYENMelmngoMY/NOGKJwGh9lH6eXAFt3wzKeOtBs1y8KSoj0TYoPg
gQJbY4mUepk4Q0bDutbrZaotQ4KtvmZpLIe1hOczWaP4Ft/CFnBZUcjIIq1FeFXRKPFCRFmpm/q5
8c/wH8j1cdum8qUTz55fy08dJZISnd2NLP5Gb/4AARPUBcNlIiKO9GCtjq7ANWs5DF3MMH1w7zuQ
obisXu2+ggujfLnvmVqp5Vj2NLnYNzke0kAyJAvyM98Xc7m8ulN4WRh3OYzQsSIM6AwJZuUBQQ1Q
mjMH5l+U9DcSLYo7PSBMbZfnJG0xJ5uVuQpF+mNy2yoXYYEVofLshcAaFzUKSX63K+7mx7JnM+4X
hd38oE359rWTgVLDn2S2TxTS39o4nPZ3eCJw7xMcQFJ5QyiMTRiEC/fgzrWwUjvgrrsFRyFEXP95
rfHD1TD4v5JiFfj/z19ZhJ4ClpfVCeCNIcTC686WU7/MfoA4YB9hmVumV2imfO2rweyw6z2TQP3Y
NUizvlHYlmFgqpuv4jn8jXI4zau7dtmHs+z4U0xepukFWB28ox2BO+CrkJOKNnyFMpvFIwfUhJvX
TxotZA6SLDVLl64tHYt+0Cgs/6s8+d92zF+JSrVCPKAQZSYCnI/dguK31llPclSisLKVCWUDKhGF
T5PLtfRN37UKUmbNdYZdyPhjBscRZ662Y8RVDNy/Jto9fyWIuEMUA4JUXiy30sJQkIKAjK2sPNmu
MaPuHxnYi8C5XbnGpES9MUPODHGpYf3YmmwaBq0JhjDps60DcbMC5io6HTjm7hZL8wxnVJp3GoVv
L/xjftAsqs91FZfsb50byhsKqVwUZEOcUeo8BSNJZ9jUEyq+xH8FMN1rDb6ULUXn7OAfSx9/oYPY
FH7pQ4IdAafBHHRW3uRNQb8OdMZmqLhMcOBtX/cKTMDifd+4cPVfKODVxZ0AajxMTaV98jdgg5Ge
jE7TRSz6Nathli+G30e4y/w2d46ILJPQ9spvRGxky/CNiGGiZHGcUv+OcM0LwLqcvJwXPeGIVyTd
wseVQhtIqwzD2M9tdhN9oocUMo/plzbhordWfMRaYzG9ODtrqUo1j/FysVWfQ449wdq4bW6nom+7
OWulGVwIwG1EZyLfNFprW02eFRt38DSxfDO0TNrjD38kZQdw/Hpm99PtPiqSkuVlJQeiMDVgtdoD
Av+yEq9kDK4TAtEPfRcTE5oOp9XFzo8BYVS/XxAhK/463oFZvYAUT0YLwRUuPtbwZCvUPwSWNxuX
j6qMq+UkOI1p8IPorbPYCOWr8SSxI8Vox+GVSgnRSTNJGANn7BL91e2f9EfQKm5E8ow0eOIJZ4p5
DxX423lpr0u3au1PAhOXyObszJTV5jA3MJdUcKWqQbwWNRrdJzDzexL03/Ej2xuTywtoVui+KX4J
1tkSKQIaLyLdy3TEXzSieXmdgxGjUzi37oNCpmLjPL5aafafYHGupboLxKGVRk8sWVTdLCI8niaj
RDqm9jsZrU2bPWQO1aPOxFSNu26HZOkqkTm8Lx5Z+LW4tV2cJyjLcaGJVfvbrJ6ctaBcIaQkS5LA
X9ovFUeJRNTGATPT1xDCETlyQHLktrcQQKkRlWjJTPKGDDho5H2MP+C4JDHClSYPgAHX0Edaq/CD
N+plleqUdwc+iyewiWOUWSos/FYuaqKidMIMkJDpH+O0NJs9CwQCiT0qO7VGOkabqmCaEiorb3Bz
tD9IL/jDbvgHZ7P2qjUBywHmcM4j5cJ/5DwkFhSVB6BmJgOzsOfxUb+rL+buMfFCQA3VUIE13Yqd
HruB+zbgkzG+5JE/dWXuMlzBYpk8rEAPhOXOQa0CPq4QAaX67t084lrIzBSjK39Folba+AJdyDva
BCHwzWRXBMokwwDhMcmRzte1sC+2cLOtOGbW0Vfu/s6yhqmu49xE+5F6NhXAJsNII8VPNb+XE072
L0zUMa3BwTodhUUdtckb7y7UfvVXn56pzxkgem0M1KMt0EMv83j302cL8hfS3Zo0klJOfj5i7TNf
LGdyMqEwBQFSZDCArZKrpu3uHCjzaUEladqT87w1q4SPyj5zFWD+1BwEzbwI02OEGho+P5MTobp/
HbeLuh8ErJMbQ9frDTUMGQafUW2xVCz0aSHmmXZkXbICsZeyJZ3MD03eQw43TXESXle0+zwocfCS
cRE9fajNQwYRRfBur9bG8cV+X19NJdv5ej5quZ9FXqD7x/D6xX2mbLVU/PPdrSCxnjhXfqI2pFPN
79+u9UNRH4+RcnkrilYOP0Sg//iy76kxuc1q4pKmRe3cM6outsW0ca5F1b1pFBHsvAkLZpwmYcE6
+ByuHHWQQmTKJ7AANe9VVIZeZQrfFssHgQON07MNerWgHDTm9cRx+Xn3HGwU6zeoi2eqJu8XMzuL
cPmpc++c8GHCfYVZ41Wx5FVHe6BwDTI5mtDqtSeoCO4vYYxd3B2IYqkB+Z1e+UKoUonZc5NGWkJx
KYGAbKcNocuvLUYgF+hFYp0CIR7FYG1uSKqtTDDb6h5GNjgwdR8R22YxWcTroKfR8I9xnIBcVXYD
qeZcWBahP7JZayDL8H+HTy6WCbF6eb85N7E1zYsZGHEYreRvYJRCufnqZ5hiyLvwPrM6SEgkWuWM
BLxU4syVt3wW/Xdl9DlPl0xADVESp0fJr9Kn1nnCcyOFWySphm2ug3UKX0ZrVKdKJeDQBZ+lnH+Z
G24aKo+t3d3G2LPIIzs9sj7tgsozpLZT2p62MSQb+q+MvbEivvFFjOPKa5dIxiY8sf99ZWKzNA6f
go7fi41cs2m7cOoftCQyphaxH01RMu6wwtDz9POpmDDS6+qrj1U5y3S/iMT95g6wVcNcG7DtETzn
3pkq47TJ9x6fSds5Y+qWaYgXm1s7DSmpprySiKxTQNzwcEpNHuI6cVcY4u0o+Q5gNVBROl2uHTbd
/cMem5qMfiGtkjarV/DV2/qmx2wDtlSFCJBvGP+yk96osp2z0B5p5k8y4+q3S1SpQg8AGiX4216J
pbRe9vhnWvE0jwa4JH+jo2CKUBrpDAni1df+YfxH0UWAiGp4V3Z2j2OGj22w/Y9t3F4EsSMGiTa7
Mu29y1MZf5kPKOvNtgFkI8ROHk1Jvuk2f0PWmM3TdahL5f2PFdadtXbQVzDUsrduJdQ2EVX5p5Ry
KkU8C01qoFrxWNR+yfMtqrdwGgCv9n29TXMdE7vrfu7V/AvfzlalIDLv0NeHjuK4yCjUESSq8eXW
gPmGyvs8tj+iCMvcp7P7s53aBEM84tzmEk2jYzIpdaNaMq58I1AIC7ZyCsMNY4zf0uFb1qs0Xw/E
MLArWHp2z1NVeicyWPHNlO9uS9VLEw+tv63T9IjFZiXnhU6cWfke5UOKFKN+obC8Ivk3bb/5NfdI
kjFyWDy4dcvbjNYSOMb2Pr+FWVDcAHefff8avY6JG31yDfxAXak0PIV7MhDZFFIp+cjsaCxl1QqJ
rKx2sKJaj0DvEuBae/mgeHQqaD6vTpcsfxD1d+oJSzXeiDS1tkw92NsJxmceprtduBk1ValJ0F1a
lkKfrt/yNZdUmKbfiTymWSpsKQFckTxMpqdaFQ/LJfL77Xskz7/69R8nCsKEdleNCzWyO6y3Q5go
aKimlvzGijrAzAn8qwj2b+APVJb9BTz7LFDfx+QAk9GiHGVEzThjx778cvJrM9CmkXm2XqdZ38ZD
hGZw1DVmVkkd74fP0+IszId9erVRrV2Nky6KMxFpsxiTzCAfWN3o/scUByYEjvuTbl9SbPdzkoUB
GEMNXmUiNswCOWCZbX7XP+Guk2uPt/KxRMy16hrfSfMnIA7Zvu20KmYmWZ965ZUlmfWHAxmHYLQ5
nBxMj80uSOHqOQZNcT3oyhWlmDexkBWoVAYVkmfla/eHtrTPFpMPrjuQQp7H8qTbusLA8c8TafWS
+p9gNvX4ZEupIyIH44kp2SVdX+rCtWRrXfTGNXACok2NeoB27zf+gg1n3B4pkGllTNJtPbAUvu63
Zzl6998XLsP+0Y2e3gBHxjHXMm+Ejo7IA7WPU1vP00whwd+aNc6PVY+rWOX3si0ELXGPN0Gryykw
+/qC+2DZq7+4O3/gqgUah538il/JKrjWJlHig4ZNpBYPp7lbGGWmwO5JuN6HFV5dPozedNkUqCpE
CDMz+pKawoKZ80G5y1aqQv2+H9+UbGUhxa+ZjPd9qbohYVTVkQguW276v/e2MZNkCfWMeuLZvPFD
h6RdKy8xOdTbLxuZyMEg4vBcX72mamMh5/uZxGpLPFN5XcA8uR2Z9To2ookv8BMzXcQYbDnCx+Hj
Ehvqgt/2i1VVw0rKyFg6jMo+Yeuw+MkB5jBvwWYgcbgVLjA6BuD4qDWDAp3sCZZRTw9c/F3XljwO
Wf0IvF8K29hC7o+jlRVjZoyG5tG8NFGgB/xldGg3M98t7GnX4hQaotPEbMXaA7m7Gu4ljb8Azyk1
s9T7VQc3XWgsnatZ8j0MCF6wlBxC8m/DuddUwf7nYThVizUdrbRWmAXDkZhtGW2PZHS79zcN3yYZ
kHt+CBLGMKzUJphxrL9sU1yaCe7tW8CXJKh8f5e01vI0FiF1VvqnplhfIJ7NXd4jCIdZ912/eSa1
5sWE0tTHitt7Z4Em6fdEEI24oRo5W51B+z1Jad4dQMbnvI1tpeSWHwGNwyukVOAnP2qRD52lKyvF
W7xzBDtif8cpX/MGLYmYsgpiOGGSujVySPbQxqapjskJU8jbGzHP16XYKisQVSjqGYMR8h8uWJpx
IWXWSKfLyOXriay3VNqrqM2nh3w+oA7yaxShi5HX7ahnzelKQexP1HhfSlxvHAHn94x/jt/SZrWG
/9fjTEcr/GwM0sOLlD3MfZtk39eFn92x6AK136cHwOHiLYN45Wwc+CelPTBbM7NlUJMv7rMl1oHZ
r5s2ni3zjrTEAj2gXNSOVjOZ4mTua0AWIzFm4bQErkZUP1badTawo95QLccS+tOB6C0YkNoVXOiO
itksS26bXdZND/MZX+dTTbrLvJ6OnrHUWpADXCtExP3WZxidrH1+Uu2hSnW40nWdpcn+dtW51pb5
0jH9FzhBLMxDPvGVxQw0g+o7lHs46RN9tO224az4kiMm75C8vROAcbzfim7pvvDA/Vh+mVcSaRks
MMKVsWTgdMxCjfXsVrch9c7xUX3qGv8oeHEj2NtTo43QOSpiYWGndm/dEwg6EdE6io2y3aIofVSB
F9KwKCrySuLwFZAnMxmf424P+lIvNf6mR9SvcR1y2I5ARBeufIxylCDEtH4CZPiLslgwiLGMQxV2
HGNSzPYl6SMjeg4eXPpxzuU/oyCAkflgd25/ITnyQe6/yQDvwB5NwhhJWyrfqJv3mJaYnqLyp/KU
/EDXwoFfYlQeLDQCwkVbihricWHMhqAPn5ciVbSBx41gOerIVxFC4ezRo8AU4CgRiiOvYnZia1ja
8G9dhzHHFc5pgA6IhKAnuZpp82NXTNVf7h3bp4M9LKqmxSXcHRRMkI7B4v4b0jadHp9Lb1jVk9BU
CU0ExgRkDlUq1ebUpCfTckkPwXhPa31bezzKfMCjPKRqrmuY3YTy64a0rhGCg8AU5g1fSMUlZjX1
Qp7ivrZt1llKYz4zZudKy7JRfe6lKMFmb0BCLaiHDAD9GipbigVk5SAYjzbQTxnreLMVTZ9+Mqrf
3elD5b4sye8F8X3pxzOhhFOkr2WZFOj6QZ+x7PiZDBPjkCQjQdJ4YSeQzQY2cQw+gbmjQm6KLq8j
jBnkBe/db+GYyMUr0C3iRRqtM/9NjStqxRyEBL0Z/Ad4D/4U2zQJOl7rm8OnUTEMkhVVL8Z+hfRO
+gVbWZcZQsOZ7I01wvxZTmjZKCWeKcdXsns9+wxElxA1+NJHh1OrRS9bHOa58hpi1CETre4KRcqo
g7tGNNLgIvw+f7I+0CPdqg+fsB9fSmCER8ACvPbuMSRWYJagPABR9UZ8JPpxMEtjxTWJo5oUzdQI
Q2xWNGpBZFurLyyRHd5CbI+rkQF7AHv9jQNf4lndxDcqHyi0RuPb8D/RXsOuXJ/9ahwI8IjIJFPM
6V63RffgHthlMr7Xn11dj7la66ILE3CTElPjrE7FglZI1rTwAbmQiqtnYHsWG78KU5JufttZVBN1
icgJqvf3kNnRS9CYRJdJ4BzIYyS7NsQ7szEy1hj8MnguvFXGHIbzfwXRvW8hDgYct2zandfmEYD1
YDyWvhobWhuMJehLslGI2+slxdeAwi9kj3lvCPDCO8ePf0VrKT8AbaHDSmzzgymXPaDnOnI8ctyC
4fynoQwkJ2QZLYKFPVHiM7Tc8akVwp5C7oMOy5IOUldq4Rr4fgpeW8tzAUMYvmq85Wkg+OwxoSVm
69Uey7VZSyo8Db+OBBvnxy39Mny1DEg/LVWoLHUEFIvPdqzh3EJqlaNyrjsXD7eAJUXFRpuXHhpq
g+lDBaByq78GeUt0lC+RKfmO55KY5ev5FngZstTpa3KA6R4oMMRrHhmv5e+FABxjUYK8lEty6V5B
sAUjRz8+5hioZV9sYFHZoP6Ctd/ekYivJ/FPfKbFpQWHg39LLYWAs2mieACUX7Ln3GHn/87goX1q
UJ/O56lT5Q4xo2v7AARXgJ246rT1+YquNYVtjNy7Wx2YKABZh9HbN2DWQqCnTShErPU38PSQkBJT
RU+4JWxZA1DYbKOc8ZcD1XAzj6H7xDP+UgAwA5elKXb6I8R6pr9xsGKMvQsPgOCeVP9h2wNEVt5U
9mIt6+bl0B15oO0CS6/D7VfAAV0jL5nZWp4RssOt5Gm2pFr/8lKNVrevCYXJ0RSKbqebymugSCYG
lti1lMjA7uUEu3KgoqWqPof50C5Yeir04aunq8xIlX+N1rSOEWaBC4jHS8ezyoHTnhIpd6Yum7ik
DBcB0ToCo/vYqMo70YkO1+/ZZM1mce54PGMHhv8IhS7SOO9zWxNtPniRhw/KILPQl/gcoDsPs4pd
4MwVOSajzuFYq2TrC1zlxaQPGhHTQ9hvcYdMCXqu7xjRa0K7zBoGn3WiTrjS4yqZEACnbQ1e7FJT
1CCaes8KcxIce/Y30aMAOlbyRxp5FO2sNAvcNhgOLGGxvlsfq4LqpI/OCiDfjofDuo84CeQHmp5O
4ra9Tfgjh/Mj40icrQjfoAix44+GdU1+6aMXvnSL8NWQ1KMseNTQ2/vcuRbXmIWUH52taDnIyaM2
SDRdjPm1XmQIYi9up5Uf1Sr2KqpkuKJxccWA5WZ9M6xzapuZNiwCH9Qak8qll+/m0I5pgzs0lWbU
3HS9s7L4SelDKH0xMwQj2JvMjmYJTN2G+iL6QOLF9dQr5Mcav4pp6Ezn21BKF2i+FUAFnkxnRRKz
NulAluJWnGikzXk9GADnQN0CTz3HVFa9aoTUMmtQpn/yitj1uIxc+EbOCfCHNmfwIzWLrdISmPSc
a4xcpwg06E6YTQhwN/D8kapwm5MTUWDieNoP3D+QGWJUzPxR3Yoa3rPMcSV2u8S3lxdFbsuk5Gpm
6brEqAhgt01d97bXpn7PsB5Gd0jGjhuALBiFdLMSnyeLNRKk0M1Z6s9oXXmFQYQXBQVHJdPAoKyb
uPrblBIdEmAzqkMQc4vyznVrzxYOE25ioJq8+RYVJdC1YSMhyMRbm3TXXyMadvw3FaX4JHwlTXmC
lY1qga6fNSa26JcJIn0t92k1IKof0Odz3nrc8IVYJqBkgMNRub/b1hS2iZYrSTTYFl9V+b27+OxL
OzQWHewU5AU7GLE278t6V+IMIXl0xpJ3uDPvt53eQOOSIBGBPQoaNSlrdotcs1exKW6ipzrQpM/Z
2f0z/1v8R8lNKtPqxDUgkJZVR++Efqz7J5lBHxt37JYyQO0Rzc0dZszSk3jpmscXfYSzBMoqeaJj
m8DnD7CJZGVjUeEUeUHAZYzf0AiwwzlesyRmiL76PYQoOKQVnCofsPtgZJXvYuH9eVznf9GtbyhF
3UCf7jM0PXCKhO9SACXNs7j4d0pKpbsF0bX046jdsJ8GCzV+n0iImZxGG9MD/ThmzjnowOvEqVu3
0bMedUdyfR9r8XbxbLvNuxsFICfGsj0kuoLqfiuxtK0pGHtIzk7gYZHZ0/rnBvWdRA4RBk+UB8vN
2TzfT3CTkwUCq2dHgWCAykfvnPfztaceVYuF/e27hbH9hi4WhxKqEc8521R2213CLBmIpDirbF77
iHlKGGUNqJU7SWu/RTWs2Z9UKhjhH6uktc+030xAawVv20gqC0iXwzHWqRk9GMZXQhxvanWAZtyN
Wa+gLRU/oWxe3mvKC39kKBNNTugZDLEoIFXI+tMLHI8k2FRkKbJHCI3jDEwP6NLi3+3s8avDsGtN
lVsHgdgNdXTdFKK/exdkIjvykt7T7UhFm1tynQn/7p2b3JqGJ7ZljqW7w7/I0BHMYJ9d/KY9ddcb
L1hflNyJ5F1RNWSDm1C8LqEViWZB1jpCkxTZXR8vALtWwu+6SbQguHktQD2NCwirloNpi+kljBRy
QytH1vBXBN2EOfnXelwcE37nzr5kvqA4EzE1WVtUF+2xBxTPMn3P1Cm1kvlaNQgLtykkER3WeIOp
i2USOskRgMynoi1mzEBVVNxJDbGYAj0JfiOkzBGvoT7U/3fbhc57mKmQxwaeRTkG6W+jMWmmLsvC
v6ZA5PKfWiCY65httmjtZo79v6BuWJJEc+xhCDw8/d0o8GLaqKi1hFFo57q5Jh8DD9kP3KMHWnDb
ajWzEIQtsPN1c5meePH4t98WbPXxQYzwPa0hQBglHM3Rulb3g24tyjFyD0U5c/+bpVULwaN+89WL
Zw0sYoRo4b0NxuqPxSwK/r6kxZrhz8PMk3d1NlApPPFL1WJyffMSoYQ1ETwJjX7ehCn99E/x1fTu
PmGWloJPs8E6FyJyVKeOA83QEO9EwJVvHRDkbr1LfFVz4i5XWnYmE0pjO+oAQOhTIMx3uyKA7czb
buadF5FGmS5sid8rStL4WmxW5PLZ26vKhGgTzk6OG3eHkTXMTVpInDJV7XPytDiWOxbmyBEC/lfO
/fQ10rLH4VDA3r3OXn8J34qeb8K4tSvAppsLEHVd9x4lMU792MulnFjTVRyd43zNJUaahugE/meh
XElJcgPQICMBipglAYNgt0FpRn0z6TY3HKsgLlPUMBWfoSG3WmLoScVRtIh7Kqp5k/e+E5cGm9eA
jEi2GaDTQLWzkRyG8xzW42XyVTSTMptTO4a4WpsiOQj7/ITrbfioNLBH1aMjk2G2xlxo2LW9ipvn
0uoUwBR0zEdV0Ow7YqVbwFv2unkfv3zl546qVEcp8n5maBzrWa2hcB9sfIR/MNGPqGnvp4BM+rx1
bxGThPJC3FoJ40xf1FT5NcfU7xBTMdKIIbeDzeO5BCoOarbXyVNmfI7h3Hab9LSga78jD6iB0w3z
lGMi7ULbA+SLqeDSAFuBIz8V2/52G/WzlfL5D7BZI3frEudiwU/DHH+ilXQ3RA+HFy4gxMjlcVHN
LPj2+KwECBagN71psRU2jnX5vQp4WE1+jbpuiQ68MKlohl/wBZVV/D3cbweMdq9wDoEug0y6zsbN
3wYCC8Gpz8l+dSVCks5eMIXlBEUKT6bC+erV0FbVZsPA4XcrSTX4EcqD74lW40V9EHY6M9SyXgoN
UGM4XMknNEKQrDrM80R7omZWIMZ8RDR+mLrVZioJVQK+C6mWtd6BSptuObyg3VtKLdL4Eu5dEwNa
qiseXV8rdicAX+8Dg2/e33+Ud5wzGvSJqqPQd+VypX2olkYDHuSW+iN7GxxeBoLvGemRBlOz+vs8
scpZ9NFRXnjyR3CKULJJgK+n+JrcEFH4jVDXiY4hRWpdGQKFR/lfUXcg1oe7Tcp8qzxjNBCuATml
3ovMZOo2vbQ4cQJdDpFpKFL0I1pNZBEBr3kndIbqWoSVCm4ixPAMQKQTyz3I6G2fBxMgxCkbmKAe
sLUBanoigaBilYRwpL2SwNApldrL0fgXHa8kAwigZ1Kx/kaR23IBiiGEaaA7XHATVzaSUImbjufD
0tt2znMkyLCYgPFkwgba3tgDiliCibMkqBYv68KgKe0N4R/sCj7rBQdFenxFRzkrnTmcFuhA0/41
JAhqnHcZo3TFLetqcCsYBIuTV7ylXSgKBCk+qUXVrvj/IXgPNs65Y2aLF57LmQncGaZLnNGoZTpe
uPy9Os/HAJr0CHqa0u4KaFpk3LVX7uNQQeXbXiKHowoFJJGkayLB0SGG1/uWg/koNAQ01nwTpE3G
TQAVbzB14ShooQD728F2CdGP6ZTH8is47rttcKmJcKm5+FcU2uFagodOhIkg7v51Be/VGNQ295uh
9s4GA1I9TURugBkXbBCkBXM2VYNbjrU6URZprrO2ziruJsRiw0vGWkgaOmdL/waFKgkxJCOfU5jE
MRzHKRlPIH2fy6oHW0qJzhJhMtMVEN1BjyzxvrJBY6Mu6zog6Ajw4QXwnKLLHF6eHsIvcrmnsGss
du6Ht7B0CNfWc+2dEJpJjDNvcpJ8isZiHaySGPELtuOjI7X5e5cuAymzUTYE8vYZYC75rXrPsUeC
t3ym0ngaVqQ3XrnRWNx58xGcfP+coPiVIutlkeyBlrX0XQDwlJ+G2xVV+gM9xgSjYRzGUVa/ZGuC
GAz98aupM6n7ZG0vYVB+p8Bq9/tyHNpPhvS2qEWOX5AG2OqJou2CuukC4Zj5LZx/fM0sJjfaYXq0
e4q98NNKTHVs3dk0cEX5JD+sP3twUl3e25ucxLsWbOEBYlddW3e4/f0l99/vBjus/2iDef9jTZdQ
RydmCk8y+tbZeZ7LUEQ5VKl8XHYeaQw7QV9n6zJvMq+8o2OazfFDqathUCop8gMEPZ4aHCbtg0zq
OZpThgN08vfe4dq/pcJYWQwo017EBYrKMk4mAxKGBT+b482Y2sFPUHEoFYIxuql0HRaIVof+oMz5
MAqhUQTx1I/IhROfglktLMcej85+o0F2KYS80IaIr+YCrr16LY6EvuSzq8Ze6EPw+x8DDkA7TbMF
IvuA97ET+mkBiKEL7MOU3bieJ69WrOpvvrA4Lj0+6+655jrr2I51ISt5tumsPcFkpt6I2ZRs64yZ
hNO8iHuSu2Suq46Dwx8WkwhTYp4aqBT+Md6En6jIoNEDMlhUNq2bIyMS4JbBL3NHvAJMXphpYsnS
8z86Bnny3oVoMDuAyDDh5gvmIAE8Cx4IeGgR1gJoONtbVUH4zcfyzh+PrP5g3zXO3KiHFNk8llwL
st/3xXvVvhdPvFm1pq5IWiROJ8Rqw6UotT9jQIe/3wBryOS4GlKWkQDKzXhPvYdnT1HDy+N7Ric8
rw4ndt3RtXVlz1OQZjVD4V+lYDWaGIXiXsyifD2uFbBHb1EGTMj1MMYo671A6bv903+oIM9XrQB3
EwcUZ7Yb8girFCM2ptbz8D4wKL7AG+3uhElFSPSe5ruUzTHDlBaZN0ahId28c9GiQ3ohHT4RDXGe
2orDKjBdSs+1sHpAsSlTJh/PV0EjCYIgRNcWu4pcvRJiIqTJU/xZOtbJnPTKrJ7HBXcvMh0QK4WN
f5hFx6bLxSvxO3pVH2dBLGi2+T/jvdYCmiKLRUW1Q3e6VFtvDsEkEpmFtrwcshhGww5wa02sEqk2
pImgKYoCCdas/GYPFhHxSACrS6GDBaD3VnoIlzYoHGiwXSDG4hs9Fw8XmKnBoNBTz+2GCcRf7bsL
iWy3IoZB4NkBMEWZXQN5pQElnNOt7vt4nYkAOxZon+A4jmqY/AbG4zbwP7+kebTkU9U95p5b2TvZ
TKNMhqcARD/4oTMiWuM6uPaJAScIbnqREP9LsW8jBckToOglKt1JNl+EjuZMUJREFl6F937medYh
1k54SaAVM9CFuE/H594vWoiEWPE185ih5lnBo5oTRH/cGR9Y9jUsVUKYnJhaX4wI31//ohnndGKl
h8FG7zTbn1pggWEhWQ2cf2+agr6YJRme+uzNR488FldbLUHehc24MjoKBM2FgjIk7MxxrHuQH6N1
xFh6wY0TNbwIlXgA0AE9EkVEXxHAYGDImuu6DWvo2jcEFRPwZWTGYxCXBuYulxY1OH3lEpUzy5zN
PSY7bHjlW7lYLmweTZdVXAwwbgc8ZC9/ggm+naPNiTlxlJ92vpAJgmyloD8WQgG+FdZOCtUUrdY7
qeJdzeskm2NqzxNnTmU31VE0uvkqo6jASSOpykmlpcEk9MjU2SwIQePOSfoyvCW8sLknXj3rha/b
4hXAXWgvxR9o037PIitVf9QwNItFyFx5c2Ml2zjeOF7LKcSUrf5nw2qdJLFzZ6mxXEiqS84IHaut
rl9fhKsThYEfiqCyFpO4BJsWO83jhMFIXbirM9TfHdrurf1SUsBCGbtNSvq3E8j4yFS9dgHhvyM7
b4fZxXi4b8tWT0P5sdE0tA9PM4prDwpdTMRpLWHbffJ38s+jOSZNwbvtbG8/CHjMHzna+Owlte7l
n3UrE7SmkAUtpo1U9Zyu3QKa804oHXsrnbE5zBIlnx23YkL59hh+SGvggbZNXlJcAJQuBgRrD2xx
XuVHiIMpNtBaOOf7ul/g2qS43l6HPRav/naMX5pWP8yxQJ0ZVHUMZ5ire7sJJcomKq/jCJwh34KL
x/p5vRx0KfQiatpZxfUa8aQwtVUWC/6ugYRninkueRwPXs7SfhplWoGfxDlYp2gak4MAmF1YRjBR
RPD8nSMzqw6U5Ijj0ZkdR3861eheTcHYCdVJqPSQJSlBs1GhNzJ88W57x5HgDy/1pfsYM9A3bqh1
j85kjkMAw0p+vWHuFebvQUOFXm2WOOEqKcykRfX71kLqtAFdMVxAQVPJPibK0C2DNesekMZLSfez
RFidz9kPMi06XR8Cfw1sLCNuF93sivO0a7WmVMD0YAQJd9w01ggleqYp8byL1CHvRztqz/S7Ic77
oozAJTRI2B1qXfevCGqzlelzcxvq3IrikL9lPTUE3B4MvF7R60DI+lHc4JssQYHfiSE9XtTxHJ/7
Yy1FEQpe3UsKDonskc++ewIZrGNTfVCQ6JOU8Tb5lkZSlJzqssg8pH40r/DzS7hlIexW0+7uLOfi
VejR3Nxw/ltDznTmlAngHkG4tAadLR/7l48coTKEecnYCpyJH4Vlwo7cWFNIcEG5L3tWklcoiH+3
ous55eOJAFQL7+ENOlRBzJ2u1VVMQoWvXswSh+39groVlpghgfYziVR44mzkF/rCXRA8nghs27Id
jEnYjfuV2uAc4qKqny36boneaQy3uwMWc50J0ghpxxkQP0GzJpVBjumDc3Tb5bvE4/kjJ4tX36Iz
mRxwSTJx6VOOkhBzk3slMiGkwuLRdSocWe8beZZNpYlvimQDKhBvHxozrl18oWvofOrvLD0TFxHu
3t8vnvypgFWDyQFCubcbs9uzMEmwbMAni8gouOMYB6RfIRGH1R/ca8i1FnoTEfexrMDYK/dG5rr2
aKjxznLUH8egUElrGLiBuTYLloqgIVyz6+tcWsFhoQHxPWeB8Px5FiLreGX9J6+Jog7nhO1stXNn
2xhWbTYSq6FdIj2WC2dfxGFvsTNipUTgXVz3GJLYdbXEaJglGd+xuJ0AvgohnuhqpD3NG45yRCOu
kWfh7RwYPfpi3eu6NUc0CbMNwoTDfAcRhVB+OE5lCtLk41fGeJDAkWaK7CyNqggq3a80E/1bPAg/
Bq7DwAHmsFIIbp4jZAJxU9LDi6uWmtst4riWrNMd8/3gpQGg5Yetybe+xvxNFqyoynLsba7owl3G
l+gJeUprwr4qNrfrZPqSWRQjKo7Brs4z+pyBUc0hGyg2rK0w+fYeOUFxnadPfIDIGxyjCSva4yXh
Kd2KO/rm9v+UpvYHX7Rn/nm+CZEF4r/lviZtdj4RkJTmBly9/QAx7KGApJEWHx9IvawUJYG0zpqG
ZI1NmE0G7QzhFNU9XuojrHgRqCnK6D5M8t9bBFFCByOJw5Y0Db2oU1iLJOoSfspmDtxYjhc9sWOv
bYHD8+Vz43mOynUyjPbxK1GhjHu/OhMbjwOO9v9YjzaGQWc3suJ6GPiASMqzykN1R1FS36RPpLGZ
HhyEluHRdLyES3HnYWI9k41fw239N3gxB9Nw5Ge8rXJNNwFn0KvmjZaYhmFnc+OLxnIN2fKDp0SZ
/Js8I0+Gtchvnb6s3dxFekSozsQi3ULrtOXeiV2ljlDmGexqPTXh/fTer7nJcwuXnTnKep6IVmuX
gIrRBU0rWwYIAw7JloEslIXuOH8vg9ufh/ZutiT3+rCKHy9wYF6CJSt72jSRM04aOfsL8vTQja+v
ErE3ojUSkPCLOXwMmzCD9ATKSq9sCU6Rl3dy1ZE/hziJkBPvkVl8Foe9EiKfk87fNUUBvoOsIq+2
meUsUGLjRGOYaPyj8kAu8Xqi4s/n2S+qki9s+917VcHF+Zy/GCUJfEEkZPsGJU+Izq+9LdSm3h6v
TiFNdUsvsRWNIipBLav+dg3l7x95x3+f6f8IZISLccLUfZH8izFi/RN2uFkMPY9GZ4Sx+LCsx3/c
imarcol6XNksXnKtw3gUavE4f72/LoSPMe0dQTaevNwXXnSou34ttjP39BbIxnoiqbhnEtsJF9IL
2prY4vieesPJqtloaQo0+bodKairZX3qjSn5t9776YZ4O1NUXuRx83rAuvALr5y19b7W+PVtDh11
TZhnrQmOXkM03Vw+wPxCXjB923CUfO6hC6j3UV60cCb/u2VG2a5IIwirwxvGP5FphMSIkZZ3QN62
wDJIYm8dACBBaH6GBrc3vJelIvvq6dciqostDDUUpG30jaD1Tu4IEsiNx0USr+I6ZA7TO6NDzUCb
WmYbEmlwD+XHxhdkgZmLz3A/ctnkwQRqG8gtTFJHdSl8XMPZDt7TpR9ZO1Ktt04EshDalKy3n14Y
n5pgCMomFn+lEFdgp2V1TbKpdBFezOEWxgv5OYvVGfs4JbKhhu+ZfRxD6WM3Jm9NxzXXN4SuSLq1
HYOSCRMzq2xyaWvWySxbaN0gUGnVMLo0iaIgFBIvbodj7sUvNhshxqsDgfTddKqgYOUnQd4Ssyfm
LJXcDg6UY90rc/1fZ8IbvZZv7R2of52Y2r7dMwOQUznnWZEYPTnIySQAVZzdoPwGljV+WwrcKcjA
JNMd6xA/xKZVJji5lEIQ7oNGhQUw0j/mVjAeYe/5w9+JEsKKItOsMsZNxVgWDvGXtl/8XtPo5L7J
IwbkutG0Oku58ChuMFaEIDftJE8xHYxk5or2jkFGRFNjhr84Hw9Sv/79W2xqg32GUXTRGPBPalzc
Co5beZMqqsXLqbrBot0Iec5KnQdtZgQwn45Du51/JT9RbChrNS1Hx+jWVQNfv6T5GDnCeilW02uj
YxT3/F9agprcXBZ8b7IbLkjgFG30WjVSd3VKr00p2USHyrFzml8ArnN5ZC6kxUDEDeNabpQYXFvH
jbegP8Avu2ZBoAP/VW6xtTM9xIGB1DEZbmrUQ3GvI6q69325dmqsXY1E+09xgH7r8BCqmqCG8FmB
OA/KXiqNJMrSQcwsGLFF01pB4jXapgYL8HaELVWEqmES7XicwuA/L8aoLevKsXYSs1BVYC8tifMc
Wi9VPkwDDZTmihDmuZsgF90aNzgMgzMxmJSxpuBnoN/XU0KNDyLtng02OuvtrKfbj4KKvZLQaF4L
SFUrxFQqjHCqi318od0BaAbQBu9WkQE2gXSVwsemVaYG8ZsDeRjnFPGCjxJKIl+VaT6w59e7X3iB
/Zza7UJB2VWjJP3sGqqyX9xMpoeuQQRQ9RKv5vkC2QNBdYcguW5iDr2SlOMUVpNuDGDOtcw7YqkN
4vj+WUHhItnAMRX7cA/4d1KmnUbeeoIeuyk0eAfVkIc2RBYpqwsZHx2k9P36JOeQK3RA0RiC56or
RWuuVuxKYfWQe1L70zk+NZBJvy1fXYGr2nxsbzfoiwK7p32yj0MdK3xjjXmz/MpVZ05OEAMSWeOQ
sP3HZJXS9I/rhQOjhz03o5HopSTSYFI2heHRimWhEvLsQ0sEfswmq9RjRhWhNsn4KuTSGjlgqOH9
SfF5PPrFeDNJ0iKs+I73FO6KNnxeyZKwk5WwNSRfJyK5SXpP2bsbfByY0W28ISLyEj8NJ4yJWTb9
FAH7+Nlw6sVW2G3TaqMKhuOMPTEpQTYgALovqW5tMpM2yl/yfU53PhrMX6klZhtxp7Q9GUiksi4a
1gt+7es6qhz/1u4LrsTwBvktXUyFjEXQRsVv/FcJd6V9q+DOWQQ2wkrak9QNiYyZMapuCQVU5s0Y
CaKxUbyLJhuNP0l8toU06Uc+XbCUovZb4I2vlQlfBzK3A9TIOgAUB4WM22wCN8LgngQVq7SGU1CE
GohC0Vg2W1LpzAXqecJse/R0TUj3MbrRix8oj48DkszGRMIq1XGlsQQxLRlMBeJGG2a4rSB+5GKb
IlbgkbX66mt7MgUx7uZZjXhOGJqh8t4j4/fDnUfmKlM4iKwbQ1N7ka2j7XabU4bODVgsKPVpQFOG
cXg3aviZMQ/p6Z9s4w2uF0YubcCHYGZdALdt3wf0jjgzKjgwSEQ7GW1xxx71G/nKRX56lgeJG7fy
LV01qidCE0gbGbPNnr8Y8yMIk4jB1zB3bmlXmetXuAS2CrdgZuOcKfOt6/BWoKlPgTf5f/5E6aQ1
+y8l/CBoyYe0ZZMEeerrtVP7WX6QnQnsG5aJY5MHU9dXyRzeMRGDm4/KE1O+JsuSXLiSXVfobexY
jCsMlSUKzbSDUXihiFS1QF54q4irrgOO4bI5Og0Nmkts7OuAibAf75S1uqOyw5z8Uj9JzosG4Xjp
DivUkkqgtHIWEBgheLXtZ71IHjA628BmFYg4ETtwXneDdTEWgp0m9DaDq1ii9xNHqcxpaKUn+puu
txWXAeKKubCWYSsFMO2xXWQJP1Ls/yfWE9vju9pKP8LBO7SY/RmsPexJZ7EPjBrcCJqVLUM4GtlW
VvwBTE+Mj+fcV+OlKLTD9qtTV8ZkwrSuMzluoBUXU9m3rIrY6MUynW6eGG768uFOB7yikxfn1iRW
V4X4CkgCGFMl4MRZWt6QUxWZF1KoH594DFHAvn5uAs9h7l5NVLCpYDzi/e2alt0Nb1mJoDwsXKNr
tXq//QdutfWpWDV3kyyyDqtDtFG+q7Z1K1WL5Dz9EXQwkXieHaCJby9Kb8nhPstdT9rTFM7VgaKY
hWBVJlHD5zvbvTe64YCaMkxlxos1gbvqk5F3KjYAqnCu/wh/WAOteYOaJT6SnzWqQWJeiPfZv4PE
RtuF0RJfEXtWMC+KgEy3wWlKG1HrX00PNSI5nEdSJK0CKbP5AXbd2del67dv/dMZYE/gyaFQjmUO
Puc2iRMV5MsobFQ2aGV4MvD5wxXGlCUY28GvIFC/OFFkonGcFoTRCCkGAVRj1fbUvUMv6A6UxODv
NWe3VSwaMecTtnfjjWz0hn+zmDhNBAjwVMjpxHvpZFyENKSFm7n4UMUdsNJhL34OCX9jX7QusC5y
cmfCjg3iXboXw31SAambEs36+fn913GBL66Eo4VYVpPeQJLjz4Ir49+yy54worZAGDn/UxSOTUJ+
6WS4hmTXa0yh9ExzhMVguZJd+KZk00ky8SnRLRhC+nNTGmaCLDDQFPFPvqqSblR041/Obx7xuiy5
aPTzeyYIfIbAE1PsuSMAlne1VcLtgVkH2kQedU59/4/geTNarlnGgIxHiAXBsHz97loDvtWJlIB6
FSSX74FgKMROYrXF7oA+2UtlLboSS+7zDSygg0kjNFe9u7EGX86yR+FEcf/HKFsLY5TZe/Qhcfz8
tZngwY7qY0GFjIV3RYqjFaqNI2IXSFzbsOgWK3X+ala5USHCoQwvF9hd6YmfPG9tW9zhUJHCZVCo
gcin9HpT6wgM+Nk/8E9HAGfJVOoXwqW8LCGwAurGYAqk+cw3CGEXHCg2S72nWK/pIBiuPkqyVwFF
bm1HL0yaKNnFKrjFdNcWCpAegNr9WYPnwLOOQ+QlpI9WAmVHlyHKMhVbyBnMz/q4B4zrkLT5yOzU
2RBBzKbVIDM/Uz67LL0gtbc5fxFrl2BDYgXpRWlCFgxjLQKFp/A33qEkCNhU8qjaoIwukO9byCTy
l799NpS+h2UXCGxdftdbowOwMX/8UnWNSHdsrM6Ve4dxsdaMZ9YIOTl5LFsNNhT51GjjohoGnJPj
BT2ABlCcCCRkpQqTIdEoa0UMVw8OSA//O6/URcuY/h55EOBVu4s7u8a6ljJTVAbNibURCYYfhNZo
oZaQLBPYLuS3Wag6MYVeLjJq5YqXddcuZFAFQhw53HT7yeasYjhm7QRIDt/bZZQD4S/Pv97NwHx/
txw3yiMKLpg+yrSx+QNPR6CXrk0zkJ7uYLGS9dFJo5ifdbFIp7l+w2XNDEAxOzLXMQnpzH5u9NZo
00kzcLW0olYv8aFcy1rv5OsL0aKVr7eb9KiF/u9bawtBWDzYE+TdHpmef6RIcWaLcT1YFITfB2rd
wx7SD1dN/cWPK/dNDW1c2b3gEkSGy5f5Zrxt5qwU5qNwFJg70jIpOv00rykNxRtRWENxkbrn5D9o
0HhgvQ3MxmDyF1+lMnuFvhgezF/WLyaUhg+tFG7aLlwF/fqwU3Jb0BtccWBdbje/26KPij0PozaV
AtiVBgXQ/j67tbhdOzNV0JGcetJw470hdoTTA1pH6Sq1GNAIxSaGpEJlv+L8ldU04M49Yw2f2YOI
duAMB2HaaSnZtgbR8ve6+2GTE30QC3sYa5zHC21pE03OPU2UjgvZi0yp7zJzpoRqH3BQfC/Vzsr0
Xt2KGs0qEle6uJtGJaSMfznOfKacmn7arRH/hE0ZE4CoaP1UAGx8xiVmeLbFsdDjxRBaA7nUySAN
tRoKOeM1nzw5Qpf3Tnz2gia9AZJviBK+nupMRwK4QyPISlhsi8nsnSwhraiK2l9lYDagXmn+FnCV
7NrEKFy3GxokiYEJkI4akm+BYQYd4qVaHbAiUq17nq6x4xIG4P2qrgviwG7luT+zn1dUy+W5fBM+
LFp563QQuigdcSWLHKOXHs04tWmn9yf4bvN49yI5TMBb+OZwfpJrrjrWL9oUbMkZ+JcXnoJG3J7G
tqFu65ROJLBB5XtA2oZgSTyVUcn7PPDKPb3DgpTy0X4m1lmIiiEbwPouvcfVZJHB9jVZ+RnLRPzs
yqRArYzLdWnFc6BPePn69ysrR9hHpSOFkqHmViYLtNHTmR2M+iZ/JeczQxQS+eoggHc5M1rvBrU+
YbIqSxCvYhJO1B/jocQeb0ezPcGCp9tKlnaTv8yzgYUNSdng2b38zy2hK/Bakzaey5jwtc/fsnbK
INKh92j5mUWdFoH4V4YycZKOvsw83smMulqZcC9myfIFZOlRqbk38X7C6qyyiaNt/lZV1XIrJoDE
WBAL3mGHr0ez40d39erP+xOh6+xFKr6mQ+IGiKvMMIV3QkfrwjupV2b8wUKqERjpMufMpOPsvdkt
oG9lWdf+3uf0gf2UND0NnGUOGcF9RCm26VDSVFWwQD9qMCHyK40/2tqiVKRcc4rXRle+yboJUKJv
Ap+MnthWsmLa1aVnmbFkYZ89TlGhgOUU3u6y6lV1NcdoXRzBB+fcPUH2+DwDWzyZzF5Z70OlFI1m
jdJjOJeAg6UKp34++IkTHLaJtX0AQBsluMX9Z6DR+iPUCB3/6NyyZQyQmf6LtuyGSMNNf6Qn9ggT
a1Xi1VIEPxS1GGpU9MPkIs0xiS0qPi+PzWmKxGtJx10OET2cauR6gr1wpg/dZQQyof2V74KIruGt
wW2sgSHAkYLHVQWMs94zfUyKJjsV/zaRnANvDc16PNWbBbxgXqKjuiiClO5++yx0DZco6QOAJkIj
+m8b8Up2InbzGoUWr8+40eF9vXFKcFg1259f28xM/SrICK/nIt2QJD6CTNzeojwt1zXCNkB4sOow
ImK/iZdoHWeOF9ziU34YNPYf8ZuLZ2TQIoDPKbLUvGer90P2rNSPiRM1uv0bIg+0PNDEgCsKJ1jA
9djOkP+Ikd5NDSRlBRBTQqqQDlNrmBZnmjecqgo2j70779g3O7vLB1VBLivy3P9f/YiTYPisyI2D
bVY0bxwXlFt/zTGi9KXA3e7JkthENlQer7nd31F7km2oinHgKuvd+MPclqdTVUxa0NWz3zFzasL6
PTgvsz/XQnc5o4H0KdVqxafFTo905c05xVDx0GTJlE5yn1tKrCBEPwI1X7jj5yP82p8rOJqIsdMr
GLyjHqInQxO+HRID3/rouac3ASiwn04qm6oQQ+yr6MBb44FwVDEFJA3xoKfnWZtyUc//rgc0aVgk
ANfbkJnIwG/h2s879yswHGEoavwa7UCRlUlFgCrTJur7L4kFvUtc0Jvfq46tq1qTRY1EddNCtgA2
3a+p8LeEaJoHFvwC2myzCVP3q7CG91/lA2WHrRTlBnPj7RwWboggeo/W2xMvVEZ3SL1zW9ByDYCq
LbjKcCB0NQ0tMNFiDy+8uQ6O/L7e0hQ5MSIYzKcTXn2b9YoaSSOWtnIvZsWtqcbYEkmH3f37Jn8u
8JjPCWwA+fsAAaL5R/RngDhYWRwikJqfB648D3+f63+/EcE1TE7F2QYuWsvVLKOH8Ts6MqA+0fXj
E2B5dyXvzBg5OoBSIHEVu9bA1/xP4ATelSIoWM0l8obsSW8X3VaNQKPpFb4Nmwh7EyeC7eYgCqc3
DvHbsvJz2Soxa83+umdwX3OORHXkmfPR2D5Ej3WTHydcraXHKExfNHTkVY5V7uhAtq5ZJjskpAlA
euEfIJp+XdJeoUtlzHnPALjqKbTjvFK9fDUuTs2fKTlTto8fJlEJynLvP8sYiew8+4Ysm/MC3SG1
4OVboUyJSZVvz14bTp86wTPZcvFpiFp+E1frmLXmZsJWHxNbq+6lbciEEKdHxK3Owl+GQth1i2AA
TAfyMKWGFKIq6hfeVmhh5LGu32N+1/6Y+rjnByVX5boMm1VTSTvFq/UcaI/2sBu2ngroCEwWcB7j
kpAJZw+MHNRY0j6OzYNP3E6UMr7pP1cUm3trEq5njwopXWAWexb6umcEcsG2UlmQQZOAz5qAxxZD
5cD2dTZVgj8Au3WP1xWnTD0zmUEnLOgjz6StTs4KAGxnsmR7lx2nHUtW6HvlqMVbCDK4S8ZCeZir
BxYr3UHB20I2efAcM2WxQqtSlsfS7fwx9pie2HjEh6hjf/ujuWwz652ESlAKtdT9kUwsqq59Hy5u
KNXDuq3vXu9GZRS2NGRhxzoRcKg1nQAn/x6nrgPuVwWMQlWjxCJxj8fo2lawe5el/audz7DtpaBK
OH+vQ+nlAWuFHVnukvL69xcCslpgKAnirMw7fDVMO7FlEkRvA/OCSCHOoAPVH/KvzI9AD9Bkqevg
21xezu4slAYJsqYrPHJEOslA8o18i3aujX0LNlrt0s/5xBcx2Qg+CAmQur+fq3/jc5rI12/F5Tm6
s4wcvp8lP0zNdTLibniYPFoPXYlLPrv0Jt+e2G3eNWgaZov5JWZ8O307l5q9DOwA7sscavwpsPng
CZ0k02TdnP4OxWLSB3Ebgx7d6I3hConXV5rh+4FdFIkvb7/3IMBrDMLBL13MfifOsfYgrv4WdYf5
iDUvTNTDMHlF7UjeOFPRG4p/8jlgOFe614DPTSYRayfvGvL//N+MJHWvD50i541A9VbenofdjY8x
Kjj6auIa3V+Q4E5sn7zgP/PbLa5X2GRWR/WsRXBLu24ZWgUkWaR/k7da15xkb1jEJ8emSh7iPHmc
QdQHFGgFGHWUROAnCrDVD+bCV563rtMOgC8js6Gm/XB6BXWKDZ+D3E7lO3un/LrnMEjuPmZZtNOe
2KbNrMYcK+oPwf3xS/EQoYHR4qO++Sfd9P7+ezIo8hkwuRWzQ4Rns2Y+QnnDABqD33pGsYjEQg0e
+6N8rUscgZUsV8XKZQZu2X7SBuMezbGZ/VwUCrGL4vpuudVjwVqINItOW58zeRXwaljx2jNmTvp1
PrpDCr38PG0kJvQ0+nP7oVmjrRzA4sdOK/bCKxjP02jXWBbKK3TtI+8e5EW+O4TRa35GBoDLXWcm
Oq2JdAkMTwLiUfcZGAZ+GqTbkmOy7WujyH8eHZGej69cELTdbij4zqXrLca/1OlDEySnpIicU1v3
JLYEa++eUTJATutEmdCBR7sNVD402EPl407f6CmN4jZCnvVRPU/+Dtk805eT/eQHxk8gJxWoM0pv
O37PDgE9TMCw2Ra+KB5KXnJFpQdTcHlLnrXtVTrH7BJTFGAK6o4niQTBAZlMtsat93XEH1qtyiBu
8SXmcICSiRL2Vfg0cz61odcnDkXRLPMFzd09SycwJXni/NfLf4w6I/FJ6TvLmb+mGccnv4ImW1hj
UbJmFDiu1OOYtPn/Kkhc4AmbERSDYn0S3tPGCCf7YGHJtyVlzvJvzLkmnpCe2v8UKJ50JReHHLG+
Jn/7WQxr9KTZ+TmicOaMJ7EJ44SzAf8QbWxjzjT+B0Bs9cBlC+T7gCoTM1a9/DVFpLqtY1c1bla0
ql0SXcAAPjv3SKkirVnehXnQStnPi40Z2Y/0Fwl1nPfXNZA2xeqLDLItM8uxqSJQ6k45CmThHMvp
Hjj1LGe9S8DYNQlm8KrSLvzrW79jy3+IkTeRqodWi9rVcw2Ix4UQfPxgjCrmTzGpCCQXUzuaZDT7
/+i/UlaCmIDuIcJRnCQETCMVC+D3ZcSPBKMKWBYazP1/2CGo+pIFcI9m6lCHSmgLKtq1UDrl41Lm
uZzYdqdZqlHb7Teo7PtDcVnXLGgyx3Qhn0FRpFWSx7ReSE4edoAlotjj0CvlfeEQy8IPSzDAzuNQ
0Cuv2RsEXUAHiEDx9JElCuMbNv+hC9CM+mVdAp1FX7buu2KeiQZJvoQhQEiet7ySFtk8YfYPEXMX
QQaqcSU/gCI48gHy/imuEhmSxmAJQRGxyQdf0VPLSIUqQjqANKMPInDY8FFuQEOAeikwkie4NTdc
kD/dLUopBZdKKeyIel1cGdriiTmoHj6bIwO7NhLD7CxXlyTYqs1xNngVByomkRGSfWq7eMr/41s6
QCrwgAZFtZc9kOE/h7ALtyg686ba1ecSJw5rc6sF/KfwrWGrJAzsQFfKl4UIK8NVaqtdLL0mHtIG
Ruzy+zK1YEpYfwAsDRm+dtEkabMBGvOVeUkQuMF+ZxLN4LNCsAtmPCF+tsTLrKm4Do6qgO9jTyuy
LIOQp5rxt7ctoHSl/FIUPgq0YPanJ7zrTfKjtvLrAaS/QMC6fa76vfA656Sz2RmerISPlh+YuVRp
ZohCVJyUMeqB2LrIrEWNHVpWzisyAjH44eKItvB3FwqNCsIzlDSXfaHY+8j2QmiM+j7PniAKLYyB
I8iWBneEEnB7XLYHdVLikdDSR/BuTf/6OWdZYNodQdCEAeFLkOTH2LtyHKNLWW3AniDAHoveT1zT
VdRil1hD5akv0I682VTMxSHuTq+ycSrs+wD12VddxMCpXJ2L0Pc1524Sa2KE22LE1o/RqfYZXobx
KdGeSXEONySQk+oTk/Th2zh4VTTRfw4NlO8/IdCeLt6vVB4Ilaau+7jcf4v1SmndMZZUa8MgWw6g
1/zsEDHnii43cLuRvCQHLnRI8pP4/1Km4L/Clh/oBMI7gcRQ7ZIcYM3Q/+IL02lBpU5Y4NewQJNO
RwF6AyqwwJulFOcW5/ZlA9cVq/lUfCA6Srg0rCaSj91oBNYhKGH3RApPHbWHhc3Aw/hrsg8iA+Zr
A/u+wduv/o8odBV8sl2Fy0O48tgasLoVaXVYo9JKiyzuafNNH2KU31TehmXPNg6Nq6P2Bek65tC9
oaiTOAgDKniUaR1yvQNSuWVF+3g7X1Z0xMz5pRvw9Cvrt75uGrvczXR8zAsn80yZdLRgclHcQa/L
ibroPkGwFTExPuwuxYiBQsQZa6VZr47oeipec8PbQNRro1fGg3miNX16+rOmYce1X8tHRlVyRKb3
W2cp6Z0SkIls9Xp26iWE/VZq3MDkY1hm9KyPgkruXsxnZJGfqs7hXdnHpnAAkkcEUrNjpz2evEXf
tBFxUPyDutIRaUz+vEQ3/eRHe2TmeyMXPK56fSwhJswcPVfq2fvIeFqAZXHEQvlU0v+MAByBoAsC
DA7YaXuYu1DxaFSrIaUuzxSYsph1+oUPWnc/h4RMfZZrcFSK3Fo9KLZrH67kKAgqLsrucAbxfWMP
2Elms2owDhUFbIc9547mkcuz5y3IXGjoi4yPrxJy1LAt95HLah+kka/oVKayRw60xekBh9olPvNM
XewwRXl6HUpVdIZMcYTP7331Tci5dTSWcMP+Id2+VdU81SB5ZV1cM2ZyuR0eK2a6+5KwtTLYq5b7
m/KSt3uKp2GrEeOyLCuCpYgp0TYzx1rphfWQ9DdgEbgCiltUj+N1zmLNA4mVWZitOQ98QwPJ3wZy
Qp/aMlOAe9/aoXq64/f0ZB2p0Tir+8ml+5atyIgXv0wU9GSaVWk+fH+UJfGnrEBfu6sZ998yX8Gi
Jpm8bPAHQSIkmg2nMQaxtyUfcfJAKB/b9KtuXKq/yzsCSP5j+IA0ucv5yB4ZCgDLUFOLGcvOugxx
ZlR7mJWTloVITQ4xBqJYdG7X266r383O/Pq+BszADRRpOzlaFdA7dj5TheNMO0zCcrdPFXThZFuA
litZuYUxdVglQnI3wXw7p2ujOF6onyzHZw2Wa37AV4wPInrG9nHsgjJch6HywL6gPq3s35Rtsy1g
kCJZkKfODW5Rf8/0gjqpQlUG1TE8bH3kphlmWSNbD+/WMQdfT7x+jm8DRkdgBAO3p4jGyxeqrFWw
Wp9n2E/+d0U7zpx9ayLZb+ZrWOb2LNoAiX0zGI3TrF3b9SfVgYfCup28olEI3sV4cEhwRYWOKK5I
E+P5b3Mp8Z/b5UO0G6bgceAoCeKb+tjZqzQUVvLmY25jKuGX4ZsfRidvkaMuEZZzHutgTlqitMiR
i/1V2PDwa5x82JUgNNZJzycrSFjTakWGEyJlAlhdg/cMPYSoA4oo2KlguuadMfm9T3fweQaM57WD
MBhEE43pV1WE5X4cqN71qRlmJFfXl1n+PzV76PdrVg4Wz4lIffxceUQYQ6ou/FYYieweFdKYpM26
9E4fFWd++YgvJlqCNV0C/GkJQqyLG09LPd/UzsiQskrQq9mivuXbKtTcgqhe7lNA7VyvkkrpNLWa
dQse9JKN027PTPB4j9bG8a+kkTszdjrBuhcqhmFH5YyHpZk4IlZhDB/hZe5rA/IX0iNG8WGgby0n
Ni7cT+nLtN6qKCuwN9p44T537WFpGTXhdXk5azekkS03LHhvnfF5XZ77V10ramPbTYCfB/n7baGj
BQl5ccEt0PjI53/PQY0ezSBV3uLF8uiyU78quiY7VimHis+m60lGbwm1mmplqyKWafkR/3y81iYJ
hu81KU7HVH3yqie0UZ8UkOmC0BcW6Jq4fWF9fYX3+e4weJ5f1Kugsr3cOtvZ3Lw6L6PtA4TF/0uG
/on5PXgjQzdMkv5YcwsV17LhEDh/uD/eJKlNRvYxTR3SKqfdLOMDwHcCtqU1BzLg+Wganr05fF9T
vKvB1bIE2I6C3NZHbHng2kVUDqs2wx0sOU7P7FoXqBgGHHpjWQ+aoVsdpdSLAJOsuM15oKW2fCwF
SHNQGnv69m7tgVfLxQF0TJAKEyNoi1QdhsHMa6NBGjcKE4Ulp5JWwo1+FSj0oZE7pzrelcC/NS6T
8BeLWItPjAXHbxztk45hpHOWa5nq5BP3Z/tGZz83h6dqpYypIUgiUlZ7EOkoJxmzab2qDOs4D3vG
0+S1Yhigo4QUE25l09NZ7cqtooP8/ptcXj8JOy+poa46x+QmC7WLGZVOh1JQy8w5vcnS/fMfpg+I
VsFoA6yclxDnV6u2vcJlnkSj5ihJZ737NBTG+tGc5/z7y/XqqJXN+7gOk/5vXXrMOKF6vtuY9p45
r4YVmN+fRAIaMtnz4YJ8+Dvr9Wbo4C0LAWblTomJubqPLJcW0OJ2oSUZQDnopx2OJcF4j7D/qpwl
ReO5heWo2zG6ShT9fbpokf+XUNBrJ3KHVq1kN4eOJU2VKX3U6eNOw67svDTLMyTg/HmMZMC6wMTs
xJW5EnCqWPXw0furHrOmufoJrz+buk09e/421XaIiTE2+2dzd2fPcTWMY5q++qqMFWPOx6DH2GSw
F7vr8UwsnmNsnMVOO/t/aYGTK8U6qYShjq3v16Y6TCVkf1X+vBVsDStg+qP/AqMXmxNW7SfiFznL
r/o0uUUWAZmwiPkek5qqy2sMrfze6dsL3vqi/ND5fe0fd+IeQhRgzlX7pXWYlYq9HF6mnYNa5ozu
QmZobCbhle0MSxrUyclC5UYv7uEZUArjr2erDfc8toD+gabFI/Hy/6tCrof9I2tSSjsp9JL/NRrj
2t/lFdKRdm6o2TlbXuOYD2hHA/HPhPmmd9v7P7ugG/gA1iqVVP1n1APTHKByPKNKqe0uPflOExHz
SYkdrAywUJGCGmplogoxCSLh4kSGDkdljCD1EHiI1vLlFqWI2slUUjPVdznxAKdI0uKFj2DqpFny
SddVrp+iHe5RLHH1aD5UP2aRbG9/hQ0+FpLTvLTmG+GFR2FFhMhrZ68FAXX2XKk9c8ggJmRnOedy
ADvBHqBFAoYlw6uF6YDqTr9ddEIlFebC8Ls3zMWOJoZ7wiiEmZeVEEATGl0+scbb/BjiZeWl+CRN
8wRrRwTdvuwIz8B8r/+D0qhImOB9zMnotcQt/Mqk4Qnx7qrhGZPNLwJePWRdyE8tkqYe5Wq0JX7I
lVXZT9Dou4MrQb6NqLenBIhYu0W5bQ0kHtEvQ2OdM2EXLKwXBEIruTCh7G5HrmJWeVTQyVDegAsj
mmU3vOhi4lX9N5gFCIPfXdV4Zl57KbSHNz8Yzt6/E1yf0Ty7qvh1T5ZGjln803DxGGSmBuZFTKPS
VVJNPEQ/9stuzjAMb/Hq6B8ZrA476GTJvBuRZs00FlUQLRcfsxpTaKzF9NW5rZ1vI67yBF2ygV3s
gPoxTK1d0HQCbAjVcCHoK094wJOj+Sf0zHGaEIHoGUhApYoDjJY1EojVBhAnzeo5DyIftiXJ8GAP
fASCxGixl0GF/9JSPPJwjJOqwqJNqVT1jXzGXfnwqPwvNMmSgBdKqC/xXzN/8F4J59cdbC/DYUDL
Q2SGmAia8JCyFSrH1U+uqzPEU2qMdLGVsy65Zwv9HlHHnI5MUQgbNiq2Apf350bHYebtVZlnZnf1
2cxfapvDF3Kr/CIsP7qebXX12RY15ncTn/68fqh96Qua8DLb0nZIsTiE7WxGLWh0ZXV6qxOoaE4H
hj/duUZKTkO0qxGAUvX67ucbFp5EUZczGL/NGD34qKw0YX4ApqrM733Sd6sgsYW9QyDFW0w2LB+X
CLQEq2eCV4NXLmFYGRMV80sLTbT9PDTTNqKWSwRsqyPOajv/qaysTnGDwGAiAlNxPvWilEVAaPq5
eu+uu+iMLVLmnyTCM6Tvk9be1cCK/6+fBaB0YyVTe5g+zlNd3SXSQmNh+nZMfUhwqsHX2pQVMA+w
le182cHYv4TVhYXTAWPvP/yF0WmMNipvLzHpD9o4DqeUKQc9BG34eEJIv5NDvdCF5w+ojlxA1e73
8eSn2rBmaNc+n0gawYsCfTKm++PZzU4RhCjp9yd/aGFNVbNnkOmg//KJb+UU8aMQvqTkrPZ4g6n5
pd4hMtXmPOcBCfs2o/MZPvy8iAcBXHfhWv0iSKhqGtPyFdbZKq/oAhksijtSBMFIAON1lo8Iovip
QW1LMpS5zRt8TvqybdW33few2y0jSEHjOONV3wchi6SqdpjqkgIWbS+LNaaa5C8RTn2URsa2gCZn
yifSxGW73BBNtYM/ej/R8zGpKKiZHKCkXW9VJpcT/AsOUs7ARS6DkvpAKkAMfURLVI1eGKRMXQwk
uzqooSHwDcI8+LO0nzreI5LitDI9nSCrdGUiB/I/J3OXrJSvwsOu8EqPhK+A1LIUGapoaCcdO/az
4q9yfC+h8ujSA1N7ha69vkvGYK7hKPPFAqwUaxOaCtVmFisRHMwPAgZmUZU8wBgf2/bKD4rB5dov
RyvsUAhRbhtUIvINdMTj74nP0TZSV6eSrXEhcS7uAxwG7/+wbYMt4saHY29EeID9dxM6HHKtLcRg
LZ5QQJ2lWpT4xHZG042/I3hpFZyvfzuXcohdxpCB93hGTIcs9LLNGG9ILGtYkEkCPz0FSzWpQrBB
IDehZYz508i0hDi+b8GQDaudEv/3W0Ln5y1JdK3xab5nKNgEk70BVo63w6QyWuQpHwVRTMP70e9V
IqPUTCJMBQwF1zbOrwQ7PKMqRXyWc8JXZBkhHDRjK8HJk8oYXVMVUQh+BJDdJA/aC2YRuEq+xhnR
6ZEiNG+RKUqTfILgs/g8/K+p6VR0Of/cgeH6lRBKySloceU3o0L23lWqHNKR+EN8++FEjOhyKHjY
AiRlqhlSUC4zYWfHY9dBR3QpHsbIWpfK4CJFzvkLysobHue5cDWdPCQLFP6GSdB04kwQowiX88Ir
f6qZ84Inj5lA6AqWE04MFfXTD3hCfRjBi4mF6JRfGsMeO9TO2wfFCI0bKw0JlsJp+EeMuamF9b+X
ObjEc6xs7aviC+Vimdb3auNK5dPDGRsfk3VvZnJhpy4uPgkQHVKofe+C2qVPZzmlEot4RQZqJRNE
2ymuistcLEh7Wo4bbUCn81bq84tPH6+aDCDVH5VbYYvAC+RRSFo+6ujASOU2pR6lWCzq29MiuHKv
isaoPIbISv37g7JwIZfcYKUin/ZuxiI8DWY+ktsLW2E9jZ8hPk4A6H9pPgwf4Fc/KHn+4cPylpLE
6RmdNW0JrqXPTKDkn5KXA+H4WwOlSK9nO8qiBhc7xwupIvMNk6vcoizDoow21Az1Kik1L6XRJytj
q077Ph3K3R8aGd2vbbzjJEHS1ZVqpSD7KSTLqIsdFzWabIpxGTepFxJC509o3XRRGMs6+JTMqTwO
iKO+m/cUaxK/6bFvo+UAQTFPSR7iM0g4YbfLyy5auReQTq2u2pfHGhz57YvS+L2DIHGiSHVoBwYm
LFjpA4EG+megn6T2LT0MNPcTW0f4yAar9YRdWsg4HRHhDOqgoojlTkxmdgYU+FePLpkFJh3+7P0B
BUtm+nLjsvsp9zrnBxyAEqe7TYiD4X8Fh7ERjU9ASAo/bw9QFnzMS+H0xFkQZ2DhaY21GagqmkFV
CD1B5TaL3LEuKMjDXtGXhBkQ7Oda6h5+4Mau97XJUi5nElvPUsDxfsytMOSr5n8FT/fVFs3ydVk5
ZDcdHkDr8Ybota/NXXcYhyLEBIIU4WvYxnO12aT5n4Txyu45Dl7XjNZa0DMSL0yfg+9ffdkH2W1T
1QJHCXyAYRqXKNCcyy94qpbKaZYDqTNEKeShv+Wui6PqfUQhtV29kUAdS9NEnPol+C6hp4tyeJ83
yNJiGiyuhXBj3iXS6Ge7qlEKX27JTQEvujfzeDH5WbLAZqxY9Jjl2/2CcxEFV+FUxIfd0UHhLSDH
j13PzjGMdmA8duYSiArvJCH85L83yMPQD3/jf4RwKkG67bbvhE/StBrqRCqnH3oCgaoYVAmJz8In
qRP5lFLqok/LBRm6ez+IL37yAecLTRVaWjiqyzoaafRmk0FauTsdRazcjNzQ44hqkWw+IQLXsbUS
zuDhIcT1uYRrsgnG8gZpm5WfXhYXx5dzBEx1MOh3Gc/vqeg8cmrN/0XQkRaBIrMc79sAzXsfkK8f
QpZUuyR64dviFvqZDSEBSP1NvwVBBb1NXbaOd5EolE8f3aFLVjoplZGeXzeQc4cYt6BNuhlywuGA
hhOcDNnm80UvvbwnKVnxBYVcaR65tpX7uhWzx6w8a7g7NeLnF3dK8BgZh5BUvIUixT48zkbjVT59
1i+1GjfIcM9txmPDSXG6QuDiIrC8hO/KKnfkeXiLOtpyaYS4q2CIeF085zULIlm9UVA7eSaDH8P9
/wVtWht9TUhAhYyUSYMqd2pCjNe+WRmUGECcmijdZ4VAXxBEoXpK91IAhFjNlsPrrWetXFUVPC0o
1K3ZOxGJW57bLG02kEssJcbYURCk8vDLmela7ekvFDlG5njTIWDEewy16VivtTIwGrHYMO1pngAC
IT5fulnOWhvnniqqxighH0EmQRY3kZAVojf44Bauokmg02PD0hQ3SLa04xrEuBL+0vtLEHb8xsLO
IrpJmW3IoKNYYT5jOVlwyf+DoZB43fy8onJIJC5CehkBU/HN/ZM5jOrsDmDhdtT9Soi52YBAod4F
9xoDkONPfiVoaEXFCZwOI/1wpjfHyzzcOyXfl1RojZrG0BZqWOsPQ7XePlIn8qlpOA8wXw9jUEvn
JaaafK6mLCMwwFhv8cVeaHIJPUnFJQQZ158TU98HX5M3WO6VunYGKwqwP2o6tx2ukhDrgjz1OG+U
5/pJqfdyYM+INnO15NbZjTJpgc19dH5MoqkWypESnNeg/tQx4TfiY9TX+JzC/Y2st7ZKYCGW6VoU
w0T64hcTa2VOl5URBXnmJEEEcrwEsw8g340CCfdyP9mpOJOaIGyEPgBEY3/UxYBSaKXkrc6WEq47
OWG7Pt3aSPs7G1os+81n+sZsWx9b0d4aQPlaA84mUkM+UCwHI1Lq2mdGfVcZzjTVnDHu8Tb9LqR7
eosIXXp9i31XDHzJun+ClhKY2MIpDfcUlnXm27E2nGj46OfRyjcIhr9d7ct+70NzCPrqW0pgqCBT
3ijUgSa/qyLEny9+rFobIWOILtHo3uGcAvArElqtk0snBTdNL9tYsQE71RoAwi+9BoXcjS1ZCx/5
vmokfT+NKLos27jkrzFK+1qkFhTrbHR09VBJ7Uy/UVoQwQepXUFbwlDk5wk+JFseEjWLzzTESjyM
LJK60H/cp19XH7sdBLernbWlhwVsXwyRdXdS93OnTn815pNIjcQMSPSMzRYXmDATJO7s5zIJBLT+
CNw4xnJDK17faN/yYN2Fv8GaMhq8LLwobffkLGBEyoY6L66bsz+JbXjaptM4nFd/VfUll6PnA9tR
0vmzROB6S9wzuK0VFaQXaTyuKJKwWcusHxIAi3q/+1En9GFFfzlz9MAWnnlAnPG967Zxq06uTbyg
z7voWHpwUyfnWyLeTHBf5BrVBxW1GALaRNJrTGWWwq76SRkdTRrTtwpiQTCEX2PHFpVOR3IK3XKm
GM6Ef3NKRhnKPVuWfecqSehzc7RNNUfoF+PXPNEK7re5ckJvDbO6/0QZaHon3/xPLqlKOU2EIUuL
z/iYzM19WhTq37mB0QOtbrFlxgSizooKM/2WVQgNKzqkm4wbRqf5Y2RZs39+/hlmwcpK0kqlKElQ
MxJPNI5XpFGK/+m989aSaZNT++H3RN3E2c0vAOQKU5bHcQx9aUhvluGgbykBXwg5MrUuHFSAhj0V
wZVxIqahFCsY+Wf+DtlBTfyvznwaQAnwwp2GcZzymPpJvpWsL6/cGtNONiDxNIKUsRdjBKBlkJjQ
dTUJoDAl9csXaCoOGzWtTzzjGwQmkfrrg/lSi2WHKIKSHScQLe9v/nQJ5F0qedFJSoIk19i7sDX+
+VcKkvQX/Nzy5I/w6fvBqX20DgqnSeOJoFq7V03K51L12d5OTN+pMt5hn7r7E2vYbDCZ8fnFgYGw
DBCepLPAiEddLQsvnfYfWDkkEkO1ljP0hA1xXzaXXyrrRklSqEsZEAsIc++UF4io9ASkdvgbmOzJ
a2fUjj5GAYXmIzbROUpfedpQOIdYtAgmq1NnAMxyubjFkMyILrHth5pmcMxPeMSY79pf7z+nzZz0
wWh4Zhqop0XGhzGx25FqYUKIHiKGn4/gvjJvtY2tlGxsVz+hobV3t1mitH9JhAkAdQEGFuMlHMi3
Vjd9sWxC1RqYZ6mPiqkWyAGXQQ+dFGfik6ocsaTORtTRoZN+FvAYXxsIlppW16l27jPuODPUL2jy
a7Sq0v6Vw/DZrMbzkKR9O6Lw4OeGzCwJiZKC/E977GZXcay+9Dq1KwApnUWZFlIdk60HidKghfOi
l+OzgQBVURJ3Z0giqxhyRdV1JAFVIiFSUkl9Q1N3DCgEK+S3FEGUnqPH7wo3LI07xybt09aBJDhr
1WiU5nqjSkFOQe7AfJrios5jMPdLVNTNgIthwo6dzPL8MS5n6nnCD5FdrtQZmyt4uYJ3xnOt1IIa
nbm1lYaijwpBfYmIfYA9l0B6G09tWDRgORwRivcCCUdsEvWeZfAle+LkfevXADCr3txDtKGSReSA
7kl/hLCE7WvGNwbbkrL6RqB0wBNnS355xJ6Hol/zKjSK+U+W/WsD+H0p84pJjP+MbiVqZx3Mv8ku
aZTSg/bw8IqvZI8tyfAuLyM5kw/l08h7VRv9wEdTGHfH+eRyL7idd6505kz9VGRI6Vkmoy0lqzsN
VnD/bCzjJS75BzPt7oLv2jNPG6bl8O3JGakz7oLLZGmjxxYb52Ni4El/KFlehLoAYmfHjL/x+gwi
kAOteswwDVHUayy0JRj72YJO4WDRIImB9o5iCVXTVFiKlr4fW6iUf4lJRUC7xPsz9K+V+2C301fH
BAHXERxlZJBuLAkkm5byuwAVNajov0JgBxLv6c3qWp7R5hIoOdxCEQ9A0sKm7YiAdIl3pCAJiGSi
28v9DA3vxeNXve7N9ofpdH/OXFc0EL0fGDNA8qrxmLgkOLnhTqVqdqys5rnZMHf9bkmdkWfKuW8q
7L5UNNav9QVdzc8UapMRc1AaCtI1fJWRsHd1GBig2CbcBLy1SVQon3crf/JXAQNgvwyUKb9Oa53J
7EfSxDhc/KyNIwVL8pcTIqtFsnLhiclKpV5H+YTSo4/t3e7bYm+mC/AxolmiU/V/JR3ofolkeduR
Bj1CIfBSZXNuxD13VB1lPrcN8lIoV/UNe4VA0yJOLREb6WYU8D4JEIcGvnR9MimVe+yDRMFIptIy
naJgNmg/SRVcf/LDwLTkNh/FizjxRkQoHQTjlGUZ5ezp9ygFOzxVu2p8x/pW+Jhp7uYP8grOMP2G
JZ8ePzW83t9X6tZwQr9NMDdK6dI2BPeeJia6kuZROos477H5a/Lq8Qxunu0NClPYRZRM2qzm1uV0
ZPNNHJ+DFIWY/Ge/9CvTscqEsnJ/6kTiv9HL+Dbbl3KWuXGSoc2eOhMiezZo8hWIrLx/ckW4b7Ix
1BY3Gi+C+EaljfVqqGnrYvSSIcXwlVPNEwzO7XN8WZDuzZZlyzHJKY8/cqhbLFgOzlW+e81XOikJ
iWnF9hld7qHzUBdp802a9mqmU8G8iC9F4MPeZTw5TFKUw7uYoWhM03Ojn4fXSiAbAkmS1CFr/lBG
y5q7b7+Jw8s2CgypaAjuOEbzYLpB0DBeTfZOmX65Sksr396Hu3Cl4TV+7SzWKUFoSKR64t1g08Jc
G5PRMvymz941ayFVHH3DVsLeqT0PboPUwG5+JJWiDd0lTcpRLaydmJVEUxxskQkR1rwB/iV/fUET
Nxs4TK17PV7QyMG3NATszoiPwg3mExzAZnpaET6QBOdljKVVyzefzBwfPux5S0GbDMVuwrVOihkC
nxYjJyijG7c6jfbmGDtCV6XvLcLy2A6gVbuKdjxlpcEOk0unBTa2TSO9cCQWGPU/pq37QdKAoOaU
+I5e/gx3WzwRIHOL4y+D7WzHZruHw7cvspOgdbycUdwZzp4g4ysFq+8gpdfcOK5Ox8IG6sfKXj/t
MpRNbrsihrsYTpXlSwUZvLjTkcL6B0xt9yPkZZy/xk9HfV6TT4yeoNLrGdrjo/ig8YUdvSMOupix
eOP3npTDUrkVblS24Z6f0jpbKxDytLb6ZdbaQlmWNL2EFHQwmGuszhA2fdiIzNAzvCwZQXCPxKLS
GziF7m0xBpSOHB4eSs8kPlyrcJBfC6V5JaAvV46i6SF2/zNGfIPGi8zAJwvvjGKAX06PZCKFS0/1
BIOhhMgdXk/TQbgKSAtG9PsVeP8zomzZhImqN0MPLilozeTk8nGkcYLNrFFm4jM+0BehHd9h4fR/
lsBV9F//X2t1joDztAna7M9uyhiYq5aOwWPJgVgeCea/00e66YRgLWji+YA6iDdFJaMFNcZTJn2z
MejyXfpUfmQnOLPR1BFRnZQAe4ZxKsYltNBuuqT+kUCJcpZ7/ZypJLotiBOU7dCqUUvL7xAmhnjZ
RKFGOluy1YynPGqJenGRszafzstv/FP/M1MT1ziZDK1LNmDOxLyoT37bMhgtz+HldtaZwMJ3u30v
QVR1gFyMEZbtTPy4drp7RQsGVGvsO4Vc8oZDdiZl898t93RLjprSR+kOEU+JIf5HWw9b3pZmGW6C
nnECk+6s/SSwb/ZLhAOqS3B+5wHoNMe4A1qfMxyJOMaVeOPZ+ppzmQ/R+DKpknwhcsetE4q5T71Z
C/+S2/gGoMqDawsLedc8mfKVzeKGVhhJnHdsdha3mBqhDMci9qLvA0gvVvRRrlrtnP3DqZHdgqOo
9J2RhHlJtbEd23wjN+RWyYurTCpNElQHLYBAEKp7qx0qaDGGLtp8j6UNpI5q/wp2+0ZOonjl+e5j
9S1m0tss1BVYuTslvzs39wVve/RRjZdgWcAdn9hmHRKAwtsX7eGafgS7WLfq/1eRDFx4W6vAi1ZV
q0Dfp30ZzHIXc7OSxBqgjP7BFr5DMnZ4PlXjMruWnEsIy6RF9s4N6aiyOoydRYYTMIpUNSFimzIW
E9YQ/Avk+C+h4a8HDMX5j0RiQti0zKWSykPZPPz2x3OC7jGIiL9YPrnydwpSqShsg7BDReb5bheg
QzM+haV7SLXzYEYhjCDqbut1bT+XJyvqV0AxsjEH9cB77mIFwUinY4ofsXaP8llKkvNO04duBgaT
in+Ug0NiuzB39ScnKCKPFpnYaDgQzI0TeGvFMAcgmZZcnYbxEF+X3Rc75f//8YVhwlJvmZezRuO6
TW+GRB4Re2EIUDcYPzi5EOqX2SLCx4WoiBOOYYDCxl3tmu8srPm7KA8RJOF257skxuf1Vxln84iV
jdSK0DUgB0yLvAYUJxlDySVVjprRG/6l6Q9RVJy4IGX2aVCSp+C4miwbi53KcoWXthZklsuIjNpJ
TzT6P0ME31k6iBpsSZmOFgK9Kdgl/GzZSsrzYZZauGweZl14nZrkkaIyX2LMGYFwL/ZiouIDpVj/
qNNm+6cdTsLKSyZlcMcZX4T1X6gJS03lvGDXYuiOG1vyTb5bXMuWzEcupRxxAv7fBwCseXyYjCZP
v0kNNvVqFD+t2bjJEnUOExRFoqJ430ydcEj3ecXivoKHgLpQl0WLXo3vGK6X3Vdl40p90+o5bgvQ
/FShW82j8ese0vDTHC9qcL/uqtcpk/XeV2/uuZ/AykT/+VNIn6D+xDUvimg+pPnhwI+1hH29HRO/
nVrsP9dpcLSNl8Z1lOi7hD7Id+fq241qWWDQg5NQqdGdtjtcupWfFNKsVFsgO/AE1KypeMxgfoBU
9Bh1XK4LIUv25SL2ZyQo5hHmbw0Cy+OBoZ3XBsqtV/d3JV5BgBvZsWDiZW5oRFddWjOaxoK0gYCY
oeCOH+PK6B7lBIhtiT6MsEQQZhrSWws41gxYSRdvQr7jNYm2ccNn1UnUBpeJDiw4dljCKcRlpD/m
37e3BKpcoNp6jWd7s0rEhv9Jbs5nYKZlcdJNqkFg0QOBKXSVI8JAIZPfjMd1hl6oMRaTsh8KCiCg
2KdX/b7cx6E6tKhDwNFYVsql4ZYWrKc1LJWEzEBjM5BxOoFHRktj6BbAbfM8EP/WbBm1m5BocYie
fx7MPRb6c4fQRUp0kbFXzFB4XAglGzXwKs32c3wh0bRkKJECcOpdlrsGBQO0T8EqjAE0sj4AlAD8
BhWEtFHF1a0tqWGuuUK5VY3q7Z+hImdUEha4dDn+XCAd4L3OUyK0GCjP6D8AdunGmD9wcA41ZtB2
+n7qf4mR29bFwvtn18cTB/061kJKBk0gx+4WiPpbYDMOMhgqm3f0TLItuY6bUnDrEvaPFRz+sYhB
/Smqipprhbt/wlMZ1JNNKfwsQRRd986fGis+2Ip5VMIxTeP6y5+m5bvLEYfpX1LNUZNW7s1x3g21
SUvCgKXYWkrB755HAt0cXTlBHXApm+Q9XyH1n8woYx73xzhI5snnB8g0SFERu2tImrFC/p8ZLJuN
gA/Shs8Y0t8Kaa+UG7Nw+S7xHHoLZNXIY8kc7vI+9m/gp1FS7iw8R2Tuv23J6YzPZa/KNL6nFlpw
xaY9UoAqLw7GKJImlioqENoN02How6wfYkfZ24wzfzMUfHyWOZDsVA1FeGa5A95/TrcxxfTip8p7
jKJVWIU1vVqt7XWIg+2+1pYToRbZq9en6dbAa9Lf2vMmWBuUMeIRIEiKkYcjRgw0qTmj2UfIll+X
lF5i5OeHvtx6MXEXiXDFrLc9FcJEtr9jRStw7+01SZvttxXmCnWrjRbu8/z+Aa71G1Xb6/fPxT4X
MoFGaKbN+iUrdk3UpCKYSqKkeDj89mJrQf+aEvkxn3MvS3MQAgVreIKDkrRARUCBOImN+C5fqhS/
qLlX8QHoRi0R8sVV4iT5lAD2VA9uK0T2WlPwJ6Xvy2GBBdUkOy7D03Z4WxLS6Y4ndoxfbQ+sq4Fj
Cac1mqXYAj8oEtgyh6Jst31u/Hyin+7CXVb3G681q4m/nU7rOU5j2Rzwp5crV/ZmrCD81VvuPYf4
8sWUpb4iNlapChAMHUX8f96zActBmnTixvY1X46Vp+gnxDfnuWnI+srQaQ3XQyLiZGT2uXCDtsQM
klnh9eJJoP5wxkUYJxJgJAnzxZuj9Atb+6jNv2x6CfnnzMeoCMZjLmWFsebwN290XO5j+NKrtv+v
S2+miukhxVU2N1uYOFzf0h/We91V4Ph6I9CdcIHNPsV9VM6vpt12ogRVIjZiE8DbUJSe7EzVcLBq
cUhl3o52IztNHyYxf8wKHUOYqSQVqu4VYyXz9zL8qXA6j2LF7B2CckbcH//QYd1AYfK+8oXbbkWp
6a1VOHBFWmX832Aa3Vo0ZFSTrR/bKgi1favdNxgmcx4YozkdfJ1abWH/7KofDItlqGOt5f8RKuYp
/2CXHqKIzdHwcwUAFAmjIj5dIZ3pxT+aIGyDrz3YlT+9wfBxn3L81jRiyGzwWcQrEwRTHgwii7we
3gVhGOQuHUU+DhqtAF/okpG2vncTEQC6AXilv9wwYJz10d6PoOh1ISnkv4d6yDNvpEHlvpXprWod
n9zyNmInrRyjPmEnvscBj65LQeEjvstUb4BtIX018HLmjL1SgRJC/42MsywYmlQepPio3FjLb0gA
KZqLD01pVB9bGORP8YIrOh2qHIzWcZfrDtk2E6p99OUI9pkjI11/WbvP7EYTZ7A2VcTdHDVjoj+X
NUu0pIn66e9gXJ5ut8Dc0d76z2abxd51Ce8QDQYcTCpfnivdC+NdT+/e3LBVe9+UOcKRGp8WmMOz
lQ6XrCtMmIhyJTUc4k4c1h4YyAfPhod+bMleOVowBSfueOj2T/dAZxEIQRxTYe9j8yjP5A2sa4LS
pS/KSmYr79md55YM3ndh3hJ66DKVazSlrm3d0c33oUpHaxShXoKRVtsLxuf3HxVWyePGB8uJ8Br0
sSuLOzeMMBohU5aav0Yvb3EBjW9e9GHHjIZ2QNl3OpDaQy3l8+b+NDqhQjr7HKC+vXAJ5CfXWkMI
Qz7dNb7br2n/e/1IgJYkVDG1ollt8wB63GX7uGhirRJfKmNLo6td3miXPa/lxNCOAUNnvuFLf45T
WLG1hHUkUY2p+VvtUPUY7LavfUw9NzuZOeowtiJhhPek3UUekKQZLFLVNnuzFWRCxTFcXEexOUkH
/+7lGmlJOrZbnDZH8U3iqblHU+XneoLGNCm9EuHKrIqIlTProY60ck0Iu1mGJ/BFqpIBxMWg5WVY
wrS16L3Ws3TvkYk0RKOvMJPj9eLCiEKmpwDzP2kS6VIrJyfuajIrTQWII+Fvt50Cox7WYjFrd4Cj
oBlEkwGcU0Q2KKJ3rxdwd1+ZUIEDrs7cgD4TeevzeW8l2432a7+ewWNrnRVkqkjdhtnywrW3xVYY
D+Xk0tJawmJDBYOwgW2RZSTQAgpYJaMD5TGVwyDC7TO9wYTrNWh2yg0ApKwL9NzuvSsuEbALgmGf
temXp5sjK1+9IaI4LJKGq6aLVMNRboO8LiV93T8bPYzgJi18iPufYXOX6IlDJwgIqNgWRicjs6xN
QJbbVD9PBweBNN7QN0Uk8+yUDicX5E4bsLzWMbW22yWdOh+cJUvBZULiqXDZATYV1+Ig3T71vezf
IIcA6aH1KbtnxUsmMmmkmti9mMuABtNpYb+eYUFBbmBUJcjikwoCalCYmGa3TT3C9crMomCM3zFT
Gm5qVe1fjlUL24Z89zZ4sJLrGpTAaZNiHwwujAx61+vhVJUT7TOcP/BYyaEswpv5rWis0szbSz5x
v1YIzTWnGgiUb2Tza9fLLxCEWTzBVzwkhtkTm9u2bTtGWKILr3Xqnciw/ZGPZm1KtGG73vNiLDiB
dpelvdvHtQvk3fb15pDsRoOmJwANaDddeDSYf4VMkVUSjoDfMzXGXdC1wpTXKcDZ21HJBXNBMSyo
3fOZt/npiYcXq2Cc7XpkKUBj4oLJkLmMzN5LNjgQyz1CXtrK5mw8xr1WqID3Q4L0WNvlZaE+M0Br
gfO3An22aiW9f40YotUxIZe38/ds+M8/jqwUxjikaBlzh2+EmoYP3H+pijutpx8SR1fGz7cYiR1m
prGX9yzytKyQ6k7oejwiqTyUZx3T3r8s0ycto+Nv0yNZ6jDytwbNN4111OGvJT+o3BN3Ns00N/XO
BsAOIFSrNCSxqotNSfn+CwxvaAPRWk0ahhzGOLBFWy0S6v56B2qnzavUpYfa2Z8FqVgdSoOuyvS4
S5UMLjMjrxMeI9jSnVqYo0ZgaOuChCVHrMWYW+InZWU8xC6yk+nj3eoM2EyzebBHj9SuyIRDUGAT
BWasn61hQZcq9FQZekMehXBtw0gCnVhRaN2JEoVWkdTbwK46Cmus4qG+Q1n7A9NABUHITvuZKaIT
lcrClui87zsdZZYrEGQoPuHuaQTYjTbJOCR1CjOYWjJTez6oxTwTCn1ginnlE94jxdjsFxCdbi1e
CATBSdXyAkui1fEegv6rLDon5eZjsxpUZIDel8MmqBU03f++EBz9TXrDl4kY8Aan66CXq2SyVXak
a0b1WwhpCL2pQhxU/DMxqUPDRiR1lqEmz9S3RROOsy5V+lbtUS53njJrM9f511ceZoK/skXzOKWH
Dw3gDSToEa1TQrmXPdQMj6dHER14kMKz7w/X49glLLtNzwSYNgeLD5rwJ8PDCQEUvfUj7Ikm9Uhp
nEOcbkk7XPcKW4jJeXLFWw6Cln2OAsVtXR4Owg7G8wrY6UbAlzAVqkLzMIa+OU/4dbhkgWspkEiQ
2xK9JScahb6XeHcvGbNuB+mF8IQw0x+oB1Co4SJe9+zfzfeg5E0uhnawPEpArxoBoOFqhDePjk2d
NY1+lbdY3T+yO837dJOpAFc+ihpclDH8ivKOANDlzYupYPgIX3hgTB6QpJhfnMc0um/HmvN+Z45H
+b5UDlsLwrKNycL2GFStfhJXoktwZWHU5zlqgSDpwc/UJ/bWlapLLZc0/31UK7It+gIVNRxgazlt
EVzeuEX3D6INmeETBXe6ev0spTBXiH5Ul2z8sN99XG5NoWBP2k4GkrF3jGbeL/S1pt6j1RzoG7AH
Yy/xM5/yzqvbteW/hyJJYYuMwOudG6XRNOTJieJn6qObOr98lIrdInSNvnLwTtftqJRs1AoGGgzk
IQh8dTQ1TAOuN0jKi4G4Dszpl63aN1TY7nZbonzMnyhl9O1SlqsG0NTXNZ5ylt67yzI3dyhi2fKc
OTqAGezse9kVeKoQ51d9vqKVOMHu4A1Oxa+jp5t6u+1sAGVFYsiKopE7G+dpMQ4EbuIlmuCofpKA
9sOnmaFr4IcF75ooCtp+sVitTQ/yi1liu+8Ohvcs95PkGztybHX+2GmteEb+hq3T5o0DgzabC0J5
RsCMSckSggyen/uamHcbXoP6OkKJxuWW0oD+8BiVuqgDt0OMtSEEhsXOHzwWOmxGNAASJY/4LB/I
wYLhIuIxym/OdBHCN0DJd7sTI0A9eQM4aMCscgkCL8caNqblhvPA1+Ul6ZAGTkSwQygVnejCyHj/
TlwT0p3QbhAvIjjPePDys2jHS6nXShVto6o1/Ra285/ZSsRXKxmXLiugTmBs/1ckfG5hz2/Tw5DD
9CMUTPZ65XYcry96G/vQFPIBGauj4f8161DmamBucTG6W58/BXTjDXFQkyjJavVVqMo0CVjvzK8Z
90qqLLzlqI46U4WUGHuVt8uwZuuleF+vxKg2RBpUPxQQl0GPiC9xQq5xEoZKg2YWXa8PY9bkum+8
o3XDIADJ6WToOFlFMxftr8rL9+PbiZeYnoCEFu1UhgiG6AYz2aR5iGzU4odkEM/ME+xYGJQdbgZv
zrIelcJ68V9upRdbWXkK60GKtwH2y/o7D1XWLMfJne971TFsddNRZS6tuymgtgljEXgkqeuuMNAx
7xTi4lXVan6I3j/cm2PKtJmj/XLzAwyoWglngt89YgFeyacaCqI5FC7XykesogKVknxIRJ2LWoVJ
D7JXK8J26zyDPsYKwBAopX3kJRBFfPOrPM+MwbTwWcoY3N3IJgZfsBOaI+fsQl3BCa09VxtLROCA
ShwNkzedooKaov7tbBVv2caFRemi49uPYmVhCiiwy4qiH5mqIAugx+mvgZid9c/fHd9p2aUKhnez
LWpU07w8Ljs+FeGX9YFFZUVREDa/G8Spnvmtihy1J2X2Du/DvsxC4lavIUH5dPt/1ZnbKPxUWW4n
a9l47zC5YpD6B47V1xvFdFX0Dmr3JO5gifDx/IvKnUAuugZmwQYHP+PH2EtrVv2j6zlHo3p/TgIY
6jZWVy/2ma9677TLA8Nu7R9OKofqf+xAxQTX3imQFqvkBzBZb0GdE0yUxEuwrEQomFLhAj54CvM4
f1q/MhvL9gkjBDX6X9SNrIFO/16+0+UMsq6RViSF7e+egkiDmmnFVpA4/iXP0qLiTGOz8+oYqg8v
Yt8o34f+455359XTa2gA/5Zr/811KpeJG+uoPqBcJ6MgfzBygvPhWve1Aq6xY2R1sMi9KMWWP7ix
CQrUWoIf92Ukx8dK4bqgkvjNhdVsAkYyLZ+u55pdcUaamSi2ByhE+5Eg2E8Uurm2eMIc+ZSvLau+
8U1De5VHu9IxYpd5YvYnP6FxhmSJMxMaLQfPnaxYBqbpZ6/tJw5ump7dvvzSPYvRKIRk1vzj8OW8
7OptEuq/3/eJd/NC90Bd8OSj+YTioxoALDv2zHY1b3KfOVfGZawukThlfoQNnjmf5VujoOEShhOI
NSc6eMGjW3U7J7cVW03MM0Cu9+VdG/KTUsN40ubi1FtRSXAenEYB+/i9Br/pbOXygWq14n5mI5F4
KZrSN+KNt9Dt4z1da78xt/IRKdjX9n8onIYxtGH1JIAZmxFuK3ZATZATGXW6bDM2uBvWHup6Evzo
QsavQ+N38Ba+S7PIhsLLpET9v1dbmcBr27d9lwkBFXjOy6lcFtoEAkO9fTCawQodnkz9R3LaQWkV
KfRFSEJh7jL+CZNxQ9m/tGHFcH/wYpa/4AO9ytVcngeRGx05NcIY+QJVB1ilZqZuhM+UNDiv9CCx
sq85NGLii2SWGHL3aMTnfo5vGYa35MUr0a0raL4cbVQYUmDgDS67Mlob7GDr8lBK32EgdS+00ct1
6sAD3yrWj0ltC/xAq27vQc3EzI+R46i32Bjc1S183EAp5eRxd2pBNc8QSTuW1wFq7CEFDDhSMBtF
AK/ARRQlIMEKqkWmUKt/Q/m4I+wxADmSEjm/CSTFdvAHBizOM09juGSm9khgud7mrYJP71qrAEPX
BEVazCB8b+RHZiIXiFaXzV+s5xkPO4eEXszrCCc8MEmiFJAha46S2EWK3+hfnrzwU63I7alTb76p
ju9rQDtdZsB9YIu9K0Skl5lHtFwkC+uxZpMthd1e04HVeFWAeVARQZUNNOWH4LV3SGjlyc6+vzTv
NyWtjJX15dilh118HWHKvS7AWumR3Vvh+qQB5xkHRxIi/nt6QMLtqmNvE/CPjdN0M+wHvQH+YgsK
7lX/nOsMzf4dZXKPxRulrRQhD2IbtQM75PPr3DkfEtFh7I1iTEtU4AiBec4U0VElac1jTJEzGFFk
gByRwPXa3qaciR9uXAGVZS36PdC/jb+tIhdC7MURvr7tiTcxCH8NxZLHa5pMbDadDTT+E9nfdF3P
Szmrwm+eawEU29Cwe9A452Wx8r6NBM6zvWhlvvVYligmo7pLIoKypjR2RHznJASIcd+IPOMXBjdi
JD6DsyDF7RaY4BzRITMUe+Iqxa+xyE3pYI01X1p+++ZOzxDXN6uhjld6+j6C1FJw7NCLx4twjJOZ
8MQTq2I6hmLzvwA9vFVp+jneZUhuBzm6wDqblzJo7TgvHqz2NoHXy17VtvYtKHbdYGV1Et50MKpQ
FdA1lAFwgakAMmWbIlx2/v5d/TKpGnRCRsikPcP7jibIpdr2vQKeT32lkI/lM6eXjkOnhEgA896c
7ExYT6h0JnCjwLHjTNHL6NhdsvTq61LD2TkOKFuLrL03axaa3YXOVXFjPZQ/l4SC03UXh5oWpIlS
G9OTAJgMHPRA5i4f7sgFyjSr5oBbR4hU8L6sIvdljO8AuoKAw+Bg8EKQamL/IM5qccu/q0GJ8bNY
m6ezzT6QJLRcne5xaOjOEOwhLkA6IdICAjvwYbX3QZV86nxYYOl+vIV+Fz6J/ESxxJtaywsHsOrk
YWgP3CrBXBHE0ILtqwg1sGyDiZFIwiPwZdMndyyb16GwlSaAPvNxdklW9hNhVar/NktZ/UZOqfSr
9ryENRinjHTEwJehYTxyuK61ZcfZNTRX1/Ww0U/HLGr4DhWnnabpSDaX2yLzWvNsfjrmDUtQ2GiR
1hqKsMjkk+vhuchPJOP/o7d//u873Vt9C038BHyfMSDVUjZijy2NRDbXIBa3Bdg39yXzC8DzAdpP
qct+GUMlP9HedXCttb+a2+WniEqNMe/QGo7E4yW59BGFyn0+p2luNPeIajMQ4jLpbmRtSSf4QeXG
Q982aGkr1s2vB8p/X7HK/fAqzWxHhQhaGqbV1w/4zkHJiVJiybS1HpI5CsFD9PhR9UCjDDvjMPDl
ujvJA50SpHSXaMZJMx1ilUXiWkh6RWP0tjJWvhCfnk3gOGkxJQRQtzqtsSVrqblQ0Vj6QrZNeGMR
j38kpx5eOddLewWDhtzaf5M+4+6wftI6Lc6sKddDHoPKnFgaztiP/s+ZSiecYJsJtLDVR7lmaO0W
LkaToVtMYS6UMm6IOBBGEtC5Q7ub2ylYWTo0a9w9zta4YfGoaO4BwjyBTX+RTwOn9K9sKBi7tqZq
chb0zTxvToiFnJScR5/wlhdh/COeG6dyIQ551fjLNHScsolE3FmejqB1nYZhwLR9n4FUUnkI10Nc
2OTui0oF6Vyd6rHWvRTeDSOGE7BEQVE4hPAtlNeC7xdsuhdRUndbPMKU7Kl/psZQTrBR6YSU6rgH
f7L7sqfjOk6AfimRg9Z5fx9XDSMPY3umEzZUc1VQdTqWZtLzB5Y7Gb2xzvHFdcSKd7D9aC9VQMRX
Qzvp6m8iW/KvERm2GnvmTnVMAv+Ds3dQ3PxAcqzNGlV32BmVRRHPO9m4lfeNsdOtcbbvxQ0Rg3zN
AL9xyVBsQzit+jQe1Ikrw7js8mg+ivZefC/1UG1Yit1KURgi7dTfB/lVdXtKiyZL/CFGDJiRIrOA
gjRIoDT4HmTKsZ3Ma1ni44PVPV78zfLlryV3f77jwXhBgSklduv1o6Sr4E2ZhUYkQuGi5TygbP8R
oH5Z8kN7pAtJZ6kemHK2W96UALgMrC29p8r0YvEcEnDLi8kgUQkfGXKNsG3MM2W3C8MdajMwHQK+
mjWQEsS7iVfq3+dXV7C3Adt0N9AqZlRPHO/pA3QMm4epmC8X+2Hfay8L8aHz62KfBDHcvqv1n2Qs
ZJGb/FTs6RJpnek1pZw43d3fWKpuW0eqmIfja5CN5BYdvZwxdhSFdizuzI5/OngQ0Ym0Ayhf9TAy
AD2APT7JSeC6YcFimE2ibKjKqswcV+XTY4jm62NUbc8yIpeFPdCrpdzwCliG+0cmvW/u10omB11h
LS9Hbwg09bUeSzkoQZZOuXEk/ZIUG2yofRZV7ir79C7G1h7HtE4fAWBNVxEwA3sfVnm60Vwy80WT
XK53VtO1wNxii9by0fqx0fSYFFfY4GLpprirpAaf58NKxnCcr1EuVoZ1/kdlqrRbW/fNBXddTdtf
cRvNuWdVuyC7Xmsgc+B/cu5v56BhjRdKYaQlJ3T5gBDvzP9GbsSEsT+xKI/vbfkAR9gg6oJnx/kR
0ybvZ2DZuhFV7sx+8vJ8XfwuOR5X4DdAjFu+W5vANGac7IYYxO8IW/LDsmOECSR84JQs08l5Q2PS
DutZwGGXqvRs8Hs2I4GT/s5g4PN4+W0vLlXGGnSjEgyL8Mp+YBDsc41P3QNvjS0hJENexlyofugE
+8Xafr8u8CxLq3R35OOZeaGeOMJlVy7m9tou+5+eyPMEfRKPQn7J7W53BEdLuaF9w2Iw+HxsZ9Nd
L1sxM7oWAOcM2fl7UfHt9hAHJL41ouC70IWkkByQNHmNzFedGqLK+vGoTzTa5gd533M5ti3HLRVI
X+VDvVSsbvFIRMqn/1r8U0kypwUeDnollMBhEMQgGersRPrZDzrKm2HLPDoLJE9xWh0nQhX+7bfN
XY+vrflyNsBGWMmW/IUqO1ngSlC3KsUJwsd2jXNmLOT3gqhICWnpnTJFEIr/d4CMim0hgwlctLWe
mQ7Bj8AOQatO1FIyJrUt4j6lPrc8N9ei/IKfBimPfA2H09SK/y4JycImgUKqewPVTpdekqPJzQbU
6vaTBYyLOBkHupytvhC3QEC4HuUbYGDR8m7UlRjo9hh1XtB8hf+Vg6FDAdZChbHCDhjMdaxZOgaN
y9/GxLK1JLftziWVRAau3jtWs6vA4qmNZUIg3HtgEtfbV65x4aG9/FtMBLH/kQlcJtbB6SEi37mQ
g3NzDXdr3Saaafmn5CA0dxLoYxJsj4bwqpVol3arsiDRN4JG9VYvx6zObkXPNdt+BLIPLypWddRU
EJVhBB3umdxjTwEM1D28R8nTi2d3x/nWnzywbzovh0tgo1/3Y51FgECa73kKaaQZh3twc2SKZXoH
L/ff1dU8jZRWAcbwqhvAO8Bzh0KfjXnTu/JFGGb8PK1FOHuDkc1Ma9vdXRbs/Iyvy2NwG9AFaXuA
li2ubfCZvVauiB08X8kBeajRH2fSYaIkdK6aKkuXEWBWV+jBxqMgazBGcn14MWiWxaUlp5mb9o7H
gN/Vn9GhMJvXOxhFQcvBKv6FfnJvzgtfYuRN6dBtxi15tidaJUsYxbrkKSbzhK1efSXv8tTbtFpQ
u2OF7h7OTm8utkkZAhjDmL00l7RQYXozLo9n+HAXWo3RS2Azq/O2uTuAFqT1SWRvJWhbiy9aiHlp
mJUREb7x2ysIa2MTS/iOT6QjS8Kv/YN8P11bO/UJSLj4DrnGr/6IMFzrUSL44PHmaG20vKfPfS3X
z4IHhkNfqQAGTsnCZRXluJpaantkfzCE3Ij0sJDksHjoV0wIB8DWobsP7IlcjK1M/63kAU75bbcq
lQg8AKmofCPIYM9oQTGL8pLeu5cw/V9PKF0TYR/YklE2/tQp6ly2gla2vvhsKvdlqah/Kf0TFHbP
FY5VBX3dW5sSTpXNNljcXPFP07YJWu2aijezaJOka5UU3dCn290rDXWSc3AqYsTw7DPFjwRyHdH6
DAxx99U1LCs224ktaUr4YGsiYNKBamKIXDhPMB7KIn9SmBEDs6EVi9wiyOIBMZuPWIUS0cda5FDc
br0Y8DTIIM2iUihnliC9f4nIKgzJxlTjRnGixMTqBydqaKcoqaGZJlNssZF6cxtr7cfKUfTHZqXZ
lYhfKolcOwaSN+OljY7VERZX7/k7UD4C/at3wkvf7TdpQUvw2MTVhAD+FlI/D79vLyw+8pxblQv8
hhB3Smx7dl4mHEbZ+UBtCZhz6b1+5+GBtN1SxpuxmUGDjbagUAMyPpwenr8jwK8ne/Q98F4VH7i6
6UaCasqZey52w3zCP15jfqvaMG/UzPQiPAfp1W+9YjvnDAo5RA1tN36VXumzd+CnYRE4MGOWigpH
cwfhcIMIyMpCt4mxhJyuEeKDpFnP411UvAaBx2dBrFEDRnbkBxbVns1xMdx2n+XjDrITEZsotrFH
fQeAJM1h6KOWM3mELA5rW6a97jhwy24sgBjdPV18IUkYTMJv/0TmiZ3JptVkRzTRwqOo75HQplEj
rIIY0um3o2w9FfWmUerTb7n0+6Hx17mEhzCuw+7rxsYcdlEefWUoB4HbWBCGl5ZNVhJLYA4bCCDG
aqm76waqb3IaO/wH2HLQlmjnl+ltJqj4rMx9ptquQg3McsSOeA3BiYGlxet0nCChXNbaiHdcaD0x
dQrSFF+iJooPDH1fTVVKT1vcxYzNVIS8yD30NecuIDmzd8VhhD9sInahIDZhpqzxaeu2zSfyMJ8d
xXxOLgGTNXSCpfk1NgMv79h0oVB0pGGjS4WBiJcKTcCvXEIuzQoOEHBh62YPQbN4arOire/zZiRY
JkTuPcKdVweaBrlbNSIwqwqwwL6Urtqtqf59uVRNGyNN9wrcSwy3jYtNVeMdE71Y15wzmL0fLyv6
vY7Tp6l8xwCpojiZCvcgIFQwjZwogSBzqKL2D+FSdfEtWM3RQ/J1DphcYPvmYGUQVXIKf4SZzDIH
tLFqRhefhjfwFrIIGvSDoehMw5i7KlP5d0TYdA9wnTdHACrbeStIZ+AoUet9h0dagOFZKshs4Kqv
/69743bwZurqhZCC69AIG4KBuetUGgw73Az34FojKbwxoygusjG9CoRakWu3XskC5NKQov2dfB3w
xNotxR7a9ZUvPewtY6CLzUGLVcgq8KLuTZvYaFcKViM/MRM4JD7kGOy8wptrIukiq/cDVGX5Qjdh
B0XvZAlhPDwmrvWFl09NFPn9Lqtiwkd7yztfdHLkdvxw0vW0E1TdzN3aQHgmXQ/oUdq+f6UYTWbI
S82N1GHQjhCU6mP27ZQPE5NncWTDVx1PP4KnRozINRNS3QdwfpK4DVCto4qioqKCNJJiRQ01hVkz
K6TkKy5LkzJi0MhzgEcLvErZGtDvVR7Ofvqg9lKpkRjdkaibKhvdMBbWRkYsSe+KvyeaPAwfcl8j
zMZspZq38lk0n8nnAE41yKlTLm01IR0l5E3PE8hNmLdkMr6pNmrnzud8HzR7Ckzc44iNix+xYcGp
Gejx++bv+qmycj9TWCRRbK4bVoxHOjipGfbAerV0sMwBKizoAw5Lyptu1SDg2KB5mIcT15sOIJ2N
QZu1NUFfKkSYrgV3H0BOhpL1YMK6pVRThFdkxUCld36dwj+ZpJxpCmLDsvRrji8h7wty+KvZUxFz
7RR4qcWFwcfM25nM4El3t8U8xTOHgsXc9eaSqFeQUyKTY1EiodXiYxC4d0vySVHdPJvL5I40lzim
mn1qV06xDKvCvWrOheneEejh+wHBvKLaG3rjztAYqGxXZL53UKmCEZw4pgUXHVzG4UXiQYKkCek7
QyoSo4j9bcyK+geZUsmJgjUrEan+xUZkIei3ixmM3WI1NCL9ZIwABmRAao/Z/ZTV7fQI8vcRIY72
UBUC7TkXz6b2noYjk14LrCvx9MbfYeQeLWs1VoCgNR228NQIAMeHvORws1mEWolHCAHxHsvnnnSo
lC5tFBmhWKRlqHxbP/dXKErca7JXOa200uCPvNyiUfItnZ2HEYsxH5shuu3oN1osRkHTHsweeIbt
6M8k3/o8+vXua624nX0kS3tnpdqKh5BGSF99BaxuY+60QLC0MSNA2sgrAivf/2X1+MFtqA9xtJhE
/A1SSJw7bWXEYZorIzKIcpAARweKDlYDdX7NXc/kaSrAp6qaWEpL1EhC40ohRYMPOS5DS2ASjzMI
/q9gN5YOpRQZ4ulrUVXcllkwGJF/hNByhzlbG3NMeQfLkxPuzd8VNI2vlvfbJGe+/Jr94Eb4mVj2
0ueG+L7hd3nUOJ36P7I9Jm2+v/YJCEcf8P4TpROClYLtU/WhD6KZKkCL8hbG2GV2ojuPJvQUI+wP
QK1qh6CxrY0/xk6F6YtYwQr5I3UQ6zZ9B2VEGYXjkABD+EFZL1/5kgMF8sppxzbUrzIaJKa6Ed5M
Mpv7eh9kSdYwwrcAdBLlcR0EqPLR55cuCK8aeXfGEozBQ2pPQMAj3s0zEpClI0DoKhZHh9rsFe9D
OPYjXZg1KASP4aN1kbCFJMZu8c8Mqa7Ot2zfq6vZHjgDMESKP/W9H2GU/hl6bbFsHL3m53EUUQ22
+IEbcbw4gPfdckRSNThhcUWXgFPwFgj9vFXewol9IfPSH4tCxF7StLiRmNCOHw0S4BJKA1RgnZSt
JT0VYhlO2lMY9snUZ75b1UZlX4Z4g3YxkUR5xU/auOKQqhk+CcUlCjl5HtfQu7GAPme8Kz93Uk/g
rRbmI0i3vyFDHa2hCW/F+kneS2xa8AAorwAHCuSe1n/48ew1bclp/r3Gp783bWFrO2lWUS0Sf2cw
dOI2GX3i0ypVS9FG+mYqIHduqm2Znff/doM5+ZOfap3HXF5l6BJMI4sS0Brm2wUsYlrjIUP5494/
GxsS17vTRvAlS9S7Bv7m3bkwAJbblarrtrZaURZku3Dbl/8wVOAFgSk/GYi7CgTa/asvAqi35Cmf
+WRruN6vUsCy/lGBI1RfegpL1x5f9o/UrBhVg12iHqTAP1GhkNc3Y5p7Z9xcIiemYRAQtpgjVfQs
9J5DoloIPV3tOM/MC9wjOK0cpV7P7xHD1KMC1gVndtUZs55hL0SdLaU5nk1tSsbmYqv4YQdi/ARp
A/Lcgezlyl6wiz3iZ+AxMTYoerMKnd5KwGPHLfEtU2slf/tPdIf3BB2zjvpNYcaXFL9m24sYhz/b
9OJwSIAo0M1W3qbvORcEfa3acs21LLS8ToEp0ZpZ31wBsDKAOKscZtifn9ug2qOLD9zWbZW0JyTh
khfZeR1gW1Emo52/RDvoz4vbxZ/1X9oB6D/0GNuAzRdwIsrzB/R/0g9eZ/m9oMtdErimh9+3XwPo
2u4luVISEiCvyNA8kVlUiUn5PrYb+tPd8ng9zqF3DotDs3HXogeFkw57eSPGj+NUWT0/QO413W4x
XK2CqXj9C4wz3ukKwJhSCzZYQFUlU6icERysFuZBnsRvW6lQLbABriA2/VsJ3hTCXgW3hLYB0LrW
C2r7XWWm4skUpBbkG1isgIryVvsVtGKYt64IEMhww+6SBCjAtwdYTkBBk5nc7J0y9dradJ2VNObq
5oY72/KAcELQG42e4PQmsq5hQmbxc2AjkF1KzMDXbihPd2RnoztDtUyxGztHUk+yicirQoISfpTY
BS5F7GH2LszSx5y4Lk5Qvd7ztxr7Ozhr+up5Xq8sMH1hZuR8tqHDb5y3wlw2E1qTipKYOdD9wNhr
wHUI7cnCWPVt126WxpeiuPVWHD8/sz+hM56lRfkiy6DZDEJrl7o2pYuG+O687GcXPPJCcnOPrMyI
NefRrlgM+PwGJ++cZqn7jKJBm1q8vigFENAudRdk+I7qvC+iipcucp0EfHOWAVAhkn4CSgxFx0b8
c6oUKci6tZPGMJGCPTb5NcoM0lDD7S+747RsXvUJDK+1CkMGdsRjJ7qlCKYVzHz9SzvQaerd+yzi
1R1h9CZoZby1xpgTuZJOBnZmJpaSGn9Nn77AUB12e3hCqV0vuVSuSSiyI8nS5uCWdUtZnDyh7QOJ
2gRTGgf5Wt0Xcwu7I+xu096a8X+BXDkkIB+MkZO+TRgkbsTYQ1WnQE0OfYGr5VgdnzuVKXCqfplU
FCIgTt99T1e4rOAFa0eOWmEEre/ZtcjzfUDa3Tdc/BmSd5TYrqukmcpKrX2gDjaAQfLSyC+Dkapb
AsS16rqwfl82Cvar5mWxTu3BeGaUbXlwSJ13s2jn8e+nLewokusIhJzHVMBVv1M0qP13h3JkRvZp
BUBKLz+Rqh+TMk6KOqP8oM8IXbiIxFB99GogUJ0n6ep5L0/Aw4W7fwzTOviDsGU3vvFvaccn3jkZ
TcM7Ptbe+xxlNOJs8vcC+RSmsQovsgsuMcYqW7u8TEoxHps5oTRTrQkwKs3F9kben5zP6WK9uYN4
7U3VSw2K2kBKLMmAp3ax3ZDh+eCHAijJwI450m8AM/nneGnkbIYrbUtMk/k1r1DI1+k1hchX1ck4
s8ZusZfKCdb7vyAPVSyuuT2AWTAGgKA7OWfbSZNd4B+kr3lvNDXMgFsxBqpi139ARyZuc05eJb+s
rZBzXGTLozQ0cKpM9f7SouBmuKB0s36OUO7JSKoq2NuEZNDxydtygQEa9xq/r8uFOSaq1pPVB6gT
Wbm96JM54LW25AaknOfVJ3J44vpCxqu9tUD3mbG1y/W0pD8CywPY2WqAi3vBAIfoBUejrCftdIC8
dBfaVMLLD28pEf6yJb+1CLiAYUQeoddPI9AGYU8Fz77DvvWrlj5/qMOFekcGog+BY4FmNMLNi7pH
gQQya41AUrm7jXZMCevcak2WZ0NaBexBBbdWahQI/tfoZ4yN0r8W1Cdz1jZKU5W2X3qg9L9DiW5n
Sw0b/Se3Hh+0GNmDog1vqYObRl69WnjMvdO1Lb+cYo7RWTdcao8G9BgvjygkUeKuJMTiVJHOXon3
oBDY3nDvbmm4gvt1Q4iqj1EHTYJWjtsyhdqThtkMaBmtFei8zqKNpsqjehiH59ro3GVsvD0Ojpwj
KcN0cIpwsF9ylRhVVeGWkYdIpFsagGd6wA9zYMsQr4RWwN0vLuUiheIWduchLXuadnFITHHa+YlX
A7KL9DCbvldHX6fU/AkBQAPZ/S/awYG4R9iqHkyOXYa71Y7VKhc2wEqwNt/PfLddWi5woMatP938
ZlLQr4PppAnEzA4G/DCSGobxYSjMTQ7Iqgi76O7/bNWVHa5wMnOtskGcSOwIooVF5Pze/DfjjbuA
d2I6EhXTyATYLM769Z+60QHSCuXYu/RAn7YMRA5aN2VKqEfXObxlLoZvA+WYRYM3ntxGvd7ysacB
V5q2uC4Alcwf7QjkjvF0Rcuh7KIWprZwYkcdjGV+I9JnXtaI06hyBL/QQylXbc4ohEnJwBcmZbug
CLrKjzz/ZKi3ncmoWaxmk+Rs5Esu0ykvJQnuVIpfOc4NQICy2QBR9QZEYsEzZ2NKQZP7uS9hELDq
pcEOoXmC83u9R0XZ+IXbklpsxGViuRaltuFqVBN/Ppm+eb3QnkjbOqOT2Sq8skr6NCbGpiAPjNZm
e1F9fu0gKJhMuPc0c9oBQOhXB8qpXzftfV9WAwSKpEM275HNJhYohg9UAsYhjazxbcOcbsz1T9oy
JUn5Ke48gOjidCV3sjWJka8OGstdLQPVKgXDgbA19G89t0MxgulMR9EEt/jcTAFPdGZPs//Bz8Lu
Trw+ewoWNXxy8q67JKVh5VCdtbiN3oSyF9TG2bVHwo7UDjbM/lmT/rEVSfw4ETAGpfAjD3tBK7L4
kxFKpqPZpzp/LTFgZl+hBUqFhfX9PNa46eV8oRoOs8WAmfwiGL8bu2vTWetzQ0FYsOchCK/sCE1u
fg6zA9CN55D7NTrwwetDUFDqCGFkBd7MBMUi+ZdRPD1o8KKmjAHrgMBqCQsU2KcsKPRZivbptKuT
mZ+c/iFkvxloH+79vTbo0QOQPIn6fa6bJVPW6Tlw5Tab5k9WxHVjdfx6myLawxRG0BrDfi3JuzKH
iotGRPYpFToMBijqkyOvWRSpN2iNzQH/LjaVacwF2bsQ+NPXMJlouMax1cFNceIc6+g2bSEi0Nih
Oa5Z3i1JYeJUZhnAk1wDcUbGhCLoZhy9eWm8YmIK3SI3GyMqJ8/dRwEU/GAWu76ByVHs1EX11qyQ
klP3upHArsIUWlInJkS5haUhWmHlY8tnH5EY8esH3Q+sKXGt+l9NesCsP7DVsRQsxDmTcRLkKLfE
cEpxoWPN91hNts8lZnD9u53S5bRoETICA/w2e9I1qKA0pBsu3NnG/y0gn3/Gp2sOXjSgeqY95L1G
L4635OFXlrtMc9yaSbXteoBh2YDa9Lx3A3RZf0y4GLVEtsYYZ55W7KKCYhjGFSKPVpWhx4Y2c+g+
8fHoNJjZ+g7gZ/vmpFt0Y/unTBVJxCz7Kt48uHHIJPC6bvxV62pdPzA7gI+kOVzs9pWXuzqa5MIR
OTtZxQzWRd/slG3kZ+vA5M5Pd7lrxUl5A4C7riTEXpLgbtXleOhnON6R1KCNYhKuNc8sTQYQAfmi
LoqX5CKOByn75Ha+L51rl0b/ocCdNNcCDTcjPSxmlzRVFwps64d0yt0H6kbVmBuEjSjZLTplPoxi
jTEnNubQb5b8K8ie3dQ4y4LIuNR8lUyDH1pBjQy+bJkvWXqSNsyipuj89/JJTLm5WRe+Xjf69e2n
WsnzooVytSxCQngKWamNQ++NRrigZK29KK7FIPGq3h7HO8TZai/oTEbePCEaNcYkQM2Zt9KEnaTW
VZa+rS8K7FggPv5GjmVanG/6avAnZYxnfhIHAOKfkImVPMAuP9bfZjYdTYIAOqlDm0anSlGdAVc2
JYGakUVIISDVWtmH4B/SoCMb9qZz6on10r27Kt41zQGqkd//daLrBeAALMsSQGfJRBEu97y17KAO
srESylivpNoQOSH2wVl5OOm3kqI/32nZhgLyomMAf4Lofyvtc2EC3kE564yBA7C8bLIEinB2Mo/M
lof3c+ngUn6lMSqWi9hU8YrRS3PAvrzVck2BACN+AyouSSnaa44yNAG/sOqhy/6SPVE13Coyw3T3
E2NHLvrlGe5AblGWdcC5Rqac1Bpw28BJGfTKmfWz0bpqIoo4qqTz3Oue83UtRrRE9NuQlfqGU+gf
izzoQK5MT8j1BMAh1+Mo3WQCfYvJJFDwuHBVZCFBDzQ+DAmkhqmglqEP2iJKytGHfV9eTb/5xS5B
t35Ai/f9XoHkhdeDAEfXv2vesXDRbsnSMF1B9hmDHFXmRxfl1OcapkC6h+Q/I3WaFc4R5oVSKFPV
nqkSy4vOlg9hl/N5JZa5cer5Q/erA7DRuFVs/1rv1Lh7Oircb1uuXxp+p4tx3s+3GkwQIIdVSdmB
YAM6itN3f5HxZvRW79/NW9AraRE15nOCpZTTlnI18OHOSZTxuwavZJxEQShUM/JI7Zq3QYZQtfvq
3Zd9coP1MRC5sRnpHUSpg8bWoYl0jWet2EN9VM7R6X9pJ2JXQ5JJJiQd2p7Rz7vdnFRD/NcJF/w7
2l9+zvaD2b1Cn2ZsSmfB2NbrhtBbEXz8XdPKqjW5oCfWM4oizvMLBf8Cf3OV2BrOpIR2Oe+WhD02
6EIDAzbarN5zT2i6Mp5LO9gUxOVCqt15QnfRIf+gTIKohuRhpinWwBSo9ZjJktD/exqgDnP432yA
GNCpYVFn6EBdIbR+1khifCq9pX4xj3x3sr6a76N/GwvXcGdDV0yn3HAdX4xErt7V3UtjBCk0C2In
txbb2/F//nKqEVzu2sb6MNDzyxdW4CYZQzSdi/siLWBrEYa48lrKDGNl7cpYxB/V4rp3Z9TNHjsI
4sUnSGeDsYDbFYFG0KuQZeyGa9LdsOf9EZ1sUYDQhuEdJylXEwi+8rewF7xwB0MahujkiZFgXQuE
bPlQbTqlGF32TmdpwmOZn4mlFIqs5LOzvrCJZyNcbDmiRTUfRKsI8qS6cGw3nfObPIQMTs2y3sT0
b9iSBruAaUJErLkmYpwcDc4Juz4RMO/nZHLwmZOi21e4ENn8f8II+RAFQ2Df+qkZIV8o9oZ3U1HB
DoJo4exqvM2/iziewmAt0Bp+005k21BXYt7HEFwwSpPet0nHr1Xc4jcgjXSNZjtW7/hsHf1GbarZ
LWgSz+tJUmyUssB7rVgpV2Th7xA2wcFZuutKEJu26dEI56HRHGeZOA2e+C5QroWj3NOWrac3W1zU
22yN/EgxFyk/K3M9glBM9xDXICiqNeRaNIN4Uesw/lBi3jY5GE7mxf4FzWyWwn4zcbtSNqLcz6L8
b3fKOEq5E2uKRYG6HRVo3UbTAdrHGXiwNGFJ+xizJ12xdRaFkdLv7LaMPgXx2f4kcMqXxopUjAgB
BzQE/OXvvDlfbtK3odnpoVmAXMd6W5Is9lDP23M5ELj//D9MibyQLyC5/L5b/0kSRsM7sEka477p
YzxkT6gu2pO/RZ998zuXwyYKiNdCH9l332pV7JSIB+g/UTfjGKOZfF93QmylQNonLGUQVRF143y9
D3h20Zc76LA6TA2rSaxQdF9PLlSW3TAY9Tw3EI9H6ghSjWfwcChb1JXa8aUTxdSxD5Z5Pz062d1k
+8uJfBitud+tbvPzzZpTLq2IRzSmjNKYl8SgaRy2qBzJB/PGdG1AMD4iEIrWrKDC0+WX23Q9iGtl
k+7N3QInDAztCLAVzL8cQK88qPhspXTmv2X4AyoEVMxC8A6bqShgs3ZZED1z/aUZvcVsv5q/nwpn
aSEkGS6wSZPLOZQjDZ2nkOPWAjqCkDw7bDeC08e01GCGvMZdLt8uDzVWdLG36cXFzWAewDhn7YBI
V0LXtVxK5kmsBMntOGCW5BXBs72P31pcyj3Fkl70Z3dsY0pvHzkMpY6cPCBSenrLoZ+NOK4r+EAA
TTDBz0TNH70EiIT5kJwk5lFha/5jtuN8LOhlHiaUYvQPvyMiSRlA/u9q1i0rVg0YIeuf/Pfj2hu9
O8xj5DVw0hhST5mDHBfGOiidllZ8dDp+5N3y4HqJIUSlth+l9sMmGfMSB1V3jxwBNNVcJtqoOGb6
vOdn1nY4CPBWtcPr//ygiGUE6QgVZOofbknUacGhicFxN6vj5Cqp49mXfJ5YeJtMtadEh0kYl8dp
hxl/dERiUrQRi16dHkKzd/EDrGRAKgP1i6GGJmRp5LvN6G6xcnhuZQKJ3Yc4QMLpTxFngiyg5Evp
CBPpGTURD4h927gq8vNNdjh932C3aze2Aom3G56afFIs0lOQGzaYCcuCS9nJ/rRA8Julj0vZDceV
CT0tXuviiMbfFrS4TWWjnMOVBcyVqNYURWtP+w4lIDyFxpxK+2JGM4rlwoM3sTBzUq+67SytP09u
1evd7b6poXPw2i11JJsggVrhGAvUwVHjbTpXTBWAPeZykVyM0YvfqGGaSbtL60Y7gQaC6qpBJys/
loLoFUPaVXeTAdXtvQT7EGLX3LBWkEf7GINXhJMGGKmb/JvJPd9NujVYGo71NqXkT4i7FPnV6dZ6
ni0EBAlghaOgsZingTO1JGt92PuPgmaiLCU9p9SKKhrI5XZ01VrDojiq9Z983YUlJnCI9glpys/I
pRJedW0svti+hnR1Qq3bmi1kujI8EuCHg69TlgL4ulYdPZTvfo1gQ9g95NNtnhgvyV9ijOeRNw47
bWbMNzdY367f2CIwlfE4I8sSRgSEpYg3hVAyJq0Jl+N3jy7ySizGwu1AEhLThQdipTSch7M7Z153
cay0cWNGYRlmENkv+oHNnSSvXJ7XAvfVYR8yddq4HbfMX4Y6OGHm8pZ7r+LD785VTXkrNiSR6JT6
wWcXVRlkrh/4vS8C3U6ui7vPlgCYD2IhbDuCc0gdreE3R66JpTKVVDn1ezbLh6oEDbmAr3CZhr8X
BpNmgu/uGs1hE0ZyvRVGLTVCPIxdnnoJ/nArRA8U9MLQ2NInyzb+vMQq24RWeh0JEJXJXwqRGYqP
S+pR0brm33CURP4yqz+iFAvIGDaEUKNs++nUL+pHdHf1GiZSTHAfT4gLP4pcWWqAcOgQUgWDNQSs
wpSKHIQrak27NuGjhpFKfnSmNVuVio5KWXigJmsETAFyGTDoMRHloUlnrSkt8rmr0J0GB9mQuHc2
1wlpZb/el2kfdyPCJ2pBVmRezRTwO+BhVoPg2DGiyDlRgPX9rgDmmf26bxg0gL08GBtkgh5LfJSh
qwF9Baz2Ew4Sr9KAd6Tk5k2+cebqzJ2vEU8EAgdx956KHzoTyivttMHIO3sKo+rDpciToQZFLYa7
SP5Jz2knlYTEjYUGKNdqy/N0qw9PqlVbWecIPSchnqN5lqcE/G4Ew9WfirlJzJdjDTbtXXfQnGqz
CXcdlX2S9hwoPBXu9lS+8NEvc/cOwFxS4xsvjmKG2Lb1/7V99pNgxVVaTBxApdHxhL98sz+ZYiK5
1b4a9uLTsyYc9azMVjQ6p3D9B+bf4LEtx1r6zQB6xQKRYhlOMRNGLTfMLwB9JrTqXRtH7yCVzCXr
dbN1d12uZmiJ2qhDk+FQD8vckCXGT9eIOgZRbSQIyTNEkLurauO95aMKpe03fPCxX2SJTbkpS/bi
+Lwmi8casVb+iQ1pOCK5mK15yzeEDQfOZ+YWeENjK7Ah+25YTnCB+Go3Tq49R3RBZrxHSlX4336B
gXjg3tSxVfuSk/V1u6TwpAIAxd1Xb8p7llueZxr4gphJIt+WWM6GoLMLTQbZUdxaxgzhqKbfFd+m
BpHQ79f4u9dljnN1rMSDYd8LSTJXSV838xt1fok4C9JFkGWCCR+z2TfU95U60xnOCldEE1hiEbzq
tb4nSY1PGVgHSiTvdagtlLO77fl2jBmhJWmBWQTl+Lc1LgCuCV7nnk1lopF18dKj2J8QHpN69wc9
9Ec6rC9C6E75RfbwsK3DLVyG9Wq8l7yKuKNSct7b8ma/Y2Fdp7sy8Gp8oovCcU/ydYGb3wvkjTBo
Rma+Cy1jowvJ+kTJQ3KoZDR1Bpcff7OgGvSPyMRK28UGo63F4K0c3Zt3KC9aeG1lgJHZUXJAzJ68
teVWRTPIVroHI01yMahBgH1dOQ0bJSfVFTSmOre5KNd694G649zy9jMF4CoEKPUtAUNVj5nD2VVR
9oVTSiTEQgVwKf165T5Fzf9xRU+kotgszw8VH0N9L2Eg0ke0IqUg8zqwqgORjZ5u66V9w0TpjZiV
GZwyw5ERy7KtImYUpbBn2MF7plFq5b07b4R3j/UG2pS26IuYFrCgvH0xvvJwkgtUAN/DN49r/Vds
Hf/m4MG2dAMPjzOkOgA4JuhuA/FgZXafwKX778fPzwicFYlL7kwiJcyXIPCi5goV6y5Yw4rEd9mu
R0qwX65nk+RM+aozmd18ocT1LgN78VpyYn9Ox0fq3ktFEZA5kC3CEmgl/pQU6dSNM0sEUJZH+nW6
hBBC9Eub9vqZFAjI/rJL/KQRvOaodAjLODLAHhQPt5ouKIpUyeME793MbP6BQfExGyexipViVSIo
PWDLXbZilKCIBUZtWVCdXpNdmPkZe0VYLIiqIjPuzAanEbx7M8NFvNMt8pYRRnvnNVwKSyuKxrgL
uRRx7QM3BLjPasACOvZ3WfZNbth5hvdTGz9iUyn+1qCwiPr1Hq97YUJhVumf4nZMkHil1yBv+Kzz
GTomzqc77qalT97raXvGdCSduRqLsaJY+TIXel5UoR9SbpHKOwW4OL9NHLCnv8UB0nOIAC0MGrd1
5/r2UwW8Z2XdT6GUm9lZz25foeqX2NDk+QkMDMKYCookCjti1kXO6tCQ7b4G5TbGy06v4kdBcIoq
oEPAwT+kMHEt2NBisvZK1QYq+lGaC1nQ1xF1Fud8xIKllFgkZgd1VDmy2IgqBEtGO0V/nHy3yerI
CkJNN1oEr8Bc84CLwai5KAB391tZevNVh3I6fTZvgSWDxrH8njfHEmxeOrf+2zYfx5m4IKMh2nns
4+RN78RW/+Bs1IsIxiv4Zjur3ZFqKcsw97Gypicf5XTTqxEJijbGQO00O9eiOum7rQnwv2Mn9SWn
+B8g1Nia8I0E+CYHp6Vt39fYHsVb/fBjuFQs/NWeM/JKFGUXNuWur0XpW7rgHGTRQEwk6pSX61d5
XS1/5W+5UQN36Kc3vW1ZXQtdutH5jz09IEtcTeByRp6KS1fcUGEVPxHRprp3o5lxfBwBb/2cjUqR
bBo6T8ZxkcrxlBi3LeXwtrbKW5zVM26sWIsPCXihevRIVOEScg9BWseFoUjcMVjxwxjqo8P0HI+m
oxq3LiwkmFVg8ybiuqo1gVkzUYa+0jKlHfRuXuoWgCzSPmM5XwN8NUmC1ACTjIMrFzuIZV8c5pWY
eiPp8lq5h5NljpnVxnRAAi8mHH01yVKfAa4W8iKU0BMkvURmlYkpJNQBakB1HztuKlm2PV464SIj
sfWJ4F3Tu1Vn5SR7Gev9CwKZ6qYAH2sXzF6JOAsgTqeXoX4b7u+Chg0+vaq3QsnIWrol8QjtB6n9
1MQ1+Ib6OfVkbu8oSQLKEXNA43DPozEuWuzAS+M/yv/jPpQ79Uh/9/SSvsyHBjWIhmrAGrXNQOkk
RMvhT0xIvI6fz/spTetYfhxY6kOHgETKErPUBctPKbFhJDeXced2W4BF+GnBqaFiqZu4VPk/iSPl
r2MibSisn1a89u5dWY5Lcu4d6kShzvb3Bo9WrZllh5hHjEfllHaOQtpu23IsUwMeAZgE0z7kod95
xtidD4oYrSFh9wKCWUDxp9IzzKz625sjwezjjBg307LUypLndZXaagIIIzkJYUXb8i9k27TPAdVt
DI11b8Ix6J+shuwpgFhhg83r+2ik6VLXK6rmfPSptFDwON/ex+zfysEhZGRlR+rAc79gqHOZtuY8
REcwN1hfMBfLwe8/qPrlilixWoVw4pvFfVTsqC6X3zHTSjKigo2Leq8AO1kaZX50IB1/3BxFRJV2
lwFFoEjaAQeYwaEYGO/lAW/QN1l7ULaq5djcXFP9h2FBHgvE8u0pctPZZTQdg7w7AMw+rMmM2SmI
24v0mVTLNVAfpfMRb/u0bjdQhfTT4jjFRWlv1ttVqKzhZaQIjmV1TnfK34dw0qfRq8N0XCSgqs+D
4ek6EiaP2vQ5FnwFLT9PdYdcHJLtRG2kjU9FNTwQSSgdsyPUru1a70bYD0Y2fTJYLTpxA8drzF7f
wbAe4HJTAE92latQ5/P537acmF2w2S6p8VxPP4ktDzsh4L5g5hZYD2sbgU8G6Zy12oP1zTXRvc/+
PktkK/hXkBmkVga+dDF9U0KmBjn5UvV8ExNAJW7YkslNg6wUTF7ZlSXW3smQuHh3Gb1xElyeXRMw
5VRo9Mo/MP6eL7dcsrhGeqZolgy0cm8g0fYaQWWTTUj352w96eqIBEHzrYtOnTafAWJSZbN7NMaw
RInNVtRBlvoPlZe9TMx9WdMI/ptX5Lcx8ICdGc8yKpdjPdd5ZYhzFuXd3GZFGM/HHKToD5aL1pv2
XRSskWOZNf94HhfxVzXXFY/n6kl+MdGJB7vaSmczPm/bN6dI9x4w833hjQMGoTsQncKZdzTmw0ck
CR1iRXB7a9eXLBHHy1QY0jGcC7ekQRA94T4cn1TUPqD+fcVG3PwKOcfS1a1LgjvqDJTC01cGi1T0
TNIBiarXN8ELx2eISk5BwkKEEgOTHOjzL4FusWtSq5F2Cv00gx/OQ7QrIymIkllB3dq2w6k2+5xX
3unPDSpfowxMzb7DXUCNItnEwRU5yV/IpjxRR3ntupSlZ9XDg6J9bv7gVgdzILghCRITBzREjP72
GcUEIsmGGu9GWIVZNlQOw8zjZFqFH9HbxjeVuFoB32ILpr5nKDf/WtPKa/RnRMHORkz31e9nMRfK
wHyW6qXJt1d+Sc1fBI37ihiiLkIvvlETklFAr6Osolom4oY9LXWInIYj2BCMhO5FoFCRu9onUpJl
F3QXo0VjtS4lokGtq9VB6jngDNiqHKj/kR5dn+920kctMohky6pXXVMq8LzHA9b6CexE1kZ2Pg80
doYO1T1RrRxwsELj8y+/it0j127wPl8bq4k5RuC9gMIrNwB/Al/GW80hM+e9iGdYbZ17dqORR6sA
wweCPMQzOMcNiXuVh7qgtR7/MwY6ZJzogf//D2fL67C6cb3Z8Xm+rOkd+m8PqPIJJjo9Q1rQF1Or
vww0GFeg4EiItmu+TgF8ASwynlq5gZWeM36F5bF0Q+l0ZXFMRtGAHpUvorWcRSrZNEAEMaScYsiM
e4WC6KEgaH00WOfnnWEZ7TJErBcM/7ABD1rpbDDy13LOfbO5oJq1TZRCxrm70txrBrD0a4ko9ZIj
546SUVv72E+UdGEu8Ol7pAfY/tNpRd925l6L1OQmm9mLhcx7fRHQJLXgjLxQhMj/iqUtJstUPZdH
yGh03TxsqXJ5PrRxxJrdPV4G9MLa7FuVygygfHQKrhqqrEny0YSi2/NSZDB47YrECw/qZTa0LyOf
OvaHawhAGsMdc7D/e96Jwd8Lve29NYIB5piM/JcfvBjd/sxiXPlhjxPtagOY2rGfZzPfY4f1uE+7
wTc8w+wsDDyOY9uGCQodk7PNkP+kJ2PwsWnO8nSH0Dt7gEhULLQCUbUrysaUkaJBGSSAglT0gU7a
3rFdf3OYfa5U7bpGqO0FYs5waTzznJxuWKdAkGRJ+d0NHH7KFbFckjqT/3x2WcEeiEsPS2O0/1t1
JsQjwOIg3rmE48V9ayeCWfOlDqQ3fQ2Rao73+meDU56bsSjdY6PeH1Xz9beoC5FTsSQmkq87Ogrr
3HtjHUS04bP3Ly3LH1bTXfQQds+wXNtkAKlE5z2abc7rTlJ2acH64rxBYEE+mUOFskXgy7/afiRV
nuQ2ysaaBaSTyDqTk4WXgMWu/yX7+nHX1268t8phE82xM8Gf/9JluOfj0H64u8Ynn/37bGWVY5aZ
87G3NE61ov14s524JalcN9Iv5SwnToRDuIOCOPL2Fdl06bm4Kw9qS/yFALRFaN6HNOONXo/kDPjY
2aklbUQB1ttDUsglI8RpDNJVtTSio1DZldUPamMYEUaGw4UgQd7XatQFxZEcqaVy1CjJVIXKmj3E
lOmuYQYXGCPdW6o15/k2Kq7JYE/KFD3A0PaWHts4XSm+FXWMF7vdyhTmwANRvD/2r2iFec6QlWBN
sQRXgkG9ZCCTJh0ZbGONanr4lwOVBj/KnBiu/rEOZ+rPk1jQdCT/MP/DG+MDHkOp/2H4YddjmmgG
61rzIMT1oCv6uMIUtkveusRzmqzEQJ7nHqDXA7kY3C9gg652PamJ9ty/Ccr0IMAtehl3tmJg/778
nrqDkmk9bYxaMwh1MvTWwrCxCwCRAQp2R4UIFVEw83Vmo85WFlCRo2rDywi1Udqw0/sh/0AdhSpZ
j0AwejVSJF9dLBXYLthph2KiGCjT7wkPdq2BcAXmDfEPW6uqr5nP9k2v7HllvSOaprEeWHiFSGAx
4FIQKTRKOHetQFDm95UbDOsIs5TpJMyicvoKy8RLrkZAOsU5nc/5aXOEFeGB3MQz7Q5qHQZUUG7W
tILh8vu1p0IeE0CpSMr0/oCxkhplphnp/mLbSVY2T4BPbqoeL9PWZ34wIAzB8KJhjM4wxbBSnK1H
2crpMoJ2uc3P1QQHDxL5JLpobVF0QvnWexGxDSPBOv3h7YtXRx/DoH1yKCNkUxgl5KhgDjIZMPpV
r8eCsWy5h6wqEGgSYBguSckHeVmYhhPCEwH9bBCu4IDtRUqaY/KXgRGig0AQbI3T0MkbwY5b3yRH
DH0QrahvfbLR/S0+6cXbe1NyD4SLqcQQcz/MZpJ3dBp+by7JQ5iCi4A4hjzA9kyCM3uZioIdHSAD
khUwfI3TaGJZMkuhYxtaiAJaAQ1etpHSxbNvYzP2cJLMlTuw1qXzOfyn98bdEC85upjSpNV+Y/tQ
zcO4EF4GUA9/DWNE7pCrZlqAZ1SdzSsb/5YubUQkT2YsQ5fBrQFlzOxic7wEpkTTd+vzcuSnFFp7
Au/fp//Jmk8u4nQByt1DWGFcMfOuyBjHTKfvQqnBsFK9LGm6C5Qpf6z69yHwd1DgPYDyhPIPFUiy
FPT1wCLi86GyDl2JAwbqEYgqh5h5l98yTEW5aXDBS3MOhGTzTCtq+CKjjBbFfs+CRKr7OFmHV9fh
D1/7tO/DR8vPMXG2oV4jV8OWSPD5EnqbnJNzVC0ZFfMuh62+Dw7eN5b+LgwLJ8HRAzNSpz0Hkx0l
GO2w1yZRy7L5jh/EfIdfPnZk/fvCeS80T33pVj1zvF3UkduRLmXbWtVhkYkMygzsQxyvFyMKMPdW
AoxDFd6NJuPc1cAgImv5fXiIftR6LMfiDx2hKGcQrnnp5my/sRs11f8O3D9ozGbT92ZUI7EjgwEQ
NYfGWAtiSXLuP7XaAGHCWICTxtXrVGOqOWgu6KWCbJypLtCbI8GyzY22ixEwWHgEwQ/qmJNwMmVG
nx+GGRcl0+djqPvGfNAq0Q7QJsKcQ/4piSlvevzbmAuTShgvnPt+IW+++9PP56Hq6ok0q+ck/TSu
TN064gF7OlOm3r0jqyl7BxEw80S7dqBMWcP7poIAuAS3crIEbpN3hlUfgCGpDtkF39xNdou73rQ9
9CnpV51vU+7PXEjCgRb3em2SMuZtvji0VmpZwbV42Wwici78y9ZgF3dVxIhJm46frMUuu1nhaelf
AjKIliNQlbWjZOlhN5YDX6RK3FXl5yGrssUL56IbWuK/qg2e2Hk3wozKENVLoaZDOcWw6CFjutU3
cRIVG1Q4G9m3VclQuKWquXKfPlLXAgDMjO7+9VLXNMdKywan5cDrAXVxZfyKsgraKXwI5Fx+/ybE
a0eSAivcfSQ6oyUVcsHc9qdXGZNHbh3xEy7NRxzJnL9x6uXGZT7DkVJNWjoWzNSzarPUIlSfXyjb
i9+E7LAVfOHTP8fTjWPgzzJWOGn7tkTUY8nUMkG5G0tHY8W5Prck4tpf+A4SJ2k27YE2YL0UXJsf
WFFGGXhwtdAHI1XHWAbAP0yTBsrVbQfO0wwfUoZ+qxKbMi0GcDLDP9XYjlWuPNxia3R3UZmqyY02
ElGYOTvNPsdsOX2O+nQy5UTx8fwMq0N50Ex7rmaAPjxpHbTr6jnuUP5mOc/MiyR4G3s3KLn2UpWN
roOlz7rEurn+o20lkPc3pFiWmvDsDa7++CAJPbtgnptNZg126RlxHIKFbyfxp7W8PRmb9RGIZXS6
BZenhVSsQYprhjSk4+/EPcXW2HczTNPqEcn2o9GhY5o1am5Mot1CveXf9v4X7yFQ92l5vYiKAl0B
yAZ5hj/AI4jFdGgZYXP4bSZkTZ9l/BttCnUgk8w7YWptCMZa9qEA3NBjQBbzMaohXILqFGNK7VXH
cWn3p2QTVPTld7o16VeEBJWPHF/Evl8Iupws0M7lyh5p33Ny+Gfv8li317g0qQJwYWutjzE4wnoC
lJFiFrtz5A02ajeYig3vt03p2jnpi822ilY9ZfEZcEd8lX3EdZdOvr97ioN1pQ3VenZhTGzOebya
u5hl7addiz7HkNLcSUINXhqjoR6BCJ1TtZcnfLzSgZtc8WdsfSaPyLvEZuXPKBsQrGHzDNuPZr7k
FeVGPSYhN/XYVw930IWoysR8Z0MI7K9xzV7Pi33i+lkenHndHLzHJkhUPb96W8ndFBmWWXVHKkDg
Y8k8eXWTXLQuT9kXlAy2q8GzFluATuGHRLWrzzR6PmwhfMh4x8ns90+bI8WI5RwGYm7n+S2r1wL+
rsJs5QiuK6bcdU2eOzfY/GusZBlQisyryu1CpWl5UkioH6xTc07zkzmsBxauCv+WdQSw2RjbqKcL
XSe0XVxStjJJ62d67VXOLcl7f6SU575RwhTfILJ6y2lKWoSPtlyAIKMhCKXCv8cqUSQ38JfpCYH1
n3zrHYtsLNIYCYpDRM/7cGt615U3nvvIQkp+0OyeD0RYbgG0kGyY6pbM3njpe26CCH1JMPBVgqf5
rXXRGyPHe0Z+DtDDZnR6JrdC/5+3yU5rEolh9WicIuH1Flhch+4WQnOyRyTYTxrgpV8zPzCqFiLN
amIa3C1wAkscfzCc0rXad3ZPzUcB3nNlrJBVdTkGM+LewhNzXGo/VRGwA1ZMNGsa4RwsYdlZXE5U
Zs9D5WHw8D/UPO2sIRZJWmvajdstWN1VJLRxl/zj+my/lMUsEoXJbFwJW4H5yiRJEkrbJAoDu+w0
gLrozNudf0/+zt9Onzgwf/31K4XCNIAcVY4PhatICyqltMxZLCW+fRFbn2CPgfaPsRpJk8BFXJrb
uNexaI2FqOyX1BdFaiPVMRyPf5Q1YTq/X9uEBijTSjM5grGpVuXsZcUXEO9+AOjyc70bYPPX47tI
IchYZVZeANE/hMtyLjY2fGfN2FHoKT+VpAi5OhWGAaXxMD5sjowB/jbphvG0ROpzjwYlnuwTL7CL
LekHXfAQUp503gFWUUKNgAcR+l1PUTnhy64zVJ4pfd4GFWt6opwVmraerCvXn4QwcKi8PmkXLWHn
rIuivei9lpe3BgdtcCWzd0fpiFWB/YUBMNHAWRHqsjPYl0hq0UEqCvutn6LPZrT7xHzwQ3MHnwox
r8op3tIwKPuIvevvf3AVJzjneQ4WH5IRhv9xKv/8jHTlELT3fXsSB06UE29NBUIED7dh/WndibK/
rPGUSJoQjxpZahkhLDf+6kjfYOJ9chB6J6ET8GxATuagU8pIlaioQjPPV2MMDE/RmGOqgT0NoRjY
APSAsau55aq+Ujs9X/8omq4sxvxCeSgpe6jj2o9jOH1Hel6XERTtdzL8a1RqfolwuoZeo4+ffdQC
koiPDPkF+7kpKK/vjHNhiISYtizAtemgBNQ4unrbkKRnZ03GTNk0cMJRyhcSA6qsM+g2GSXg8m2Q
1DYaoe+9ytcH67CbDZqtfVCLhl6J/ddAhAAMtLbbA8GUF4OKZuIRw0oZOr01isi4JW8BwzjdCAhS
sQjS4xw66Y7NRkadDAuvVfGMNR5MRv7gFakyAckb9XRnCGdOOhcP22Q0flm4fVRA1V0qJgCzK/xB
z/wJpjnLtM4uLUGEo88ldk4r83nVrPYUnAFnXDT3VxiIeOQrIoiqr0TF4LmjZ8isA+nmft1w/h/v
BZ5XoBXz92a/6JQX/xwX85H6hqfBD6pn1oYeuEnOBCh+f55ib7YtDc5qVofeYBKN/n2C6SLxlyRH
i6flvdPkb+uMPeYVna1UVjLLS680c4wftPIrb0fu8Zb2IKSXKtSQHZGlA4QIut0zeWEl2QwAnpP1
J8itE+M+bxd/Wu2vh762QFUwsCB/bqWj9ThlVv/7t0b9sLcipTJj+ocjCaoQ/nP10lWgQC3sSGti
ByG1dwUCKnOElkHGRI7JZUd+zieqhlUeD86hYug6tvZEEQhC9DOHFHOUJtRVJVJfOgsmVYvWK2Fk
mXh6irrmlQjE+WQUksJnHPr4qLDL9oxi70Uq1O5638bihnk+rWhgrVwPjSzIDt/eicjqAXU48bHa
ATXY/HShVqn5IoG7MvTczc0fgLfrMqBTYjV0+TAYNoauUqg/h6DgVm1oLpFrxCUhAplmmkEEDxu3
SzI1cTg8n0PgOhZShYxQWPuzEZV6cYIu9FOwT6rM71jOwdvYwYAh/S19SeT/d9AOqLtR8l/5oeqZ
bBUfIEoVM/Htnfv43+x/DS+SdXXYOsDfSXEay+jyCNhTc5QQazH8HVGFTImIzDKcJDYfGxUFSHeb
KvzX2u2ywYwMJQv2nAZouuKqofyKrOoeJRRtTrpsndlH4kKvwsgVhZjHeR19fPVdSn+j/EvZQS1g
Feru25/Uo0y7mymBMthrq5k4QsLaTAnGloF1EoZKQ//Egyn7Fvd5YcpNy7kTqPF3Up63pPg1n7Lw
DIYPKrlScpiTbV4SwK1kZpAGKBkLE7ge4+MCyrBk9qDK+NIxg/PFVogGoQES20GfMsm9OC83MjZ5
5czXxDNGpAn+qgd+54SBsSzEJZ4z1O5hpV3hmGiI802wbZYyjftARo3R5b9/K2j2Nt6Z/PAGccpn
MepBbWGRQxOTeRL96ybTkmibXzYUOuJThU5Zkw5s7CBKadkHZoowNIU2cZBVZYyndVySF/70wN3b
nFtJV2eguE3hhWHA2pfeg7TeWiD5IqHZi29NLi46NQucqstviuY7cYyyFZLZ2psVrM84HAWGF2y3
jYXp1V8l3e4LUFRqZHi+apqgZoqBMvSf3F34GdIyyp6iiR5/0PrCXis55TAQYDV2ePdBYBtspa1V
RObmcBCz/hLNVQoKn10MmvW8S/NOWHEgWVF1zK4mAPAIeGr0E8sl8ic986IW6EV6cXFlG2BRPsIx
UlEbctXPGI6CbXnhccih798ZRsnZ1KRptNtcLXFE3PddvfPa8ftwGXOIdRjK27FBRp3sHzewFXNw
U0Q1bgF85U+0j/RQYUIRolyFkpjLGxHlhZ1JXDI/pSuLCg+C9tnl5xpi2W3npEQFGxwoa4mgiCVX
o021XW0lEUv1NLk9vQm9QFehAKWE0RcKdhdp6Ca7Se15qzlJ8aWvYGN2uFkzmt9Q+SbRaDOE52Qx
geBaXhIRrL1gz1D9OBxo2c3GRaZgqtipfdb7vYbP6JShjREO93CW8ERvQQUlhDJ7YaXlFK6AOWba
JLUqnhdfhCDfHi7rnMKnw6Gez68Uf/D9tAYQsyO945hnbtNT/Mlfsm8xmoKbEl9C78TnYu8LpLwG
pYl4plcph0VF1o30gpVj3D0mFrKhUJ0LYSkmHF7VXuFJGKf8dj0/Kcb12DLaif3ldeNlOjI3gMJL
BoqLZc8EpfUrQpVUTemrzHWaI8jRqIGWOdKoZfPlVWxMwUfvzxDsdc1amQXP7eBXvAkU+A++8IYb
k52mTpgFAFQ4kRQIOj0jNdJHL6raap9F4s1JcS6AifWWcjCOm1H97gW1t2leMNKvv0OJhMD2Y3Bq
yY8OGFbFUklsdunxlaq5QwrltikWUWf0JtqCkUKlRQi0ch85RG1sW8aonpp4azETh0VHcqoNaS5U
jyjMvKv/TgKO70u93yUxZWPZ9y/DTnYVoSVCTa92AUGMe6BQyW5NkJ8meIxERMAWwk3I+3XAmek2
xsM5mHWPPyeJYiEcNr3ki+3Q07iL6M2mzMLhf1Q0D11dk69egtbuZCr2cWRSr9y+gIzvv3xSkr21
g77gyswVxL/RVyJSrdqh40UItmgAvfOF2AuYEblu5juK5ALuQVSo3n+AmcufF/iiSAzxFtq2W5bt
u6vHYPVnSqstAMIUcJOcwaT6gc+xA4VEq5NP8P7fFYfRrGK9+C8Z+k5Y2SU+vq9e6/6fuFn0GFYt
0pRhZPsrKku1LKXDMpneWKL+bfuBtwOriY/VjKwkYioWZpdF4hLUnJp7mYAEJJcwOFYs/qieHqD/
utEyOsGMOOvX1tqZ6H7JWJiYmeR+aLr1Lijom/hwsi9qdZxtKXuGR4XB8JgrqHINGcVEWA/2F2vp
FDJ58bYoC1LAnFMkoYi05Bf7d7C/2/gD8rMysuZ1G/y8ifZGCKBy5H8358rsHeJ7HSzbwz6Bsj40
aSYll+0bNjw7pilmj0j3hNKZ1ZaW3XCAw3+MC1Kg2X8VHuY+XGSn7Z61G3sB8d3/tTcvFVmOG8Rt
3k4Dg/OavdONBeZBdQIOfzCcxKrCuhob4T9dTs9sFyCy9SELLIu3hGOonBTm2HU5GiCMYAZgl9/P
opluxqf6xxEdUs31R4xRsFkukHYotnzua2tprfez6YLnWeasGZQTJz+jKqCvKkFzY4M9zDZxDsIl
LqnMcVNLtHfmUkL7QETssG71JHqy/vNv47+FBT0Pv07vbxbpaNfZd7lhrTzPxTU+/qYu/CUUISTB
0F9h6kkOv0dd77AuAPDUZhCvpg/vjf86hQ2z6RIdWpLaOnr/WLaEgbVoUetsF3tDDp3MkG/q7aZ9
9fDiWrWv128N0ob4n5FXaUoTakl4n9AWb1K6SWyG4Bu0GXehYAHUieUqMIGK81ClDWtaJCxkyvCp
Z23jeNgVpuHB/j5h8CVVQ+dDEkrgWw3tQVaHBmUDKZ+hJWSM5La6feBSGp4+UkDadZV+ZwQfC+Zb
Mp+RP/IUH2pigNN+G+F4dDOybswhYTY4yMG4KpFUkfeFgSVyC1F5ChdX/Bh6DLV/l8BwnPvv0O50
y4IXp7wPoJ5SG8An+l85lftorwAn14Qp6MjlRzto4MeYL6S+uzLHkqO9tYyQzgiZ+HtTjMtzJEs1
DvO3zj5kssggWqwTaWpurKTnbUIphDVvx1v8OFMtG8w3bkyAuJebfj5aBfiXMxdtX3hwZzcwvCjc
0EVFkeQZO9iwndJ07fuSDBTCWMg/H6qtagz/NTT4BGCN53xWDaEGpzOIGAKVp2g862XuVeBAL2pE
BZs+XLKcQeu58ZY2ZLh88nzDJ2W9kkjgTYMDpfUZSwXd8aPHIs2fgCL47TsCoqAq7hju9ExyX5Cx
BNd1MP03txVluoQPePZoQFrV0Lk8q4HTIMfuuRKeDuIB2Dm77tHmpLkjB047BGX2Y5L5D1S5vzSM
cTSSx2PYYMl5Yc+R+hTLNUQYfwMd/ZvQZhvD8UjRFqKeNA/P7KVN47e+rTJ1wPMD3BeoNEzHnS6h
Zn1wMTDex11fHvWD86VmnJ90Wo4CxdzEAjyOu0A8RIzPDI5zVFvkFrw+L3DwK4jOgEEwKG3eCxNY
6m/2Ca8eENaVDZAHd1XWy3UMLKSOtswgF6wQTHa7KM5o9CoBuvDdQfGAx60mMX7wxHqB3+CfYSZ+
0MsawGkhM428+ez3hy+MlXxCRe2eZK+E6OhOfp0rgjUAS9jYBEruYlNnB6YAeyYBXVdRFEQUJjtu
pOsFvxF9ozgzMrkhuRvHuoiiZ0iHGNDGxxJ119SKhRR5Ep7R0FFM3ZNLE/hRMckSQYoULKKgVvbl
+UCRW0SCBFGtng+G3EipKPEfgBMZOe7PoP3knDWR6VjhOJoTnnTDYG9SyG29SI/kyfMlftsn+RId
BghY95MZe3VupM4Nf03m1p3XcMJC/hgKQ58sICTG47OQZuuJsmwEhLcBvLGjT/2bZrl9fI8hj0o2
KdG9kvXQ8JvuJjkwgtBU0q1EggfB8EOqIEiFr2Y2Vnp+MybyYSNl1973OKJtQgC+7O8nPHImCovE
nUdNzum+sxUXO6WNcaCmkYI9oTJiIzi8JiVboO4Lz+k67is2FX/lSWSNsisJxklLXmqZby+RCbJW
Q1cT+R/PcWkqEo1nHiNKnM/D6MX70ovt7suqa0tVXuKl95u8ebiuYmyyvj9vmwxWecMy40P03f3d
g4aJmGB6h45p0IJ9u5iydwjgj5vDucYWk/EgKbKxWpQzacE4dEFIDVbVuPbwU4zjk0w8/OeOvNkJ
NQGuATaegUJuBV4C1w3HbHbgci9pIY+tpFSeKzZsRaohrAouGqMQXPYZGM10wqJoP8ckL8hhu/Nt
WsDpXnEh/XUYZSZROk01q1lQ7NvzfE6eNRp35YqHR7gR1N/yOnlLeXhq7te+WAyqtFeRgI9S2vL+
pnIrkBBu27mgM6Twe3IHA+mS0j2mCt9krb9uhoOxYVgWA3SjiahtlSMczI1SlUN8pAqQEb1RfkIo
fTnEMZIYBm0BFLqgr2tLeRWyqYSdPWOGeMazQvAIPYqGb1yxEAn1dfWNtTTN5ZAdckqqs2lnKCCt
VhfZLKFwqEWczSmitSy1G4UubfvgZ8nH08O0cFGtUnW/grwh/OJN+sMUtF02mWWsQPjw/Z03O+tw
b36ODdOLLjP+kznGloNYYn2J4X2TV6mz04fI23W3YimHIolos3+QLhCHe3CCADU4qZ39cQw9GdpT
Xe3fLVw986uulsXaqPE/af3Th3BazVnKn6JHS9nD6xg6zwN0BxeEyRp1ADSJxn3cvk/qnX8Wv5X7
rKHp39ijYb/e/BWPncZ+XzAOjEPc3ZIbH8x3/y1YHuETIhgWPHz+3cSeWxYvYWbyxqwlM/7n7atY
kgzNEn9D6khdWNQh9XepGObR97TrCcNQJfcNwaVy4OpXx8/b0uiNvlrgNUoqqDoXbGRqqZ+mcd7H
lRhpCJEsH1brX0GejzNHKME5oWZMyrc82ssp5Y8O8gNk2LDgDSrdYNyTvTRQuuDswS0FsR3yV/lm
Ua+wNZ5rsu8Qh7GDZzCAYuH9NZ/x5wNUkDJpgvfTAij0GsNUVn99yK4TItqK88X/69f7s8PgB3j9
/gyw5P0t+l1TehNCj9bV4Fw3E7tWVA0vcBPyYvTUMByeBFjaTt1M1/dQIPm9FNjbAMA1kDn4f1Jr
lFxYywJSnbwAqfZU7Thrr7ods4SBjn93b9nB2OgQh8XQCMWsRTFRGRYMJR1HCuegdeP1MLpZVEev
wdJsFrrv+DIfVTF3wp63EF23B2VB5rngLHFxIYojKYIzLNks94kAWNhE+ZCfc7ZRfiHO42anrEag
ZTpIgUzCnyfzg0to4JVtyYxiXITlY7ed/MuyLBmxI/GVcRldMTXu4yMEZEOk0SR0QldINZmpZ/VW
nwb/URtYNjpmsg4lB4GxF088iiyblr4zL3QkG4R2sdf6pwgicNZQVslZjNRSWF0dq1M4iGITsSDj
H74hQTWVavVoTUXuPvxVAY+pJNxjtoHkK6vNYE4rDB9yLTxBQ8zYHpiH+bgWvY+PtD303r+JohcX
sr9SF7gmeDBpPCmkhYNK3Snnrh2WJnOOtx+NXluobhj+vahbT2k3v/+NXjiFJ5yJikz//gVwU6XV
Vbdx2inr5YbEyU1CvMAjuIEaSYfQCakAvXEojUXgAUMerq13mgi1YwzVgQDeRMzhtZDOnmqjaKat
xJmHa2sfA8zpccb6T8cn0aG8tp6USsGZQnaGrgCq5Grr+DN8i5q5bqDf4SarlVgfl4524NJhND6K
GWD4p6Lkla81ut0TQmz/tpKi53Yxf+lT4IKvDfSXfje0rWA8pwIeEXDXyF2s6jkNlE5EkRkOLbcJ
X30CmxECHRbvvCuxZ5iz+v49Ij68QEadgdF7z4b0jlO/i++SZNbE5Gn4G9WLP/kITKLL/MjDQFoA
DpOBZCxDu6wzREaQWd1gxa8KsXxPvYffm1iIsIGzooM0D0DMI6wgIO+xUA1KK3XCF+TNSMOyXN73
u1+ByxNt/971qJcYDHpm78QuVw8ZwnWNlR5yCznzd3imO288525CKJfU9KkrlUTqnaBXJt29gQsL
KndkjJ9dSoEPDuWYSfaQI4OYJ2mpqW37Ws56J1AxTo9ckGFmj4WDSgguO1YUXmIljFyK4NHHMb4h
zK0fmsjleYybTBWbVSjuArGrwV92gg6YQcOUA3mY6h+w5tcwqf08g8bO/9u0bkmJ0HiPQQFKoLzO
A/nbihBU1/FK4rNkgeg/lycWLvwCY55KRh9Pe4mNuPCOh8LtAGZo7sa797q0QERK7DuA/2UrpkGQ
fOJnwRsbVKsN6K0NXz6oFSNRnByfEsh2Gxb7z6Os3pyN91EJByc9qsv1dhpdMmTy6hqQMpuEdSig
FPPD1XB0AzQOWIrf5DvgfDFfDfx49638uwBpnnBmI0nI2nU+QhNpa3ojel+9HHqrnOHcqatPJiZl
7nHMpihMyX90WTe+iAgauhPKLBffR6EgMx8yERwOd2aseOiSe19zFSsylTgyBpnL/p2btAVvevYQ
ZNaX7QMUWsxrk6K6MCDmGt+B/rVni4vMsiCG7YtILCCLWP+PTZNiLkUJZ7rMJ4jLLEjFWVdQ2Un1
fOKzrL+thIwy6NvtEVoBaR3ICrOXhfo4hryIpGCmxq9lgDKeZwV2Aobtgcdxln9QGAIetpg9WNBa
eY7CiCLn72GjArwmi4fKMrYBjXxv/4aRCEbJl8uAzBVvzBF1x8j/nUjIlZdMREcZU1Rf/vnBcITj
vTgmU1YK/Zuvj4BJRV/B1kH5TQmlU6lni4Y0JGYdPDQ8pvJVpp879gKQ6MDVbQvPKagY81fihrvH
sC90eCgiGqhTlWqxpdvc0MYADVP3KXXGiiFyAFIV8I7pQfRhBU9tiYAvEs9KSc0IU14YmBZCr/uv
b6jC8fK+5Xn5dgKxMo9WV3Ctd3fUeDqxT573qYJd4RXL819CwGhGfAPf5m9ASh2mgPs6BKNDM8WD
k0+wRHj9kzwBjOwa5sDTXxfiBeKfy2DyfEybvcZeBlBocrK6mXR3BmQZd7nOVCT0PTgZe+4orjwh
pQw3cfBcQvbJwpg2pRjUrGD/HZD+0bhdPmHTZNCza7QYvMsqYMajq60WdY9D7IRUuJR532EIT2q+
0NB4zqCJQQAerV4hWC17Z2jHb2HG/mneMnp0c2hAiju7KmoWXX/hGyICNPAl6JVmpP2Fwwsx0A9U
qVGcSoyICGiK1Fv2j4w9KChf2EW5WKDdJC44YzJfMFG4h2XQOnS7yDFVqLnDzfLXctC9zfGC2gjs
I57bjxx3PUDOKjSKTnZkj1LaV+eE2/t5PpL5zGg15qt6tURPdojhJDeCrNbbLAOl667/CDdnirTU
uhgYnPaVEFdK3v7S+5VsbosWqIi8BEQCjK/X7JWktSXAuvDbOhS/zciaYzEQcvsVfFnANktRVzSx
n3d5QTCRKWxO9itk+mEdaLze7QUtaUzSTB+shg1kbok4tHAAwSkNKt+VD2X8uINZ5D8srwQ83TyM
+aNVr12XN0xuoT2enx3cUzJqLLGI2tmcvVUej/kYpHdt3MI6hsJS8wGePrixMyyja3m4MwLXrYdA
C35gFQnGTbclm4ziOm9+u5SZZu25QPfUFjP15klTjOynUaAffU6CP9LtmWuvTwNxCN0loNa0jKI/
y2M47fa8fum9nefIaMmJVbKBtuFakIiVL6H+53eM/tn1v7cyoSwo3wuIlQTroRWald02ZWUigteE
LOSXXjXjSvxotHt31uGkSOS/DePxU4VvcFbZrhPdP2/cmqdUmi+AIx5SPM0Lkjmha2wUMDYVmvkQ
X7EeQaTGe5aOU7P4gZx3sSK/f96tj7X3PGa8uGz/i+yjvttvKRC6f/VY/6sn6TCq06363gh7GKdR
Q+VBn3VU8oUDNgMiB0c+3ln/Cs778G6YQ+rLvZu3lBePhb3U3hR1GB96NBL/g72Pqn5dB8EqXOs9
Lp67P/X7ktuunG39fgldNB7BqxIe1pCEAnocbi054p3dBVFHQV/7Q0kvqKM+CAWfVqd9o+0rOQQZ
2KHRQsjmqcyLFl2aZo5ME8fLQYYtqE2HTgxEX4t3SQcwPKOmFPHzhqN59n0i7jVGcUXBTBDriadu
uT1Dev73R4olxzDnp0S77zmLJ7De/vWU/HvUbca/dDT6w+1EZlT9G7ZBlt625K4XgPrUCjlg9LMg
VeUMWXHSYlKh/X0RRxsarT4Z6curhskLZL5rArVUu2d/Vj7o5m+elwaUXIZlJHHhJ/ov0rtfeCv3
LUG78IBajKPaiX4Siwu9cqwWIQtbBtT1OnB22MUVB73tQwbIiWrQ0nPrAsHlOoqqno9R8rCNIGPs
oWCHDPinlmDIL4bkqs3RbKQPQyLwG9mkxXSiA5PKftufnwK8z7eZ9z5YUK7jsfRSg9gLzgoQ2f7k
KWtn2xdQ1duPNAlOfjL09QdLBEUKFwf6zN9tFrwPs3OsvfSqHDDzksAIHuuE+5VbC2rqtlPvD5y3
PkBMSatKCEDVLub23OkWnStR3tsX2fnJdxWF1LaPRuvRxRUKNw5/uHmiQQNJ1tNx4USXNJi61Igi
uqYnDBL+3ZGM8S4c2hTZDwlhFbvCrmzzL6CPMzkfiz2xhRj8KZvXRjsC1LOGxAvuP9997uxfgsPV
2pircAWhRFjBnvithrXWv9teKISAOAyVOAZlAaebuW5UpQReHFYnhrGFmENgww1HrcI8UvCKnMxC
gKSLphjphd5ekQqeig42v1+tY9GUFc0l2NblbbJt041Bp9ew1R3ccQnBgO2aI+tuc0DsStW2Y31k
oSIsWAHrLsYfK01UT3eAiaKO5Sh0j2hpPcdaBkwoXVxkM3aj4vydZs4o6zneNesXgnxnCqaazNzd
nU0Nae2lhBU++rs7b9ehR6BaZGaXoPSq5VBuv30uMDRXlvC/32cwxenLeOBzH095VOnbwosIU/yS
R8/A7O0yiHubFStklIHrySjk8ZxAgox5g4VRP8e7sOz2Ru++S06NSXuJbxLGsN7rr/611x0h/5dM
gbQip1xAxvOVeez3H8b2XAwdmPqFJ5lzlLQJksv+jEgsfnrHfSC6JqlxLx/xcP8iZVzU2qOoAAp4
nNjHx4Zmy4pdyMnJLzBVrU07dqbsK8hNkvdIvFa/aUOyXO/Cpmkz/ju4klF4QRfmMnvnq5u+NoaQ
5a/Uky4YVTssOVWIMBSuYXZTPa25hiT/TiZ/JoMwvJylqfZv8cOL7tTDVj5i/zNW/4GpTwClAtGV
LfCTcX4Va6lUjIui6kQVSMb7R9FDJNdO9XrNTyhUmJWaw6bp4tKipiO7qTRlVH+FTFLdnhUns2T9
VsKGM5U05wN2J0WHcM2QW/x0Ag7k5/3tkjegJuFdZGjEA4Tkpz7xcPRZLUaNSaZdXtZ6TlqtH7Pd
9K8zExkODZmquvEHvL6JZZkGse5z8JdzjFKC0nURhCMRoClUqlxFxAXeOjVm3CEWLSJ1JRW9/dty
gOgBVkHOakFWq8oDle9/r5MeK9rahu6AQ/9JFOwPpd1653dYu7BsUSl8HvqPJnnsnnhAt1p0UqEt
f7+/bXNNXEudH6Qprel9EU1aEe5ib3LjYIH5GKVTxUo/AbNUo9jZL2dJXUvIZhZZt/eSaVloDpbW
mzzeMz9MQxlZy151d0w6G0/6vEDq71w0E7GOxdjSjilbLPr4mA/aWBeIKLRtE8h/YDZSBaj/77n3
mryZp+x9h4V+UCC3QUzLXkmjLFcxYnqusHF3sWuk1wD5N8LU3w0rQY5a01LLDdfni46H43To0i37
DseWKo2zFuFU0BIVrNoOaETDuc6z7/0vSeCoB7ftPw8FEiqlu9DSWwabqwfnNEEQZ/CA17O4iPwf
xzSeVMbR4qzXMxoaDIk81XjMO/E/+56vYyypr4leiykS7/0OzAYiAHjlfYZJCqON2tG02gur7vYX
BdlpySEB79OCiei0FbRYtpkiM8v9gyMP6USJhn6ETjZVI+yEHWvjsYm1jNsz43ZDYOio/vl6mVHJ
vf3yIbYOimCEiQb33ryHeNXeQE/jZ+ZVtJcnFllkndExt7QX3HiT9/nhh4e0G5+d1sbq5EFddGVj
F+yR0FoaVp5OHOSbZ5BQ+6oMux4xZboC9gQUn9VI8M7SXURD3SdeuDcZOBgVhDcir2PmYT2BfCtI
sbIHRr8RlEs9VOBMWSizzxDWwrFCWA+CKYG+3ZIhVOtP5NCJgeN2CTCn2p76+7+hoP5VphCxaJ0U
IvXViZmZ30nLRezt9IRfM1TRfrXNhvrspikWYxfhwfOVnxoIXOxShUCI1sGeTVUjPUW52N8vef0/
PLBh/hX7EngjgRtJq3BpQ0V89xByAm55o4T6tb89A5Gw2zXbrYgO8KGdO2VimTqWmYAzn70ewgxK
WgGBKo6Z+TSHL4vvVMIh22exZiO+OCJh6Nt97zmC0OMx9dSi+GHNHjz/oGMajBHQIFgmfZfZNPyD
0hH3n2HMNrF+aPrvocmQr67or9a0FSJfSMTslQ3pTKxzx3AN+uVMMwtmn+ClcgwXqyYPPUo7oJ8a
LYQ5VYqFtTbk6/ki+NIR1tyMgNTigL+vimn+uk8R6B6KL6bzSbaKV4Jr3ELPOnvNXKrAxYAHI3rB
45wAFTOVKwlvVdvTvswcNhHcIvVNGHvhr28HZVhGZznmDNxcG7I0uQgfAae8qf9U5VRhdqInzP+I
woNStNvXcz1RyxHTij6JytCSnjB4icSX1c74xSfmciLqLLQeHEbMFh2lJJBYwfwONCc7Ff2Nb0W1
COJBh2F9VMjvQvMtWnKBHYhbC0VwEsVkN024veFy1dpOQX3CxG8mIrluTrP4Gkj6MerqyIqCqX+5
9sHLhfB+CnWhIkMZrtrb3886po2p8vhINeutux5kdSXiM2fIoLGGcJkCnKwAv+N8HJthn9rwodo/
W6bQ/Kd4uSP0+zrg6Lp1s6KZOGTSt3Zruz7YA3RrwUNNcHkN5bEO20KXuqfuX3LLFSRbi7p3QNHH
g/odLAfKxXpQChWgxBP49bxZ1tW8qtudn9OR3FZwP84tMTYpP2lLgI4u1yRUCTgQmvSpniQMd/ou
u/Dw+xdw1T3mTI3UAs5/A91dPr2+LGqL7ptkiDfMXvr8fnRNC8jq3j58fXoHmJLiI+pgz8y37vw4
//n+qNvR1o/BksRqBIRRiebVdTyHzcccty3BXrxqWyjFRpLdTX3Y0t2p+mQ/0e1xU9S7nhPDY8O3
IAfl3UYxxDfIXqh46lm3HsrnQG5LK0EnarTb1iFNwtv+WzUU7SOs0kbl78Aa7QrEyDNomnl5iFdh
UmqjUui1n4Pee4wO0UtYd+/rWqcebwL0IiuW0wextipg1GygGM3u2K0AY67U1LT7b6zUXENDc5rs
o3B5uEaTzu2WsizwQS01nJ3/ojW4EisVGwwd+eHmj9L4FBwT5gD8jsPY/zTEwRQdr2e8tV1e+eWz
DNFgkez6rQ6LofqWt+ECkm1kRD1xHwklxEuiolwUBYngAUQrYLcc2KbNuOCwYno753Pwnhdbwr00
lGIRguF1+oRQHcgjNMxKht4Sm82DnjJ55RII/pHW/ofZzcU8PAZsGhJfDmS7WL5bQwdtRcPHi6nQ
Zv5efhaTGwsN7JdRohOwAyyIcMqVBC/QuUjauq/3+NUbLxadENnx6R15aOLN2UDPEerBx5IlWsXn
oo+taxYz/WTLuah4/Xmjr/cTFli9pSXXNP0n9ImvX3oip1Ry6VU+BQjwNo189ty1swAHhojww9MK
g7io7O9P6JVFob64poL/rTWgasjz5JXFdPrexSs52yMK8c2DvHYhm7KpGil227XseWreUOCJSSA6
K+Zmpn9BAn+kN8YhlqNjynZBsAGx4ASmSfhTPlha2G9j0AQCAOL1O4ovMMJCFK8XQ+XwnoNoMa42
hyQLccP2OVOiUhknjeF5RegffQD3SlsxIg1mIghiEq9T2+4HNS3Sz6xQ1uOc3Nld96IbBVzVbqzt
A1GL6rxl9CIEuLl3/U+PX2KAmVmWlu111Ri/NlXopkM0hck5vZ0lz6ubPRAgOI25+0+XEbSQ69bu
ffgeUqAUfY3OmiXcdDnGpezCmxTnKTIBbxqiYu941VotUMM7IDk9Wan9tlhGqrQyAhP3vCfnzq7U
GOyhueH4/RjDpFMrWuijRYwVpdgUZdACqIgke739qMK8c67UOmXsdNkDklloAQr5puy8aQCYGfF/
Dmo1V5rfjJr7xcn31pMR+S88c9nsuoVgWWQnUsntUVA2tHDMdG52rLTy+fToVe7BA7a1igYI4I5m
BlW7iKJnWQukg05us23JfbvRFrp5sznzSleVsnK/Kb6ZSfNU2Rhw0yABeLAMQdTccKrfOU02UC9B
NbUaUbWhpKEmJT1T3E0axDPVeSCBsLdaIeSKIxETN+eMRCCOuFnL/UWps7CxZhFdfbPN1yXPOSHw
zSkn38DWsFCu/dZSBSBi0MBgRxV4eBr/iAm41H3w5oODn1KVR5sZcHm4/ZwcqcWbbDs7wOmzeAwB
jUsplv4Nnlq5KbM5hwMEi9I/RNQ+RAanQscXNWNi3shR8BOa8NJ46iaEY1hK0kVPk8ZcW6pnrAuG
ngVFIujCJ/r3+JxfEBiJMJlkIb/iSdaShoIdFGSvhUQB3P3JH5yLnXqhfKTCxabjV9k+qPoYsc3H
cuDodtw8d7W5rCmdXTURABrHse8wLsuB1jpTjhZWLqvyxAuEgC90xU6Kjy2TZ090W++hhdgxQpB1
1rYAeyEeWLdz+WFBZ3UbT2sX8zlDCpAnke8kswgLjr0RwawUYlk1/ZC1L7AxF1FlfMUTNVcPKMGJ
bCsRKo8bXUyVwR7dhzgDDUCmcVy5EKLmdGGZUYIyKa8EB5u9PtMy3dXG/X/VPeaJ4mqFO+UXzUhz
8DmNa/e+lSEt2B4vl4OpdRrZrwOo6GemgC37rz/2PlMnowgS2ZX8zl2H+nVBG0Lm8R+4ZetqOC2X
B10u4gSNPeR0VRXhmL+Vrwy+2BF8xj0pzdxqKMFyRCfQy05hjUg8JMJSQcME6MycvFFXvSrZdumU
gKBUcpZmfVjC3Dfpd2DnIK8wEpSgeKpld7/miGn03ANUAeefpNfsTuOQAvSSdO51oo7Vqfo20FDy
vYnWabQpDTxtlrtGx1/4pN9aUff4rBBk8ADlnA06WRQp7tclVzX88I38sVpJQxfPCIbhsdG0URvJ
pGdHlFc8xSn55mVrgJ28/YrcpERRKCmQ5+uFRoLChinNs1XYXBqrecc5b6SN1b++26vf6P12hJjD
K8Xuc1yiXZ97Hcu9W4M2DLpujYpW3TVNoqBJZ1FjR3BuEHbWYV296tkFFgB0yWWNQBiqbxxQLe3Q
082vRkrxTJb9Kjy1JXT62RlMp45u/KM0VGu5h4O30OY8wdOiUVJQ77oNQiCEiUQ2Q5wNNnmtukjr
eS+kfG9PDT9RxpeHtFKgbH3UCplcn6SixgYuoJrDn1R9/ebGDgIf3oSDSaRLhWuBKceCnZp3XBx2
V4RC9GUcve1K9Vx1kbGm6yJj3aV4kTbxpmzuT7yAgvFFODY3Nx6gDjE9ND0eggz9wTP7OZ84Vu6c
/83A+d/zF6ewlgh0YsX5127kLSjUxRDHDufQHXN/IqQjsBmuPhyqYddv9HzO3D4GcT2aBvtbUmRK
yS1Y+xfZkUXD5k+9XdFqFsDzC8PWchW+KWY3WqSIOtpggpOjqq9vu/bpJOFf0FMB2fGi1Rx9yWsQ
0WNkT6DD6W9to5ucK1sYcYMaXQZ4zB0V4zPwVSpWvSSQPI+T8xtM9MYQBuxh/NBWKQNlOyqL7iuQ
QeDmkcucjJDhMEXl4npWoMNu6WLB1He0LctoU5cWsNxB37Bb6fWNNVUnb+ylmj3AYkrBMF870pvh
VerduXFJYTmU00JPJ/jNqofVdcqzyVWY/e8fdGiqkcDHgQskCq3+EYB/1dttkXhUZx5vgxQfEB8X
Cv4ngc+81orU9dFl21pOavSehW6dlGyyUYkbd1QaU3hSbarv4CYlvK2z414RN2hLM6Tf40ILs0he
go6ICwMritfQIZtKDNgw2b5aRMtfsVxjUM7HqaQ1bKlIfbary32cfCUVPKeKzdH99kE7Ra3PAcXr
6f+jVzZi6uQ+O6LFN3kuavZ/NJ8KFwYSfYuSlO0AK0S5CgCib+joBShLxTYJwVxUWp3Bo5jGmQ5k
T9EEL9s3Bt2R5A+A9yE5upVJbGVB312DhARDwBxEs36h6aierfifR5bY/SKw6AXLnCrBgg/e1dN5
0FeEfrSLhfhXzCp0kmN3wnODvwKaQIcmpD+aHr0I2WXN3zMdTn/h6/MojPhLVFjBOKLEED4MHZoT
3EXgSUXDN6H0NsA5O2EcLJLNlB3OYT9S5bUWgsjteCVKalkUjQJgAzhyqNKNfik/TJCZRK6Qx4pL
Q9JRnkJ8BdZTwhdJA9Ijd1Pr5WvsCNDSk7vkee5lp1sk2iOAzorlkOTIyC6hF2Es03LVizePnsiL
azQyxtUJaVCjO74rRxa7SRIz7/D6vikxpYXoo0thso54w49VikCJI34juXN2WRZ71cMKQX1CE2PO
Q8f2Ih0cXkv85yJ5HoEbgwcRihOelK2JtrIt6zhibMiHc1FvQzDIR5UgQ5Hlmfui1oN42Zr3+ziu
B8TIVPQt3h4+Udux/s9vEwJ8gL4CARgZFWnr/5ecfFViwy4aqmECC75gtik/gWaf0F2FiiiYUVtg
t9dUCI1LYbgfp4kf7cwlN4rkbOsp9i7E8Dv4BTD8Wz78tiL0zXB3cEUDQJ4fDMB30jIJBE4v7Da5
/ym0iZWv/acP7eb3QmKQVV6nsFHef3JKYK3PMidhQmrOeKeq/50QY78Zuw0LonMhxhnSfERu4y0l
sU5TNkW+Dbb4wg4C2CmyuDJwhH9GAYSXNQ03vyH0rDe2l6gYg7rmcjAoE2Y3FLUTbmBSA3vjJ5AE
1Yb2ToqxvCL3D+uJsSIA0hzzXwPr77gZBOkrJWyVwwWwlq1JFK7i/hvONQrP57kY/lxvUbZE1OOi
Zb6o+tPZNfGW7x6DjoK3kP6x3Ut3cryp9f+IyhSt5Sd5NReRCdE2oSiS8QSnAAuahdlxIXTRPny/
BuySnsYWf9DqFzWX26M7w60JMe4KCZT4VY+f5UvWpmlV+vgtXE8FppoXwTZez0JQCf2tgupzt8Pf
n88keU0dFJ4NOiTZdpeFa0FclchFwuL9rGLZMZ89+3qKNIhyrUmNiAVX5k/W6eo3OwFu9Icu9CZd
zKfACpVv14UuR+qTCLmz8U9OIbDT3jWXgYgkzdpQ/jRdnJYASg1RP7cKpXf7l23U5B+Mpgl/s6Bm
nwVtIof6zq4cJO9iDqozxNqXBadb9KMI32O0j0HYHUjlhRGoRPEykY2WBATVMZEc/oWn7f8gUqHW
SlWRsYOm3ofk+qmCjWEtdtOsFsjVjdUze5iVoBwXQ/tu9YlsP9KguBMhsmH5N+vfBZm+/uVJmuhH
HwvzX9aDKT08Qmgz43dGe88v0gicjXgzoUky8HoWc5mRN76a+VAt1dbWKb4tIzvNpn5wDVl8HxYj
TbKSUAit0DKHf2WcV0k30+hopmTMTW4awFBiNDr6m4ktZV7tWpoMFvFM3CEwxnQOB4k/u/FeHYGo
ASK4YjDwfpxrzT8w63waysxrdOtuhzgxnC6ITFn66PYF47eMELRgGLRBcrXfMLyNA+3JEKESHDmm
jmV4YWG7nu0YxsgxOxBHHFAUCUgWn61fw8oV6zqcsC+gQqos9crirougXLBEpyAMLzOZioAZ5r01
o437r1GdmA3miCCvpZ7OyySVn5knhAgqpC4IpO28WcYqZpaWeFC23PiOqh32qQQnRggRzRUTEv0w
ik7wLLhD5DkkPoY5j/rrihPgWHSlyMEqq8TuRaqGy35zZcU8hFwrM6sN8Och3q09r8VGYq9VrnL6
izrILn9OZ/FSfX+KHhtyC5AcHnKKMslXn6mGivST9Oe8QZ0/kKT8R7+COiJUW9mqS6hidXPENub0
W2F/zahQXNTKt+PQN8pcEq0PJPCmZQ/IeFOb+yLxPviIG1tVa3w2jnZRBbYZW8UY2NAxjSVDiS6Q
WBVEkLhWkq1T23xPYO7u540GoMQBGNqdNg5BcyUJ8eZwaGQaZUPbxu6Q8k3iOM+R3KgbYUqLktSe
n3xEkXhV8kxGVbTiYDTrGbmi4/ne8j54BTTWFhu2gq6/0yT698N+3gTm19nkqCaVklyGXKdlA9xL
ZK7M1LrRGl1Q/fTzzHWukNW/WZQL9+Qe0OwTRP7xDxxLiqHprdQoTg8yV3IxZAo4popGCEJb4fFy
Cut6qEBJN5HNTGpgPtWnx/8BFKcwTdha6k5qDRMQz+ZYoIwaKrFrppzKegMFkzgMbW7Ul/EmYtyW
isZEycCfl7JgM/xiPMSx22K6tTdfoRUdhbPd/hV6AXKTnaOEj83ojsTSdTI3jkWtVF63sgfZBplO
tNlHzn3JP7kQxDYiYSgYt/E3hGGu4Vp8wuu/1B9d6R10QHFMxBTTtRV32NeQzF/AnmI7brCEawgI
lMLjbJorWlfWDGSxTwkKF5gf1XEz11pNMCy4XqQS3tLzGzCEtuDlR9ImKME7lNnKFsyZ7+5d3B0G
1vOT7ePlYgr7oSMcS3h6Xuu0yVkuO/CZElMmwS0YfBXiDHzQVDuXu3GMQzye15yvXLPujbyHu6WK
O+op4DL7fvPO+HZ9Ud5GzETgRPTlFg1svEqw0HJRiZ5Ass7R21bVg04q4pr2sshrOCIQU2cQEF5G
YuN8ikudFZNgObjCoY9tKyV9ozowzt1l5EUoatyR7Ea5bYlbtUl2UPRu8iubyIHN7J4WjGFvZurB
6z1Qko+WNVSX628ObH86kKj76U9kLPzP7lynoXmQx18JiXqMx8eWg1M1Sh0B0eUOMP5cW7wtcpH8
LEetX2CwvuTwk+vjxhEt1VP9I8NadA2CHPnySitgnwqN4p9dyaOAUOoh+INHRc1oV8F9803n/zmz
jAmn9G5SQ/TAcZh35PgSSRYqQaeMKjfscRDbH+Gi/Emz4btR8KpqtmeFAxCeTzObhsO+GbXFRuXZ
GY7vGU/s1JNDBt9dF3TR1bKVibMMTAFUeE/KZ9mXcfWG7hMNh3EhwrCuV8i5fs3IdcJKuDYzAw6O
4Rkr0d+UN3xOWu/jLTBgd7SYBFc+zjZZZqhd95UDZe4lgnZrXZDqWGHieqsdOJ11M6nZM1WhDzmF
4FpovgZNnoG+NM/nm6t6adIU+MZYob3DNsTLhdxetTNa2nbcTEbhhw67tsrlLLZfrikJJq4kjR4W
a7rHkYr7j4KFr9QE01p/6d6Otp9SkIjIW0Lhk4yCY8+C4ySNDXcq6hItI+UZYrcmshkfFnu4MsKN
lm4vimaErElSiD7mXD+aDruMq9ocUP6HvQUslhHvrwF/nt17zkGRtfUC/VFnz3gFXntC/kO+iNGc
uPIqmTKJ0EYVkmPEyp7T6DIE/C901eJsbTkvnF8KU+h34BgW9OwjboYHLKtrPEb+6P5AaH6pHXGu
9G/z6am/gSsz2ts27ddPzVbi05viO47JHA3wl6OceMOJhUJamgsyGAeHWJdflsc833qFrq+6AJBG
ZbJyAyzOPMMfxJsCsrNDT/8W4emkSZ5qg71BKUgwLcX2Vhw5bzxZfiEICQfK89NifAUKdiNOtRV6
KHsYcTyUFDAYncP426MrY0UB6BDuq7KNM7PjAYh10g6iSRspxHxpmoLLSDf5w1g8OAGLWfagpj+S
Yl34T2mvlHbbVP2ZjnNvwNZFRHObbVod+dji9ueAvGncZGyxFIzuebLctr+oHHv4S7ssgHZuogFp
fZsvtT1xMqA4ttHuSUcQ+H6Ekb/BAigbsyZyWPRO+4zks0J7Nf6CyzhliRXFM61Qy+lMkmjHJbcg
zVkQbPzD+Fhufsbkc5EnvU94m3hOjcE9zg7e7Lg5ReVj17+U+LjDeKdatm2jBpU6IFUD9OnZOyhs
f1vFelqLeqxilDMWMhQB9iPfBK/vQnlueBW2sRdI4EgLzpa9wDJtY2OymLOGciHrvfnPR/8ZPs6c
NzK/BkXQZXNXNVHxdGEr3F9GyR0BEkEzoPQcoMDh8s1hCxxuOJ/GOOHXUvg6ZdmvaclBokNWSYtU
lw0Xy++Yr7CH5rlObxpKxCxjxEeShNd/CgyezZkm6lhb942Go99FTiQyEK6pRJeHudyZP9+BCX9R
CcvH2LrvbYATM8Dfbdt/le1xjaq+XLeeZkPgKz5KbivcbZsv3HDCBmxb0jnXH3PvIdym17/EgXF6
fEw/ze+TtQUNQ6HHQtI5Tg2baioqX015kuE+MraI0f5OZyCmg5z4khWMapovbyyXpR9JDZRzc+8y
a2bH6/8AwXtwhq6XlN1mUP3N0iwLLu3h42KMKYZMMOpjjCETfeIV1hAiaNKFLSoy35NLbR/RJ/pr
dmWs+s65fGt9nhmZPutmFFJI/C9Ob8WZSQvB3YAP6VX/j3mOY/Wj5SMGerJxQdR72zD/Qx6rYfT+
ZRu0fq2ioGODDBhfqjoxmIWj4j35DKEXaKKwEQLJfTfhCnPnilIakUZ18xNZRpY3gmnu+FvoXPwS
4Z+hmbyRtr8Wi9fqBm4efBGE21RUCVeyJzdgzQRsKUTydN2Zb/Xp2q+yJhb8lWOPrcKCtZVCmxVs
ciX70Xpf5ZRnOF+tDk8lJztxONkzw+zeFh1uzl9hU8hDNXhHw7E7MHuHAwYSq3K91aJSsWaZyeR0
JIcNXUpgmqLR7pNicQ5ebFYRK0qNljMExYfSCYhzCmjKIqZfLV2eeT/BexXhD8Q9rO+W5bIQtkii
7xmuMfwcvCmjbCW1kh3lCSiOqE38nwjgSTq1CSr178Sx4L/ZIGMd7G4bxzvnWXHEYWD0pNLKsJ47
ATP+E5vefrd5ThARph/VtzoREbtC2ayFz5Qn8QYfVqugj47EVCwvgBAFNOBmkM+XyJhOSii+myBe
jMjedQueQ9kisr/OlD1YL9UzL0gh5TTi/BGpA58iwKne/dnjgGUrBgyErXjf15fFOTFYa2dXk769
MLj32IIv9/hdsGT6UZNEFCHGlch93bhpI7amMWIEw4AegPaT9z/FveHw/+DkyJDgRVtYJwkBBmsW
LEoso2tPo7sGsHU+Szm/5RJHCNyG3UMdIm6HLuMkyjh2D2m0eiDfsfGVqP0u/gLU2qp/OLJwNf0w
pQoD5uuDM6Ubru9AnfEb4OtNMQzniWmk+9ZQU1eOqeUoVVpDqChLsBE/0HZvROlhcoC9wmxTRfhG
9Xg+vrOC561Ek/Vz2QTj6SQE1K+0Uo8ji5LsxD8EbxpKoEaFf/GxM2hTlBvGF3OrfEaELPeBAE69
GOo1faZH8ZiNfqnUnDpWjW7uEmDA/y+9l/tWfSn1M4SWG+OhacHRyPod+lRZwrx6uIzzpiu8Wx6a
G8CJqKJKH2D+rgSwNuMUufB623uN2xwUFW92d8jxiWwP72U4bPEwMk45BcYDp2r16WE/t61YRKCg
cbshnpibxKEN4ICdje3t/uRDL9YNFltyNeGdp/LeJcf54kKnr867qtNSKCMIMGZHKqmNwzJC35KX
If6m19N+X3YHUL0eXLSOH7zMbENum49+uX7SBWFw+t6D7orMUooOsbTwirIl6OK0iPnfDgYxVaqD
WikUPSPLdmsSuPIlG5VNU7ztfCfC7SE+5Sd57h6Fi+xhjqgCVlYl2RtXeVg8C1CT9/387ZFF6HPb
+wiA9Jbavvjy2t8eTptw8sgMJSe0Y4jVPDHLiIrqKThKiEO0n898IY8JNGgfJsMFDvV0zr34Vh4q
oO/qchQcfIKzuoJ+1ujsmlA3yEf3USebOKWuWX8T7hh4HwQQbEVUi+nrQYmjcMvRTpDMkQNOUWu/
3tgvq6jVTW0VOw4+Q2TanSTy2MRjJhQjNTmO/Ozxum/OjUoyciE+lRX7PL1HcZoVL7+O7cO/MI07
ows7ammWsa6rUTluhFKeQqrSs1Oq7iS7EeBs0IvSIPs8ebDc258Y80mO+TdLbfFYuFMjg2KfJjSH
Z1a5Xzkj8iUskm7OmygfZBRQfGf9m/DGTEBCyXNMraDmWLVkGDQOr8mSDxrvgz9Q68rxSaiaLnvG
BLDgEb5+lWmhGJENI5ANHNWavAg805ZV3hG2DQ11lQnkDNPsBHQtWJvVGrNIaQyom7DWGYMVjjVG
OG8d+Q1wbsvnAa6fsnwrKpM+RLzD8L8JL2ojPWzmVmgjTeQdcCBz3f5IDsKUSAkRs5l0lfaQI1ly
FxCYdhm/cfuA65dpTLzxdivdQohghoqTDkJmW77EHI2sef8IpZMoC2QOUFugeVwtgEtCV7kVFVsD
HkeHzgDyoAC8Omr6bK+02Tn96g5Qixzda1kV3DjqC2SHA1XpHBg1BUZR2ibWMUwws5jQ9gzf7H9q
mjRwDBL7cnSQpN722sHMYi4eLe0o0rFbFk/SwTXlo5zPmqMrB+d2jsbBHzF6onO1uu02W2fCEynE
ncnxBatVivEpVM3khv1Rh/3XViiQctiClJxrtuCgXR3/k6V4XWqMWawdXMn0AjARc7LS+JE2zRt0
nUzv2x+IBDSVY99EbFtq+JXeYBwgcsEiRz9YFuPKPHwQNGdWDh8iMQqpU0fJ3as3K6BFIGTjkae+
aR8AVcZutFnXGWwR80Kq5fAHQmQDTRwCEhJnD2uYbOGfit6wl5ajh2M+jhs2lnwNt4LUUkvy3HDH
itq0rdBoOeObcwwA96KCNfIkMRLikJkc+db7UuwgB2AtCgTX9MuIeMeUsDBDfSRkje9eOEk9QUnB
Ba0+mJm1gDIzLKAK2YIRJaSunF4GjDnS2NtyVwdGTP6DxZVaEyjY2uNV1Ar6cdTAYde6jXEM4jSm
/eclU20rGgw2+yD9TeQS1s9fRaLwXwg7fdyqI/uMc0A2m99aRIUV0Cwtya+yP9QEYKOW1K8CuiLM
KNH6M/bSpIVGXf0M9ZLeUeCE7GgLLVbrMsBxbGbxOPJdw/84lWCGX6CRWNCgyI5P0Dwz3s3lVc28
6AGUMm9Y3oK1vCTN6fuxQJB3S6Oq9jex9Ha0GsALEqbqLc+YURktq13j2+PZ2wRJ/eogZpph9S8C
xVxCaSkKCE8ZHpOEScS21qV6frGpCcmtlsawv18X8dRvJNuflw05/POecy+A1uNxAeDsSkZGAQjo
Gzqpn0Q5JYig12q4hj+oVK6ZbC8rMHBFFc5X8WA9+Dk6wemIaTpNMkvlNsIsKXdttPFdYfIdD5jL
N7Xm45E6a8HnrR1BZZFydcwV52Mw0chOKYXByRqjPfNxEFlYvZNePCA4CykoxYpdv2NXUyrTWGbR
4Meo9NX4FEB+4qgCbTSBxyden61vVIAHSvKrgFs7bsv/Uz3v+CA6TsJ+UnieE1Y2J3xucMrs9xlz
EMbZ8mgsRQjVU2UqEFTEWZibHDyJsrF0NLVHBVSJT+jKuMoax0SP0NRWRdKLFtNXIS0UDc3uUuRX
aSTwrxNuP3KyPXEIcgfIFO764vwrfY7M3EdkycXi8hvyfQee+4LKhud2v8GaPX6+gr3rscLagHqX
/0mD/wM6UuCDRj8Nn1wFzJ6JTHkIOqjVUjlqvYB1nmZRUvbEmi9O6xrKtTpoSECD2JQJ/hy6R93Q
1QuQeZwFmaS3VRnc4eB4shi1MQHCjvWcVzYWTZpMTtRdVA9qQxy0H5I1CBKhEP2m/MueGSb44XdU
EvT5D/uqs2ye+2KdXVfT3YD+zuBDt8XeGRHoEC1yLgj8UELjFGAfDn06AkRPD7tfUteNV/EoRqx+
rt4jCfcbhvvrr4KK9BE4YDcdWVTKqsBzZ6WkfFEyIW2Upb5MhND1blF4peDrbZvHQtUfrxW/fZBn
Ob1yLV+XNja+acg8k7gtrFOKuR0EAimVwFxIy3+5yvE3r+Zxb28xJZfaIFsNpptzHbl4qRTPGivC
6+/eZXjP8C/FG1xH9VbIYXTAm07D50JKJ/R3eOYn2upSbRYyU/yv71kkxj9SVn5CvCunBc90d06K
VVxqpsufORVkt1E9uv2YCQxFeMSPg26N5+7gmZFuynduoHVoJf7FzDUaExNrR7siv4wpmaiLC8Iz
WhSHbzplIv31+HoYxMB31C+JQulcxgya+4aCT6aFHNsbZaigQKauLKDJMsbDq1r3XPTUI03Fd7GI
FP+p7vpwgZrADAvBbbOidI47kDAPWmVXVvmJzEBayb8hu31QTAE2+iPaDgJuDWjndKS2ibwwqnoT
djowVlE5oNzSAlE6T4fGTAAlF6/Ks0utTk0s8Gj/rk0w1zqmEG4qAbA2z8RcrBs9lBSYy8UY96Eh
EGgXhBJ/1yGbpnAAiLKYMNooFwe3bHmcFJ5GghklEDOl3e4dfEgZEsjfw4OfsDy0FpcoaySnS+mV
sO6vqV91h2NO9nDzL6u8tjBGTIQ3yf8/PuRbExIj3jaX5R7Bmi21WUgYW0xJqmXz45UpUSCMCQ5g
+Jb9Fd+JdCSkLXzggZRpvA4qZOqjbSuYnhiNa9+aRi4q3MKvNqNqnVkgpuzTxXRPmo+TH6epvUKt
kvPiO8FqxrxZgGBSXlezIwAqDcC7wMNe9hNczz3U9+OsCcPCSVFMlYK2CBIYfcGnDwSq4jZNOuFA
+QHr6WSDjvPSomYBbU1f5vF6vMY4OkIeXVYvLT6luO3KIiMUWJATo8HMV9JjIbfK0rG/9rTV3MuF
IwXupfugZpgQ0G/reOy1VYNw6EZFWHuYlmqiKHPr6A6FexYH1JLDOLb75uSfWM63DybEnZSZgsV2
nlHUVjAJrPlBVbW1yy48Hjw7039urAm2Jyvi/oSB+qh93z7XPn645eZH7xx9Nz61QZMMYNqwT7h5
KWi4tA5XjUafuHLx87EKqqUgdh4KHpXuJKvYmnaJEPqCWXIzFN5m9OSYywfjywbg2tCIKaDuqHFd
OwO3HcPWFw5RZrK2P5X8Jo6emTulgrewuYLM+0crypgHLmUehS3Fl2hGlGhYgdfoAQ7lBdzOAvpg
+ZuqypFyCIAEaggfq3EUow1/IBGSInvL0yRSTdt2LLILOOf3cN+dlhN6sE51drcOFfheTSHsX3UW
hpx0HqqHu+zgkmX1bR5C2FeLN2rMRmOZvYVanz2JuoZ7k7SyJIuDup3OApVNikhTmSUTqkPmpUkn
adio5WHF7lzrEpH5KJcOJrOBaqrVZ6V93zv3M+MREJXh7pkuONEDeSq5geiKi4VCNfBdGXV/BEFr
dAiyvGUoEELf9HANL9KFAAXBE3obMK3ETROTuILN/FXBZg5mXjWoibBjlE/l3TRk6F8TLhsMvtMe
eD6iM0uI4SKNfoqIDwBEyoKcRrfy1nQBCUCjYPbe2fQuA3QRP2pGITdLv64UT4C8EO/Xndu38NrB
mHggVS7ZulrxUttNWVEZqaM0scdBnUtmor56gMyHnLDmiylsgrNEzQndnePZ6mmazttdzKNvtuAe
YCIbSTvLHG7hsIhSapS6FD2/sZkGDwW1dSHayGA6qPXlRUqFGiGi7uGLeQEGZxbTuyNjRCdSLpCt
7QKuxhm2woqBqqKAYS/0vXxrKjQ510LxZHmZaRA/iiDu6o32Ro9Sk/j9dZchwPZw1JYGjs/bNp0A
nzGeS6eMhHqdTS4tOxW9AT5aUmrZzD9pxWIBJUUGG28KcDqAZSNF5uMHk09/Ow7+zMsLTvqL4kmh
DseIrqYBlNLXou5U5aZkbQEDH5SJHnRQA5m4f3kIQ05WaiZVmpcGz5B/+KpoqjCI/hsuMPYx1gnO
TGApC6HGYaRXb56VZ3Q3iY5/VB8S7M+L2WV+xzWaXBHVYM+xq+6W+vDSeqq9EHktNgI/vmvKAHu9
gop3OMADC8ys2693c9Ocrx61xWKnvCBdyzTCMZKqGD0dGCSHR9MtD9fUgI20klBlsWEKeRe9F9eL
CZWU6dvXOnzwhHpq94+7lH3gafXMyiMdE6vzvhJD41igEQPB9WAsZKpVULB4mzJ2mVUIA3+7RWNP
rhY6W8tKMAitemylQIDYF+oxDulW4yBSGTZoaBT/EDS9JjWAC+Fnrmjj07bBjIzvKz1FXn7BU9EM
zdNU1nR59kLhK8xfj9FYfLVlbOI7++0UOP95BNBznvZbMlYUtFbxE08uc/JhijJvIgfrpMEoUAhG
grPk7X3mWbiA21+f5Y89ZooK04MsfuEB4yQktQesyPtnukSvMYOOC2rcJynFaU0sRgSx3Kb+Q6VL
YFRklaie57vw1CU/iAXey8Ki5F5UIG3GOBUu1mruTwdbZ1IdGbUF/bLgdXhEHXysUMeLjnDJa/r3
40lL4DXRJ7gy4jbmRRqJOqWpI0/HzryTWZjsMUHEY36ldkszFsP+zBVWRYgT5FvOTpaII+Jek5ea
IpIxECVNpQWkgZ1JGUeC80heUAgaw6SPIFVK8qGzUp/Sty40kMQwX3w379IC8y+7vVO3dduS+ywm
V5MYDtzBxpYHUuu/5Hf1rO1s/i7dyXX8aR9upGDyjJ/PLXKJfSkkzy68CU4m1X7wiSSYkFTNwxNo
ADuBZtoMiKWx86Grf/oVBI/JcKehGtp2+5TvrEzb4zBpTG5gTCuRjdN6IgkOp0oy83q0uIKEwNEM
44Urv7rOtchlijqB050fmTTna96jnVtixBdf6Zfed1YiyE0bXYF8xniIKLLM1/olKn5HFhlvQWek
0wHlUjTIOrVo2MQnFvdHOrdcK8mBiNPrCcqc1F9946u88fASsZj1sgzdgd8BGc4SqkRiy5Z3sCsp
I4s1TiygbWWUS4l43/AG6Oibcd5EqR2No6oZaeeVbXFAtC8UVLTcgGqXRKAX6aC+hvqK8V/kPG1u
3S7XwYw58CDd55TrFxz8vpEVNofrnvnazptvx6NYBNN6hi1u12hF3n/XO8vvZUvUd7bhmJasPLSM
kJlTu08KY1KGXIo6iOt8lGd8h4B+6dV/unWIrh6Fw3yF1517uQ+uuXNuEwku4knKYF2lmCm9xqAz
DVFa1fcjqB3fRGHRU+BPWBMqXeIBnbfRBB8UZa0gQxQriX+6JDRdfO4BjHYwSQ9ILyq/VEMa/+oM
JhCLiR32yEbeRwV7UyDeb1OlDwZF9nVHpDBi9CX8ZdA9QxIC0hpHA+itMecs+jcU0eOLBHKRzpKJ
Stb4AyexaHpa+lOm5h5sKGVNjEzIVSlfZlgH4NWV4rS0jtBtOpqUiN56eeg7KH+hQ06bvb5IQpSQ
iw8dSn43U/ys7R/LzhMtHuOW1hCpUyBccuAMRyGGaKfa88q5pB2w3zzWUOEZgjt+AaX8Fr99gNmg
SjXeAuwz/pz/LhE3c9CfaxBXF3bCOcl6LkNyWyPbonVNDSrDZtBRdRuBodNBFk3G4APiC1b/3xMN
+rbSfODYpqbyxGD3eMreTMWuIJdohurTJLXNAgWdM2QPSsTKGrgjGn1ez7S4qdeTIbBqf75OZLpj
fJSLzsM2VAIsMsYP5h+4Qiiq0eWGL9KyIUDdsKZY8xrPJm/0YMQPopMLjVcIuafgLfhpbMHOqZk5
wqzGFZBnSrCl6kA27JK43dIzIfENnnFGWqEk7TAH48urC3vBacPk7LQVtqNAyd+FhxMVt0Dgx6q8
XXuIkoHueUB5WnOLxr2qIsKoGLaizsx/2nstmpoUacv4T/IsZ+MKEwVYNkJDEeE4/EOmUpsJcxQf
u0yLwOSB6iUH1gW9qMHSnh4pCE6LTRacCrQsgyAY2TydOc/rS9dTwLDKF3puNA3Vy6EsZVnJ08T6
qn3WsSD2EdYr4T0HNVWNhkcAOGxnD3HUZQERnnP9LYWn1LzhqTVsb+G3rujGDOXcko4AbsJTgvHu
6evqdHu/iKlJwpZq1mqPkEa6HOKLgVaRoBW8Q+uKCJG90mh4mUHiqfzZNp9HGudYHBYxM3g17yur
LiVhTYe+bRofsuB9lF3NtUJC9zvtsD7y2E/V2aAMPlHiM/0A2hBbosPWGue9iPMXYoAt0ktdRvQk
mGamW5r18wbWT8ChHtM64Gc4MEuYelEk/LFXuKxL4Q8G2ljukAt4YFb6alWmWJLbrGyR8ZLVRuwp
56VJ9xKj6Eh4wlLHfoHBV7yYNDySwNjDzRC2g8j39dfYpVwa0bxXL4u96BAwTYPx3cUBY0nzkSRo
y5yGD6uTSV6SUU6lfVWD5FkDBr7XDw9AmsvvhQQi5hxDMe2EybDyW4lMk0VpOcgyF0KLWcHpRmYX
9l4BocwVj49ZXSl55AC3COvXL8lfJ3Gn0PZJWebQQrvIurmLQ9De75euNjSPyxg8BLnQFVKjilBV
zRTIFfLEbUf+V6PASn+NHx9hatgqStev4PI+Osn8Qz1RxImQUTXyXEh9Gj0npgDXSO9Ya/spUg9u
2Gaer2roClvNLfWddUT3fDV1w6lEWoyl9GI4ZDBiYDqwYemKQlJ0XHwOOf4yOXMFx3B3xRgpPRty
mhFB4HaS663nPlpcxUdig6mrW+37Kg9EIeMo2IVzZwOiaAVafJnZTU2onZQ+DY+GvwfvQhtYNEfY
N4sFdliz7Hx3speqEtCN93ntarYGc5CM1hCmP9TvOvkmtFJ2gSAYeWGqkojo8FTtzfx+GsWyCHtk
xe5YLdphd1eFfPeHbjIVH+gGF2OmDo0bll4MQ1GzXaD0chFJAx/Np1vfjTdcYToJcycqeGL8auHi
2guJRQqBMFTSM7+qX9RJ2rjX+2GWrWhwqEYfB4cLkbiSl/9EM7O4KqSgD82DkuYNoFI+JEq4zMp2
XdfAZQtcm7sWgSD3ZBCRtEMJlJ3dO/jO+wCs6Qto1k7sZor5WFB6ulLsPXXokvKUlR+WyD8GAnH+
eaMAkwC4AXEvl0pXUBNEy5KZKE68vNHpxCKHDo0ee1DY1upomTnrxkXxxPLt2pIutBV8BMSjUyb1
9aog79NPOAagYigtn5C6VSIqjGJ/bXp30YwrzR1jkbmdLau5XPFwa1f4++sE8eYIbh7sL2wC+R9D
jscKWl3DYf64crFAHmEhSFn3G464kZ7cihfcPA7ZZ2oGtm++yyqNzcwi9mFIc+CXJbs0Rca+qmQ/
d/3mzIygIpkCLPoE5HcPQp8SJMqZjzRh+eZBmgUXPatJZ0FejwTG5GDVS36R1dDbUad/08m9G8uZ
Jfjb3Y6y+n4Ei9zdIheEG9EwrKfkxJhN/WITMi3bWWQ1aEAjwL80xF2IDTyz+AfrXg8nm752UVze
miLhwL/yyCe3zRLTLbtshqSnVd2j29OlpHz5QldXLzd7YIqO7F5xW3etEPAMMPZpuggmo7xNzaWL
+B0HV9eORLRTF3ycQbIrObKPl1K/aG6jzs99DiDGNX0D8rjz7Y4Qp5gQ0SI0eJPCPlj+Ezas+Xlt
FQMlGep+SkLoMuloaZHitzT0KGICYMtKWulsIUw5/R54zqTNdfg+FBIxeRcZUbtfk6aqX1TrSAvX
/fbIbo4A+qoQ5eBq0pjXx7F7TAKGXXzQkhhyBLwfHcsXUQxXppw/ckIUHMWH63ssM3Fv9oVoVu1z
MiTpnJWPYeBdzUsN32iFCU42M/dkJEVZpbYrpgQZt9yPh77DlYLsNP7idp12b1oxoLC+rS5ymeHo
Qo1jIbVqlPw95taSjectMimEGcYg42et3ojJWP33rOUKN2UbTXSeArBkrfA8LiknrzIVlzl5A90D
rcvouBDezwojxpOsGT7NsTqN4EM1REO2zpjUvcgvNlEXXAIlXVohBuHvybvxirUbmQ1kKjV2rrdw
72aY0RlJekFU1LXBHn1qNuT95rIopC35VC8TOEgzsHLkU93XTMi/VRsr1sNHbDcseQSVKwgs6aPu
PIvD+x3COLTxlQKWhN0ZOYafd3YXQ+cpU1vw4cHYvkO/yd6QH5pz/WS0viaff6VaHfqy+nHlnWTT
MS3asXs2hwjFFAnc9GyZkxi0anJdNWEOMplGKoEQM3/p3SLnAYTIVRhu2BpQdI0OlA8aWMS7zp+k
9ZYB1ipN6oqoLOP7N5uI2eLoXJUSPrypBFvDUbF0mmAIS7D9QKRyCinjljfACvUdEV3vK7D/bce3
5s8ZzCWaYkRn+1b96odPjK/jFzEpk55esSu4qs3SQiIB3lzmEQHYSfhoKUhZF9m4LAKYYkPpHP5k
JRRBzvfyAK0Stc+I/P/4WRqNKrNyjqL8mtbmWzm4ObxoOq2oa+FUGOuah6goZiNxKyMNeT3SDXBi
zGA3ZkoabLVFwvc4vou80rEYwOPDB1h6jy7L0EkC0GLPchHeuZ2s6rqAxWOprC1QL0XeILwHbdJu
4a3l2tQFqYZj8+RQj6JhgS1VN4xCxfs6U2wUUjVFLDJDvAimWigaVoLsPqn7ZnLt+VZ9z2q3mvhv
w3G3AxscbjaNsiE2WrMOjh2o9mTIHA/2ouRFCXDFfOH/BkaAzHmQiUn45VSwfVXo6PwGYlM/eaMG
OOnpzeQFUb94iTPwfmrTikFmUdsmu39eyeu0T3TEN10dgC3BdTUGI2pevZlbztxKbfnxrxhMKMpL
VSWvNvjGblzVYdxWRCNHqymTqMGMEkYYFyVSTTqcXzXG6Iki9+AcVDiZBXv/hVLJ2n+/EkeQMIMk
vQYn1N+9Mpm4H8K0CrPxjTIXkWOHdYWrkp625UhLSvsyek/Kiju/gcVObBBewMcmTyZtvo7uSXxm
QJK6liMpDT+buUePRW71DslmNOvMtyI0pYvcLiSBncw6JhfMfD/cQUxt79al/GDmLT0MviK54N03
/FS5n2swf9eusprUrPzeSJz2bOy0DpEsFTe9zL8ntOM8WfmGOPGZfwVzegp8Wfu7Dn3lYbdMYKtg
uJjyv4pPz6674R9hgKpheFLIdm35PaB4A6hca4WKW6cLmwP1HzCtOAnYNq2x1IXV7hM8Jy/Iyf+3
9Ibr+Zx3ofCENLgXYRPbdV1/NtXbeCmrjovOZw3amxeDsfzj9j2Ca+zRGKsPJOWs6FZsFmVOC6hh
Y8YNknVfEtgqYACSTqGDQBHgfHxq4X2X092EaBf2u5hAJ3idZ6D1Opjd2/jnSQR8RbDvElky/lXs
3X3UkJp38jLC+QcdHbvXQUA9uplJxc1RqwKz8ICctCaR6K5G93TdZB5Ab2stylKb4C69K69Ircfo
plmhfUGQkEa/NNvtFqzv8gSlvdaSikBQynBYwLTlkxw97PAiuFPyu0MZifQ6C5N0sz+2o1Qo24Y6
CL1T642AW9PPJbwIK2lapUbePZGK00VKu+m+ZI4124jQtM5R8dBwEd/K9gCXOMb+gFp9vDyo6i51
ArOP+YK7X4IHKqcERAEe6mbilNGTSgaBq1SuaexSaPEppzfxYTuzECs+Tz20DVvD/bssmWV3K434
64g7EkB03ST73dtGrW8ehaK6xQbYNxNvY7CienUhfXk3Q2ft0YdQeeXW2/aL1DxDVkAv76G6AkXc
wZ763Y/ERWzoKcaeP9zteb47rE6K/+isbqTPzst2TShjqJqCtJwWB2QC3Z0u4N4P1BEykIBBanCd
8TtNih3QETxY06VI3bq/sjJe8pjh4zQtx/9VRwKI1HXTbYHnAmnCtmJkYO0fVg78pd1peG6YN+nQ
13rbevOLCHYLM9mG7FaCv+xw8vZqf6lR0aMBw+E6lmr3FdahPCTEjkcSOz7gNCWE+M0rdvmVMzg/
sPHTiCtqND0BJ16h/zMFF2a0OvVQpskOk0kDyJ1c7UFK+TGOAsvFUZ1BOOKr92FtSVUS0en9DQM8
NfBmCBy6ahotKXTWkBufOfbfWeDSkp9PEZKdlC6TqYTykDt5Fxq6FO/1eE+GTqYMGkHwU5uVRkao
DorG2Qhi/4K/KaBjVc5Ckw5OgNV7wj282zk85/pFX2Omg7at8YvECJRDb5bKHyhMDWrqe0dletXv
Sq16Nh+4f6H2O5zEH6KfJx6jjwNrA9EgybJPr6fGO+caMaScRfCaMpHtPEBvp/K4uSFUv2NO0bYA
wUCCWHt7VvT6pEvalp/KG/7Tr9qkM9Rcz/S+6F61cnQoIdgXG2XUXW/KmT3/9qeVtQ4NtqNBVdWA
VfUuc7/+aEKlg279sVFhnUSO20Ji6PRLV0r6DyVpQnugi6JEnuoimtjj5R3TYMfYavAdJadOpE/5
kx/yWwYXoPvuvQn2rG+rMtueoIYMnfImD98px/H4lrexbnEkD7YzM5N7Von4bUEvKIj6dwow1myL
0/dyuW0GCpyJ1GWfLRasw4MgvbcUA5jS5oeOoIpdKkUYxfFeq8nvm7Xiwmf0rBdKR09eN9IrLzSy
tQIQkhsl+/KdSztDPwhKMgD+fqCmy+XprP0WY7IvWy03a9aI2wKQja0TwjtKhBd/E+NzEOrEuLfs
bXReVpn9T1rXmyxu8Xs38wmoK+dD2Iz+xc+fLjv2BHzNGXjaRSfDe9UqiEevKfluB3rBlDYctO6T
+wB9Ij/HXG085hfeMVU0U/WACE4LlCkfmUzFZJX3Mafp+AyQusMBwnxDc4hJbfuWMro3WhStoAUS
Ph8iDshFY8PFgj9X8KNSyBEA1It4Zc5AzUtYFJIlLQcnOERUUOBxKuTs/axLCtdvVSpTU53gAMAg
QeLFMpMHSuxLu5HNMGx+JfQhp8rT8SnNrLLe9L9Zb+g9G/lqseyU9uWranmtddTnY6JBTJN1cZha
CZBJ+7wTdNj/v4dCKH1HIm1ztxEIVnicom9KW2JkfTkNxOm9v0vov/V7udLaNhc6B6afKI3JJYhv
GdHCWeGN7W14HSdimVQH7YTGSZZRvntYR7BeD7H1zd7+TTHxXP9OuR3fsT5GBvOxXhKR/tXdZymj
ozmEhnP+N0GmhqV/5j2MXGre1AjwEldvzptY61oPxQR+x1spdqIBacS6aeYulGUmnaNv16ySeBs2
alLQ0eep2/xi8FwnjXPfekmMzeSOMaH3Qq7M/OXnQCdgKikTODLLjp0CQ5uwbNejXFGpvc8mEEYg
i3cYZm8NtRRqqfrAYdCReLsXlnVfUdsepgPq4dJqM1VcBlYxyKa9z/wGUuDEQcophF9+1fcho3KH
ROqy1laCExw8fgjCjGgDlY0kYAXCrTrJr3MURFJfsJ7XZ7TaTZ7YH/Ys+5bbm8bUypKpipyo1QS2
9HjiustiB1Nkfi5/Wv4XC+CQqGWbMd8urihG3WKLcyka8gJpz82jGkOOtsTAWOH/EYBSKmnA+ntq
DWgRaG0MrunmOn9SnstN9bo0QpnZLg/eBBbc9BPRMlR4pgptXaIUoeGVXgsc0f+u7pkFFzcXdVpR
Haby/OdwMAZuYD2DrjS05W2Ig6C0kCNAVKNQoGUAOacci+EPVkq9m44Adrr8vcJY2XZHRQU+iZJx
m9lSBsXyTPe6z6kFkzCLyYtcCkKHz5Pzi847VqVKchIXNHZXwvyBYneRtD9e/qcGa4nfGWfQQ2Rb
OLhrxD22bvIMMhD81G8+Ufe/IbW4+y9VdG1OYO3ieg4UNDAXsd9XywrAWLn4ScrwrvlPafS+PNWP
TIiFB9LxWtQqGI5YwkwPNnliZaK771Gvr+PLPm/YiXvHoXTMt0VuNE6tuof3mV3+wHWzrKSKgd1K
I/O+I/c/cB8CnXT8v34yyxG9EsoKIBMXC6pvUH2wxn7iUkv5rs0MwwtburBsabbkEphwR6p2u3Hh
ws82+0AS44YgaCusZ+lS5xf/lCxHryCfBgliNGKJPW9IK5rSkB0NB6M3D8pfGB3bUxewT7TMLAJa
FZ5qy0tPA3V/9VJ56Q6rxuDgTYAFY5UHNPSPYuxCqs4q2fnmRpS20mS3x5JJtxOEKCCiGMXlvpk6
FlIZatkRHgIc6j3JQeKJAOyqPaNqKNZu+r/Ioe+6Vd3LsR3Ml6MZD6u0FswbM73c1LzkNHXgZFrI
cLBhV2K+Nu6sSs8l6ZY/quNn48Dom5m3ZO15EKDoO7NTHk5BJquafXZVuFNthlxNdkgK9Q9jFI/v
3RliPn7wPMWIi5w0ZJmAOFxdk9JVK/WP8x5Jr+Hhv+Zca7cMD5U3L4kcgyjfaWAL6mKm9bfe3oqI
Q5d2c4tRxADRzwu8UeAoM0NYrHzklaT0+GRkrfFWN+00CdorMUQQ9JhK8OakJh2WJqE23Gx2TW1K
RYq6QahpK/mY/ExBjWiq1ig5X1Ro3k4btpBQ221NmkG8bXlS4+7ClGsZO71Ar6YMCUOs6aol9h+d
NyimkhImc2WnUvcADX9KFzl2U0Dby5v6+SwDgDhtjEzKEQlOUVfw/HM/PVNEyEV63+ci7EOl0MOR
pJ0OkvDTbxc8DSgP/8KRfeDwVJ2jMCmxn3OnJL6pkd3H+ysijj8iE7cQLP4puUDo0L46QuDZ1Xcy
Jrri1ZcbbUvfA+5I48r9haFXmfxG1mP6d2igeV8WLWImLBvYk18MSneKo55E0sUekDilDR6GkljM
HgZ+sOtAftM8U+f2bCYGnKaH/nFX/RLwjW8POLiLp32FX124/9PzkRhYyKihuWEdWutnHI0iG2A0
qaodWpR2akL6j/pQNI6/e+cS2/x1KeMOqZkAJeJi9mDThAIueSzdLTgiHzV3E8GbFEz51nLh2NOW
iAWUYoQC2BqMJBq5w7sPjcjYYVLTvK9ibO2Et0s3LN/Y+uSQ6RiWnoiioa5XUze11nbsQg3ygeb6
qgx+ZLrAw2o2yVs7vlCHnqVicPcnE0S8utfqNxmk0+n9iN8o4g9bhGXSHsN12i+7GbUXRr0wv8tV
83A8OnBSqXtEjFmqxgTlUEgQBm3z0cx31TzSY6+uVmCa+MREUBu1nRf8BOoZd1liWozZqkQphJ4u
NQgHENbicQZkCmCia1aX2FaLsDTBh/ShuLTmopMquW+lGvnFeqaKQ4UrMUN8LSoGdGvZ7GmdYaYR
+sQcse0xt3v5Rqw0ZcFuy6Wu78ZyFX+olI1yBTwEgZSQ50utNOXgBUyMisKI7b9GAHjEgLaSS1rv
X53+HcSr+VDIN8tbaXWYoumoCJpGJ1tGiCSFfPFxEKT2aafVHZcX+LI2wHzNoMXP3GKFBqctEeNt
996gOxRBLLSErTmlnVkTwE3sm8+A0HXt39BtVveBmgPeao/X/01rvBLrrM+ObwQ+RmPLzmzk3LCQ
1srQZc2udjHWv6WFo1ArqQVsI0ieviPD8aWIDMxDr+FaAs2rdNj4ANsc9N4UW38htOd5MSNx7fhh
qx0O07Arh1r6OiIaUT9RvigwgRuEqIEu1tOIOYKkHrXVcLGJ7cOcnXRMYLEHpCQnPvSWk4Uacn53
h/KAd+NoaxvwGEn9j44dd4EpTVHGqdG6iUnfFoGnddecjp78uGhZsHFBZu2XQiYjwdbyRBaVqDmq
T7NLLhYhbthX/RsQboBEHiOvD4rknFVFT8IIX2ZtrEFI8Dfc/fPk/vA9AVpOdsFrfk+MsxbpKpM3
Z8VXPAHwCOiKsepc1uwrMuGLQpaofZEQu0r8rtZqXX7OUntY9gB24m0qEX150WcxA1feGyho1o15
yzJlC7z9+nRcL8J5WrtGvGP4FzkIpXd1P6H+VfiqBFJt/2Q6yjiyyDycINtKQOogRhtwlIJpqHPE
h1sZJn+zDHxf1LDwTlwIWr1mfPxgBN0RZxOe5+VB0kpRJ5XONLMyp4Ms91vo79L55uHxvS+DHLM3
TXHK1ygMP5jkdONs4jWyPAVSzlvJAn4n+5rTv31+ktf5l7Kq1ym2yg7z1rMlUo2kRuvHCifrwlo4
+4caxyvzm9PRUog9FQGjE8n7uKRHa5P5SPi98bgqEGcjbzItJJhzfpLlniC2hkTHpQe9ik+kQ6bp
R0qLp7lbLdWcvxuEBYo91zcNuNf7Gcxr8r/5RufZQ6UntQS19nVfj9HLMVmj4P7aesUvtk15H8mS
MZbVYB0rNuMZOQzHpaO/Cf4VKpbwBy78EhOptZeTkVob26pcfKr0roMCUfaUcGDT2ukLl8mFSrDf
J74MXIO/GK2+K+bjq5SVj4LFgohLXmQ8CNlksiIMpWUD8LY/dj3UQCuYAoefh6+MDH/KTM7lOEXv
zGT2b7ZQBcVSfnxGcwEg2b5Rh5DwZyDEFMa+sA8MRfHUH1+72WPH/ihe88ZcIZwacQ+8Zgud+i63
V3pynyK+Z4n3xBtr7zVBHvPa231TpYbcXJ9ABqabmLvy6vY2/hanoMXDYdFbWxjqyBqfb3T5ByfH
H956A5eysaURIAuuRe+wFLDQwHEtySh2Y/9RIMGVLbiXtnhznYyIz/KIwxNUt6hWKyK0+uGkfkLy
GHC3rNZjhJyzd0wvVN1vMMzMcUqaed/Yq2SCDEN5s9zsKt+dt23iaqZgAu4l0olcZj2qKYrLy0fC
Bq2J2D0o3h3xOZYo0wDcC9bUdqrnSSy97aD6IQgNMJySvaYuX0hMpuTN773EZPtzSGEkQQKdZSo6
pvnRDST6IgZywrInVsNKziFNT1kbsICNCMSKArrHTRrqK+zAenFXud9E77v1GhB9CeoljQHyJEQC
VkIFihZXjweMAFBZW6Ipsob8/+eSLmLQbhuAsQ8YUZDodUn07M4BgHlnHSyt/bt38j3nI2zl/PHM
viFahiD8UvtlCO1fAHTX4LGBln4b6JDDBwVknZD98EaJMQTkaiqW8zavxV2By58SxvStIEV6Ck1Q
5Wy5eBQjirJkJgrfcEoJvdgaewr9jpPLu+3RRL5qHlc1VSZhtGrNCyY0OQT9BRRsnlFZ4oIGZ+Nd
p91x5H73cXqDqIAlalBodi6gXkNgaE0LqcGTLLKMiMt3EVoya+W427bqJExsezNbdd2kNb3yPV26
nLPY6UaofAFyJwY79oaAwLjwHcnWFLKF2q6MpTxTezSuJ6RmV+xZWHa16dEeZ8ftXqois6MALsXh
AiUxoKibExmB435y2dQ4qCPp5Ha7pmRtRGYPBWzu+TzS54Uyk7JX4icRocr11VRORBNQYPndyzbp
/mH7V/Ce3GTvI+ASO3uuMJGhl5MHoLiMIcf8kaMG6McSzQcKaJIMJ0BEt0jKcGF5D/5kidb/KNgS
lbKk4HZidsTQd0dRB64z1cV+MoNqsNw0YycWEqoswAjbXNRn7QW4/HDU4iaBFfEsyFWgBEmuq7At
ZUuJMO0pO1ZxweCyF81xZhw1dgitCSP6qcmwJjuAjgdvy8urr2ioj1gTarCMKugO+OK3jiYSTr6a
0QJ7GUu//0kZxyTTWvzPzog67ln2IxNrifnLFzbaES+Cj8CcZv7ryiH4iKGCzvKVSGx/MYNK7Ylc
9d8Ho9anf6E6/Fw3PGaYWwpjj0OcNdoJt/LPmCeLRGxttBe22SqyA4i0gEy1TStIb6/l017QMS6Q
+DXCvQWVtCymeCFiit8WqXyMt2T2Yz8U6uGLvmdaaEozI+cqQOFy6JVqamW7I8RtwZTV9wUtWLW/
zgWub1fpSXAj6FpLSCFAe78WOilcDCh88b6qMRdNyXCSA3IzXn7lPaTz93GFeqd3vywAvUS0U/Gj
tMROpITt5vdE1DJphMw1nj2LDGtDgXcQzlNliRSoIPa2tRxIQ6qUO/Nc8SoilftXeLzyudAoed9+
ytzt/HLPgH/PWxDSdYathbv1EbiNvByieoR624spvbAymkNAokJDA50cxpMxPi+4rOI/iF3rFSAw
xWxElGlj0znkv3J8+PXzJADnG1E4E13lNG9bphOzgny7c4EkzozrMoxy8JpzlhpO+6KuZ4o9fsXB
iHdhIxlm1JHO80H86IySMR1Cb1PGdG1CZRGfPfu+NI7aSVknJ6KzVjh4d69+gBRjoCShENHogQjP
gW3RNKY2FghnAE3/2y4qWHfusci6t2ZMb8P9LPm3KWnX1tosS8oZzkdCX6rzvfuovG9InTc+emuf
ndBnajulRcj/kSsk6osAV65T+FqLsy4H6esx1lAgDJe8BcqAtdIWiqfLDPPRZQsFTVN8qcrDz63i
sfaiV4n2fnKC9fwuvzhEIGHoe1Iruy67cz8EJdsahpKRBPe1MxpkSlvJ+re1CmWn/lUfuYclelS7
DffJ1VFqmb8u72lG/v3Y33Q7A2hjZlzjJpJDNiPa0ZZuXm9g4GITtYNAMl7NMZcBtGYdSHX736d/
yQ1TGac1M8hA0If82g27lapsLAEoMMgQ0rCsLhrM8Qgfobd6aUeqgbc5GZl74MVK2bO0rYsmGc10
SrrKm91y9lnP/LcEuDRVySiJnJgPmjQTZ7YGKSAH37NqGPPV6M6JNmguXqsJz7hfr5RbxGs6XWVU
7giKHDZtWyV/TaOYj7hX7h35b5EJI2Y3ukcx+QsZaf1stM9/pQgn18/F1IzrRXcjxDqqGORJc88J
7Uw1RZU4TQa6+spfnwmjcHUrXq0W4w0dnfp9KQ0v7Q0gL6mdqPKslS5QSIeExmU02P5NSvY6WyuR
uqc5RRfuGaESU3/gvxZB9CBUwLCFtbsMS32WlSkOh2FqGzaRRIwOl/N94xxEMgQgpv6YkbEhd1Xj
UtnuGSilq9k2+IbrV7DKzwr98d0VCHl/nr4KWfHKuu+AnpF5iZ26D98c9eQ5urRYx6QJxp583uGK
pw9PpLgh74wuze2RbNuMj/VpkeUgHGpKM2E8RRYNnr0uLqmG8knYU+Q3yoOOT4dEutjdFQmB92Lm
C0H5EFqF2LORdVdHJsW8P93nf7zagjt4G1YT1ZQhmFTAUQqdByAgVHQXUuf5Hh/Lqi8FxlETmnZp
RUHAHBsD2EGNgcwBSIp4AGWmqY1g4ElVgv2UZtk9taYbGLv1/G7oXfxAjyp+AQOTJba14W8/cGny
C5gVp2foezDBuRCkSBZfufqyBXVReM/+OiFj8qrCLzpW/syVvZtE/Ja/KlIQp74UQynFmue8M4yq
JK0kLZwsV8r01ok1UFG8osT+RSvjWimLtBS6krtIhgkHnPBQDmxGdvdFR6mUskbW5nwoqeGOGLru
6O5StMf/F7O2NuaOzoP2pgMHEOpCIiRVGsS5lY62mIrRgpAD/yPWbo/gKi00HAS37/00ETuIjgp0
DOWbJWrm8qeSOXAx0PCh9b930PC5XWwsykoE2aimAS6ORKS2AMZ8rbLTe4bSNv6wV07RzuQVilI6
4isDMqSzvpm1Mhxa+z7vNF7x9GQAPe3j8fYW8+RJ4iOvaID6a2BFEPIbQbG9f4Qd8DyXGEYDjnMI
00sfTDGnCbp3U51ZyX+460qEeoA+8Sosk1ihWjBb3x4PYkf1uk1MPh4U7g8c+UAeAP0qWr/1GCNt
EVqLFH2Kgf3jztcZjj/X0/8V3QVxIvGpHqKxLNoNFokSYVlcVaot++XPwIgxKSD+2u4TsgmbMV2N
H/ERzYKR9hBjdmxTw3MGZVvvlFW4Yz2/nsiFFFD296DXXcentc5MH1gJ0wN+Xg8GoVzmCzM8teHc
v+sovcu3JORQv4pjpm7XJ9kZjddOg71ttBZimFnJbTLUqrJx/Y9G2gZHW02eFFA0u2hZV/SCyJD5
P9pqd8aeoHACZAZazVrBxelMAAuLd009LK8fFVxMWKb/zfBe0RccrqW0USNcF/4XuACS/bHBajkx
TaHDEewlVHjF1iSlYefCpqLN8YhNKZ6GkiNCY8s0wbJNGXMSSn1QahimcTRAx4sUpa5Cok9SU7cK
+XJGYqTNkr9C9uRZ5s9kFH7XdJlpEDBUjFRPDJUcSWobkpiLvO8AR1uOkVgVKj9c9Tomwro+OP3D
JGP2WFb3LrMSCH9umNVxmdzKzRP5NmpUwmMR9KZaVFw3MnPCkOb5BfiOus1EcKKn3cYGeeRFogvz
zTJzhzXMKy3PQ8hc9oxBejGNPkbnqjxOPejinHb8ksPbo7CpEEQzsriaOylt2sGyWI+EK5K30uxi
VKIim+HR8MZx0TK+dyVN1CxWW8NO/9PhC1+34IQTYgxAFm0eKx1+NAu6nFJ2YpaGgaeHLt8iaqJj
n3gUzZWD+dw7/yAW8kyJr0Doj9lW8313rmAgoCuh8JbtFZwDroIrLmSi/GU7ho3qA88pi4V0J6dg
4zJDvx8qhYxFVSOJoKo7EOc/L8XaQdd38KSzKg0Wu7F86XxTLUV20EEiJcX3i24Jf2v42rHINgUs
RfxoR+na+dxxDACmAdDcl3O3/nxPJcj1ZSsP7m4P1p95uNJkYVLGEME1qU2hNH8T3eeT1ekmZsUn
i55hXYsINipwN3DPL6nWfVEOS9/vh2N5JrBWsFMuXFPIeLymPPexGnXntUTzmGf0jD5RcJvZ2FeP
N2U5L+ViZPpZOlSCWMAT+KsZN/6gXUe4zEZ38Nl7zyDXmYJ2TH/gmPn3gfI4dElem5tV+J9GOEq8
faE46MYF8YZ+LbOXa4PZpegAwHlrulohxO7VPySarzGBeCUrOpQ10lM1F0qEaFHKI//kvtyRHjDV
zrK7vGbaKpRIaQeyxPXS3KMvq3H/NLXl57pYe3sR1oW0u+d8o0ZB6RxAalLEOqyk34FScoL/pCFF
caXOb3q6vBHdcpfOr+nDR9I2h/FMAnlp/aZedqnbvHLO595I0PrVGfTHXpjFj7ElIdepc+wV4CtN
pNwJd9ALjsW6wekSaNhK9i41GxbDZmyG2swTFMBZS8QOaQzuZ4kDGfwTTBzK3K65exwiHCOxKm81
w1wx+2HOBTa9CcJ6Xcc//mGSXkrRtaxNWF+O7zjmqWJ+3gp+zDAylRPKYXlG+XVFLNxdgPBv3GRU
FEi4hw6v5fWmq+APih2iFdXoixr03ldIK3Up12/iQk7MdznJJXgNZm4zQEQSSck70mtlyqvSBuqO
q8hfUNTwhl/SrWWfJOPAcgK8uqb42wcbkga99ifMsuhkicx1mHOF8L/6OZwOnx/6w8QXoN7I73w/
SEja3KTBLSL9OclJmqp5G9DZ0lNb+ptOb3hAP9s8ckinKnwnKOv7xIRgqjT+gT/pW23z6awCzdub
frz2z6cVr02UgrsYMmLDUl3fMx95xCVPeyJII5fXDBvspbXmixG1sBllrBtSE+EU1sNjuIaxjPv3
5tjvDCVhz9a2OBwCLDS5eFYQ1+pWK08bRNhg5Yw7I+/z51VEKZG+c4Cze9aHmu8Ymi/omJ2bC/aZ
4w0lF7rsvyXa7tVRtdyaLusAfY6SHvi7zb0wC93ftwSRzvqxUtoGP4i63qK4kP0KhedsbGCshM/X
7k0qhm5Hv3CBOe1bgMSToYljJCrJZxz6wrnGGgH+kmzALUKQ+UKSVRXb2yNDh6TSoNYOAr8LDOiq
+Dk3F/kfpFsUksWQOG4XfB2q+oj80UNjFB4o2uTwgkEnmlyLdGutvpx+u7mfKCRZ6YoK87cZ6aOr
FgdB9x2VntISposMOEgLEQd4L5z1wGjPZg/ei4oco9xoGCC8M6SPR1fKePSdtT2FbUv593DGfNrB
c/H4z2GYsXYbf0OfQSj23weeFzOr6cg3JRlKIybY4jNNrJiJPMfUD/reSbhDMO6iOdOCYeIMRZAa
E1FjyCunPfFFgTuIVkOl/gX/UPFG97+dVIalkX7JIuA59pzLjOayNdk3gciIkeDMHqc4cM0YM76B
UfYcaavlE9Q5QG5ycvIxL1PqVU+QCTZNgJ6Kw2+5nddJyaKfPV1qHbbFRwdwIkNMgUt5idIoAcbX
aLh0h9Qj/ng3oVtyD/5GSd62VNwy1U/9ev1xErGjkAssuypWMYmLVnYa8YXFV96IYiw0wAizGXTT
uu57/fBgXhwz7pr6Pr2lEmjiiir4zryhDv9rKQ/9PvUIKixUF84/xOZNG3cgAX7wEToD2Hb3Uj3b
ETTz2skmYUcYJNKPi9z2vgT6KzpcLm0DvdW/Z5pRGO0gRlq7TdP4XMOeNajoVjapY2lLASpwycFh
ZH/plpR9VkaYOhUs4sQfiTT5ChLnBax9lZYwORXyJFPJe3XYTVNiCgZx46VGOUKj5ygV+0a6ChDE
YLqV5/nFbh7gqbGnBdcimSiS1lb8QhgJuRMt2Id58HFVzLuOPfk6gZohfgF6iHDeDB0ak2Lx1fb8
tpciuDaLCmwmTBSWH58rVB5WT4k3LyLCbBpetg30J3eCYdlJNXb+P3oU44NdsDUtthptAQ15jYI/
oDej8Uh44W985nLrZWgA4olQPs0ijDl54vkAMtl5OLhYS27VVz3clPuVIveHEqzYe7InKnHUEipL
q5P69VpZhMuAD6gvDmR4O6Wi4FrTKyLIpEgYUQYXZlK1oduVv1KPPXvl5IWSnf0oNhjG1uf7zJID
7xHPpsx/FHgz4tzHeLy2ildKSTsmw6gx0SIAitMNeQhLfCBuGQM8B2LEFH4q4djFMQq5T+Ntg2YP
dY7eJqGCYO7oIJXgWAql+UIWXSe9zNOKQJOTIz6aYNDc4eYjKC2XWgoZ/PGSxAB3dS6FiRZh+OLh
9jyPcEcE5cv5agHiHkNFPc920HJ33OvxUnl53pWkslkm4fNVPn3Ezr3HrApcpdcB0R+K3nGhvTyX
kaPa6jw6Ue+vb8t6RpWWSV9nkwpStz6tiPfcXiFcFqQSPZSqa44blIkewER3mAkBL+POsjwhHrNd
d4DN96CSh1JGHvv1FgdL99PsSBcdp5yhvaUUEFNZaBkaIEc0npJtirQ+rEx+bfZK+bAnSvQLKbZ2
PdrsLEicUBmiPIlZ3IQf1O/YS3j9jTI6gCVbh6TCSirdPcuFapqUbuM+Gl3t8RGIf5zU5kpgrWeI
sFnMMQaIpiTp+tGtQMkOLA1Xx/4RKRUuInJ78c7ai7JqdABFH79qWUDYxdR3mJ+gIIROXUaUNmly
iBzy16x+IiYErrT68Wag5DwMYvmSYsKUgXtbeH3ITAsiiSdxRSKmX4NyoDBTVzbyjVYoHgiolVla
t9esy4SO6iGPkQ8+b4/54Eothg6i3jKaE89pxKWut+5Mk75XshNAVLopXHZ1KkNaRWWzRGDfXmvv
Bf3cjN4auYYYfj8UgVMijNodLLY0GxQFAXc7CFeMYTt2qUWiCMCmYk/9ubP3RWS4LFTWQR8alo9W
4i1m3jqE/pCWdjSgz2wopb0B9dt2ZFKoxHv2C5BgHgr36lmXrtQD1mp8AZLic6GplaxTsU6uBkoh
MqACvdD3NAvhXHeAvH0CTi650tZQgWG2oBc1itBcM82zbuBaOFOyvubYjHFkeQ4p0xQ+ofzJLYek
XmDZpFhifdB/CDaCJx5ap1Fj83WCDKcKLFd7246NWxRGK+yGStjInBwwO9nHa2YPvl4QllyM9/z8
RbGE81nTHp5nDssUdQJT+x9BXCpFG6iE+uc8e31Ln+M8fSMsyBO0uAkfxPp6GRALY+exuL8ERJeQ
+lDBSkNP44Jmn8dYX43uP8e6QgXWcGIKQV0xl8BPf4htA3f2daeRShnxgnOsStCZo/NnxAvFcRgW
MlcGPjRKXHEsiXAMyPKuIKLWI+URnQF6xHvNj5+KrNxIrjT14kfmMMejkjwQ6O0EEHybubSWz0Ba
rxw/Ah2vNGpug+Gc1/QSmiQp4m6lCxzlN4tuhNaOIVmQv/deAdYQ47TTsiODxrss6LvKpjfNY9rv
qBLYitPdy1p6VmOWevlKuQNurxeSMkPYjKcR1/RFXAMOrIFdStQHUB6ZhKUiHlEIzh3EzuWP/+Ey
lJV++a1NrVJey9YrtT2zgWmBi3SDyRsktLrveWkqWBiQMI4xDc4m/yStUL5L7conYwFS/HNfy7va
a9knfLEUyCb2+5LI1Ny8lkdD1U5ZRMHRc+4+mcUbpbn6cVkkZdVHlTAUBHUh9Sm2wsiZIq/gUGoM
tIr8aCpej2fuijARGPs6/99OiUvmhhcN1hhkHh+cyDa62cx/7ZNGm7MEDLOcslM/w7Y4yJip7txT
XwA+UMP8iYJ4a8oCTxM11L9VFIekOws3SG77Yy/0+LhpsWpW6cJqWCqcrEbX2nwWLuoulzMb8USi
fZcaFArXvbDpUbBgx8r2nYNeSTGP56/y15uy8JhNuxxMxCFt4FxcKx2PMAHE4uXY/DzsuRbs79BA
wqEJuJLoVBDeVe/GzxfSVY0AF5lc5LoU932g7qkgeTydyXMafRc+vF2tV1LiBjIOZWjea3VXCoRJ
6GpKVpmHdFW5J8QVv57osyE4Kc0f6mQB7JIRTFG4y8AXuC+f7Zh6spabX9DjdVSl5Qnw1iHjCBRa
tV+luu80h1RK0oe+4dPVb2bLjInGTSBMb9Mq7hSltPgftnTEe7/kRFc3vEWCChiHxETTuTBZP/9b
p8jtSbwEY1J8fZo8ZhlLHjjXw7tkusG/G+HNv+7Q0BFnTCl/pHKaikx5l0R3LtTt6X9Bj7W/b8V4
21HfpvGtDN0GpeTxzY88MzTLdU4kiwMYeERAMtbJ5ep3LeAZua4LQzDZV70JNi+onGVv2NjT4VfR
1La/GOGVH1z5dADddg2biahzidApUWhu9Y0D09EBWofe4GiH/Y0cFLIwpUv8hwBtvJwcyFCphssg
WqIw0fIIOAGS9avbXjPnUeqXq6rPJnFc/DpMnpPU+PORcYGA68niMI84mdI0m1DqbYAgg4xnkQE7
OzXAJsqNVjcGorKRlMDpvyGEVL1W5EmMnUEUr2jkQD0eIRj6IHxMdQort7FlhIsPZZGXckCiSOad
StHu/icVMejWvGXdlvu0LO5ySo4Tq99NHa8ugSNpXHs+vgHpYejngUy2Ys8Ro94hq38JEANYbUl5
020znDIYPSv5N7rwJJRh9sy9DqzrfpehjCBwZSh4mOWS/mlbcpLwyqcdGrFxFQz9fGI3oR/4YBev
HqheHT3jwlgCUeoM6HFIgWhl4wKPyWkj2vdOiKmJRkJWxuW9SBblH1K9YEJgNk9wTVj9IQtnoEip
CmFH+M5C00d908wdlc22xfOjBGjasG9GxdJ/tNiJAJz3a+a9vXBfnDVWjwVKTROnCNj0oewOlE3C
W4jPHjVi47jzhKq6bxJDyaojRVxUamKyzC3NO1L5pFmsBGSFy+QNhsHq0+nGHB9HsiirquEyDcBP
lE71GNVaVe1HojMT4qt5rqvGObZ61e3Nhha+Udhf0SKcReHPBPjux/93I72YusvCWhGyqYXKapDH
w8fyQNrkvhtuzDkcQQh3fB4P2MK3GaFyniwYzewPCwda6BjgUSRnpySk/UqtFK55y9Dtw2qXeX6D
FB0E1fJarvjMUDv96+LpDCkLMsHEt+BZRnhh+GLLYyr4ebJFyHP1NFx5rcEc+6FrgD/ZvVcivtWM
j6Z2lMPfD4EF4vf5oSGTpY5c2yceKpwZFSyaCb51/JKQKHN6HkeDLFucS/Wib4W5WavPn8JZsmgd
QvF4dME2GoD4iGu85tqJo3Gx4kTswMR35gosK5SmJbc8jU9a7V0WPRfn5o2i2Kt26FIKqFks/Xa5
pG+UY0Os4BPFmM4Vz3y+YJ2CgJPUzHYA6Jt0o9aa80Wr1yc36Poi6qcuIk/koIkr7CdFX6kPbJuK
uYnsT7Ahwnt801ar8FyetFJKc1kdfgRAmlF259Wsqytg4xGxBp4Bs9rpcYbtnY2KAesnjZpbzvEn
p0qV3IGJHzZBndgTP3fNUG+WgMbqFfLGLco2f4eu0rF2GqOpPY3wBsMMeqJYurdJJLg41isTnOgp
/91rj49r3o0Nmahg925WSNEvamJctL5CmewCHYZjMkm4VIvA74oFXOSNVIe4zoaqDKZ8KKnYAHLx
tAWfUnCJvAeZPj3NWDQU786jRp/xq4UCJVlvuLwPn6O+e1oUbUxADrJkVyV4/nvOPkUmZO5+aV2d
oHQAPpxC9MR2314+wDB+EITLimWPFy0KL8wkHUd2of62mdczjBDs1afAT+ddS44QA2qZKKfOM6q6
1fDaDfYK5Jifu5rcVNWClr5+n8cMsJSgm53z3p60uFJOf2qs6mYz6SapumTTC7/uPjHV6ewIzn6E
78Zxq+dn8wgljCDfsAficxPI4CmeGjfFP11BHal77Stui10ztB9Zz2yI3D/9PhsEJ8Au1b+xL9pT
TtlPFQ9TCa6nybHwAW3kaKlc9PqBWDAAlWgNODsg/+v3b3GNHThbN1YAE/fOwsXUg8E0m61CPkUl
31wXIpMohWiYESlwr9YB/6Oe2tKL0T281fKkrjyJRjKwDKf2EIYeLJKDcWSNAoaubHcmom4TNKoQ
5HsMBjTwZOOB94Q974lvCxXQ6cMJcpXIASpIGjzvp+iUSSAQHaHgFrSgi271ZKlMEFps7YZuiAio
TsXRqe3j1Z+NFKQMsFiRXsw7N4PHGGVyGutHQOQvz4B4Z8fox3rdI64Lz6kLKOHceYeh+lfa5Bb9
Wem+h5FbyXsnRY9gOQC5/daiqVHw5ZOKUtIRgTzEL9k/OSdCmkq5TT9KhDekSJjBAeHkLe/Iy/sr
+qHDyxFYJ4g38hkkt44MoNmmzH3S6ycVXUBVmGaloNQkSmSa5PzhrfzR7bhTSnQMwipeabNuyFdV
/0ACZ7S28MNOUr3G/fbyUQ0sb0M3QcP5ghBGq6YL7kc6OOolCH6eY3JcGM6zBfVmW7jVSeH3mbtd
BCEUtUmjH+UoUmHWyQRP0P0OWLicb4IEmmj24LulVioJZQnhyJ+Qv6QN2nYYahFZ2Yai4jJ9PLXa
C0o0DzvfQL650WwIgexWRNdShKzne0Tlnb0RhNdV+ifRA/33tlLvmswcEsOE2uIOBtCyYsolztra
0izxh6r5iTkHt6RNyjJQKhoAvaU4JKZ4v0riShxrf/yRdIhWQZR2FvDHgNb7IniQ9eh54OlEuxuA
MVXqh4zCmwwp3LIBVkD73Juhc45VeGHlQ8dV6WM/Aw5h4xS5bccj1u+0UUJs+ejOgB8hniZXwNDG
g7F4AR9e6wpUcv/aKO/0bc9VYJ8F45iElmBZj8h3JN+eNEyqyqc7+MO/M53mWGl1cMb6gxJ0DtAT
DRdfLiIJZB81e2V72Ggbm65sdKRi+W7/6SzMfL5I8DQjPRr2pHxQwVHcqS82E2sIfryAcSgIjaFH
LlKSZp06Ld0xqIAZH7TXGVjDoAmdczPsu1EIVbdMtbA6y2DkcN+N4WQ5MNXdym2mHVYflH2svLen
cF8B2GommSeyoXIH7oF32C7XeSuurlfopygdKmw4XL2vZXdyNZ1GaFEP5xDtCGOWH9jFH2ENei7R
rF21DseoBzDMHDbpY9rrMHYhhhxTu0w4hLlnlI6M6xBikiiUcnjuMUyfNtjRdVnacIk0/UBrGcTt
L29Q34UhNlq0iUElBEvm3J2cySO7aHReyutO0jpHvjcR0+CFi0whhQ7b3kubR/sHNGeKN6MfkWjx
WRhp1tN/jrLPkBbDwPZE9+9Caj01V65A1ZpPzd8qFPDpJy0ifaut9MnEQsoYhzFZ82MD5bQNj3eW
bi2s8uvQgfIJQGLdKExJcHpQvt5yoxfAvbMwGzgSD1iHeT7D7yNRQDYkvYWP33XcX44Daxo8AEqT
jDIKFbtAcFFqnWIfBu2sZCEjo/7VQo7EkP7VU1BoTzVzeP9taOacwADeILXlHOl0hwuZFzyrmioD
aE/M3IadwHcEqBbFq+HSjKDFdbpZ48B8coxletLAeAe9BuTkWppautdNrGymvKfqNgSqq4SJqC3F
+TJS43DY5THhYbtaeEMElPTElv5SLO6w868OJ4Ziec+ArA1qoo6Gasyi3q3uuLyevemXs3G/Kavp
2LKHWyZ6wHwww3xu4+aWW3cRgS/CnOIVi9vQzQbUyggAyI4fdSENC6LAOtMXwkMd5S38Hyg4PYTV
DkW8S4VHzRfNAA8Zmr+8tMM9/LRzDHwDYQOLqWF+lK1bb91A7qJIdqp6G3RSsCFXJwLgSyaG+uPH
0btgigFCZP+TngwLVLiFv9GS8GF7LjWTwBA5XxMGN8LimJI3c9oVUJvSVi25uTMT6MH1L8YXWtPq
UX2TZErx6ef3yIjhG1Ip44QZb4YT7YhM/FiQQZuC3xh5NZ97TVugfeG8vEjQVF+Yb/ZQGuUzEAvn
9OFPBkpuCQe0oFsoJwYpWdUxJnHNhYTcaEC8FRBoUoUqfpjKJg0KckN0kj+/UPzpPt3vriycEJWq
9sCsDPfMORMyHHDSYqy9vqwnCcmGwiTsHojfFFJEBmqkWJEUF96WfkUQlXRyX6dHrz6gALAvH6MM
kwTQtehXE3thyfqIy9xHWYc7fPSTdOctuHU/rSjmPeDZ+a+cBXUOu5V0uUUJEPThr1Zi4rgi7nNJ
5q6DdQuKRqMXpF9M5N5/MplJuq7ZBmHtquzO8r4QBuHYDV9Bi4+up/fLw8lcCr1J/UI8XIXn4TmY
fIyQC1ytPOANyRCXlZeTkQeWC/LiCAFdQo0HbuCFZrCXkYGr5y4RQhm8ZDvMBobp6sp5Bl9Uvtqv
1sNWeStxoW2a8+w81/XKTOiw5td8Dugd2AB7pkefxzdRnEGuhhJBeSnOSZIsxs3rGy5K/5+Q/a7K
zmds6eN2IAgQvd9PEPa1/zrqS7hqxNM8vHG+gVxBIx2MDv/2ALPWGv68/wXegPkYs0k7lL2g+v0E
xGQOXX5amH8oeo1skR2hSdGmG5nsEAp8PjBMLHloiUGdU8YkfuAIFWJEz7jSKlU/BEbuPPIj5Yxi
/4UJ92vbXGF+fXrG5dyXOK2T97GS4BwjlYjcSVuL/nzyfpDYGy1u38HJEig8MyCBy9zLrjBeWicV
Yadx8Gpw2YDWqFRZe/86Q9r3DLYlLYG7F1p8dv7StFZd32pSTKQUTSymHoPIOc3Da+BWFfj9+CMB
A+93OVQczq7fVrcOc3b/rtcUOhIMG4lrBDuFzzVKeF9ABoFL0JX7eNZzB7tcKy9ORisjME3/FT8T
GT49l+2qHczzN2vIHEOLizNMBu4N3narj/CI4TNMPSyQ3lL68hynXAYHqbo3kBU9wA+bAfoVa2QC
UFZobjsi3pnMHVxKcjMcaOnLhadpfbPFtmCp2kuo9fyZ3UJvzgXq785mPbelMEjgC5DJOhHH0FJ4
8iZF0LiVYApMLjSmWifH7RIpgGmoUmci8xb/2XtEAy76W0PLGv1/1Z8GVmIoO1WFR7y//sVQUjBy
ZMAOsqlhRwgyPyLMREhyzIg9SDGQ+27odKMdRMz+k/lh/3+v1EzHFWmhIgZSK/9bXlOo8SwH/IoX
rDZm9b9WRGuF402krvHctG1bkXq+nTtogT7RU83YCxtcRORJX1CBqjIF+BcvqSINyJVnH5CbGx6g
wqt11wzDgeNrnZShhMbcls43ATjHmn6dkA5a9St3k/sL9Xlz6BDRsI3O6av5TGY9gSoCQSti7qrk
G6+AQM+0MBb4jENuRX2CWefBbkwf+q9ah3Jyk6jk7YUcDEJ0hv0b12jigP6h3+XRZqoCs8PLxDW3
A5Q87vZMEd5Lf4+JWDkN66e0GAyBYhNqTGxpLcUVYAeBAT4hQA0jbvrONpGVpaoYONoi6CHAGUwN
H0ST5cRPxawQdK+bN5s9rOVSxDNbkFoMlUESXPg/Kvwz42SQmfLbMp34YlXZhs+53rLjUGpwjmXl
J3+BzyMcjzsYuHBhnPL+coPGKo+cjk0xCRVyLUmbDsVCopPfHZ3j4kxJKk3fYeAPsYT7LISOEt59
VBgm0HKtoBn/YOJRjYPZkV6bgUup3u+7llgsQRdhf1SPPlBQGNJNsOwFjHl+/LYGDjaux7yPmuiv
wetbH2vVPDJuQLroZt6Y5HuEvQcwm7i2VXCXtwRvAulMDI7Yo3KUQY6VMzASC15BQkeinMkh1MUf
ZrQINrcXE2xg2FCpXtaNTuBWA6enuwZByEQJKuK1BOxU+CUUoG5PeMIj90D6zkCw0It8oP1spZ2+
xqrcWYz6bBkPlS3nN+LsJKUOdHTZsMQArh4IgdOmNg5esnlzEtel//F3Z6aoQteV7MSW2XcV/+DU
hu1Y5LOop8xqinjUw6cMNq/gek3ZoKIgQiVX2RBDgt6f4lyzQgV1t2rwAmVGrrtVf48NTjA9E5XA
5jJO6IVdOjj09hh2scI2w/j19/fppnFyZTD1Imn04/lWQ0S2MsqZrmb6lbzKuKFGR9L7dzMq+8/R
2n+zslk4DVd/JxJm6WRW13wHVwD09iNNvAWbdMsNRFezIkvREXhwERUrLY6y848/oi0HiVpBP1sx
4QfBWRqp+BC2Cq5l9vXvBpsRMJDKhA2MMGQxtxGN9WuQcYf+MH3fJG8pnaoc6wtLjpVgihUUU+Bl
RfxA+qYuld4s3aVbS06kCn2Ek9wdT101u5uGoIIlJ2aLFEtUDVwimxhG3OlLe0YBo2LhCxukCZoq
DTWfcDIFd8RU51b7z58U1olaPpekmuU1rtvZZVJz5jcIbdz+dMpnOGozqbAOquvD41S2KUP6B2zQ
lQNcY4QUULDZMJ4yPSdvh6AXVaA8Ms56a5YgU9h48l258n/6taGAL5ySncOqTl2bDdg33GWl1aJK
GK1g++O+hbOklgDftbXEPkPwHbxBPvKmrVrf5uChEWuPZPBLrFzBjxFExJ7JyklaC9tOfqg3rrPR
Fiif5l2pHmpGCW9MYss2s2k5XtoBmSlm2CsiFBAjf4iN1MDSyW5sTeUq8sUA/PHIlulXoiCCvaqA
niLozX1M18BHhgeQmR45ajibb7xsDrwrSEAkuH1VA+6VG9ZbCrHNY7BBS9g1ke179Ki0iPlUw6kg
5zinb/nwp+YsHQXzud7av3/wCvSxHAoSr8bNYp6QLVJdD4VtCsLrA02CUUFRRreTN3A24h5u4ysu
7Kigw+gIZEEkncbZ38zN0tCz6UZP9Y0zG58kydrMhTH9YdigOiINCs2UDFbt6bsXizHCo9Ib23ze
6O7Uy2fm97ZU1t9mapOxllqmXfutJkffBGOAFEQ6DXxBUS01+G9sRHymk2WMjEYuMuqED9KBuVLq
Ih8GcBWdUTppaKCKGJnJyOkKZjoCQrfUEGpv90vZV/uKsvQzFuUSfk0ml8VsYuxAKn314ieWQ6ZV
DzMK8zle1ksYac6A7p1Yr/OnzyZBDDbsXwEm7ovLIMfv8OWeWFVpvVzNmeoOfTIKsSXe+172Hnss
9Np8vxcXzDnxTN8/z9wtAeqkZd+4KrWkwh+WpjQTRqxdLTuqZ7bFEUb/5u8+H0In7BIGU/NfjS1o
5CyGEm0/k7xMYB1FxIO2iPFrPWVlqRrtzZvVqYTIjUitafcjyECBofxBdvm0SNFpOkjybpdnlIRS
33ZC7k5mJyqUnhJ/DrVIk4xPZ7sm5IaAQjxApYFtlEKDsVYDHR1HF2H+sDpBHe1WDB+rxoHE2lCf
9GUs7KoUJmm8nME08yaPhVNzAcIxgsDGyST7wd918vlike8/C+mAxNX2bzkdTlbwcOgTe3gRIWJ0
apiUrSkAYQsn3lfWtdnBpTL34MSlbvrLo4ExjaSwuoRoCTRCs5q6tc02hSPFhpA7Jf0HHU4t9wHb
9iHv7utY6LCNefzK2IuUI9M3Al4YeratiROPvjnZmmb+Z4moZUBpzArIOK75Ifg23fMAQvDiXyyl
WM+iZ4IuQgDswiwmnrn4HCOXw5akian5HglDE5FSoo84rc2QQCtezXrt/irHVyub5gNkPz5zBR3f
brDQIapjdBV54TAX/Wq6TcvQdPLeFxuggKWHQeawYF8/f2GnZ1VbsiSYb9S0lvcOHOaVe9p0SsVf
ZhDEqNV+ucbhILvvrTYoJpXKDgK3WTV0L8sB/eGpznxzSSvwScNZoXGm0RdHTNbfF46gnlnWMXMp
W2yzQREbfIoFOA/URW6/2a6Hh59wyB++sMYmL0BauhcwQB/bymDSFwZGT7HRvnmHyK+ghcofzzh8
WfLQ5GUuwNYWY6OTGqiUvxvkMGxr1GxLqWj4cAJz6+/OYbFjBTDJNme8GhE1Nha4JhogPM3D9YNA
SAeFeYtaFXhR0ZRmou3gYM8CQUrqbVPBcRGYwwCNpXTT2u4Aq9L2AYaV9SWAPB+DvJQoBxipOHYE
F1YSexxenZozY787arclEfJKVgVzIC33pSmjUN6II2TJbrDvebqk/TaV4+zHfMz/308eaozewfBY
6MbVPOUQPq+nreP5sydQlfGOCjQmwR0Mj56jhrG2cex+V5yqHZcme0huMpzaRtOinUwBeva3LCQL
Fv33wFtDqE4+1xCNFW/eBfxmp0cSqqIJ2BqtBJU6iDCkJ8YrPRBaCb6ewxNkRucYBtyjcs0rEXoJ
KmxJBQg5g9P0s6K66XOMwYX1jnF6ZwXE+kImoVgrZ8sG0l5IRHltu/mon+4+esOGzAP+2r79c3TZ
MjEG6lVBiylyda8uYHrghfzO4x76HT/gkYtpDiF/7p4liLx56NfOvxQD//6ylHbGGFTfpmh6rzPt
d8J5i+PtH/VlwiQgms+SQYWG4CeikTfPet0dVoa1lQZPNdgSnmDFD3yOJfy2v/AfZUdkKi5XCQVv
jPgmONZ9G65kq9tCMDDHy2JRzm+c6kS1k2PJFJsKxhX+aLg9oxRz5lsuCJH2c0F2B4rXBScMguZl
rPoP//u2rO0I7Mg/Z9uWn+f9Kgc0Xm783+sysS2zcrtSZDY42H7PWxB24EIoeHYA9RRAne3ZBnuP
bQqnD+adtiTIKnLmluzEL4Di5xsb174yJuvNrElKpphAO/K8jlNsj0qF24DzAgKOWAwpg4/XonER
p9fkZiwrg8wTWkrlBNb6ZPrKNeSV6RT1FUo9ueyou0RmISL87E1zRiwhVsCxtGif7zyIQkg+KB4m
SSzh4+8FoeeMSjnqfr+W7QstT4Bpi3awnRgJIS8JfadoP36Csg6eQrLb8UORzSd2BRo7geSRo+dw
ht+ulutcLuxJCM+ZWmZmuL2YcY57KHXzahEaIjQVtkOVfWmqTehEc9zCcA8Ws9j5Dqk5AUdMII3B
E1snobu4Z+zfjwa4CoUqZGN7GBfRbJla8cMRXdNwRma0RTe8lHprW1DcawD9yA6RIv5p+AFBnuSA
BZgQLvgrsdBrxU/aBHlL424g3m/x/fuBNjN20JpjTs5PE7cAZeHHpOqdlS0ECfZg4FflcqsgtNOb
VkaoynuUo2WZ4eiAEQwmouk8JVLVfcF/XprFRRA9EjJ+I2tWj0EqSh5dfOyE8G0AKWsSpkX3nJq1
AViCnbefleUhlb0l48Z/FgBR6/w8SrgIlghbZbGWJ04TYVuGScmCf9JJgVVeEB9v0u/sNMPG+umn
O9I0cTkusA2S8UDAelApDCgH98w+rXyyORIcb7WKkw0vk35iGbauYvAON87Rta5M8zLlXRE3l+uE
3lsXDjIZxGu0CloD38rdZsWxWLXJhSw35kIJB82SQbexWI14e3somgSlGXMoflb2Bip658hKao9o
VY6SMIOAJ+oahfiAo2uBvFs+yU8t3ERuSEcI+c50tLJXaENKwQb33k0AojRJg3v1Fo4SoHs6pWnJ
CdXLvN22SDjnyVbgsENpbm2NHOvXqSl+KFzB6cPIwL/u2SDlvHHZDAK9qmNEGWXpZhLktVvwFzgC
KcjTjAL8HSutgke2xpOAqyIHnYpCKW3KlJ/mHVvpU/Ok//o/0llxiHBeFZ2qu7iFI3xKRsE+h3DS
Vh0FAsRBbK+5GOzM07slGTNM/rowFZFlbrJNlUKhqdqntqFEzrFrhkgv6T8zbCclmkQ7/MjIRmcN
HG64fg0YdC61iTlpmqpxL0Oa7MQ3/mU765lhwhbET9ZBW1DUXogOX+G8Vp4UDH2hDiP3nRFk2gtr
IKh3TYy6/Zm6eVrJjbRISO8FWPqAOib9vSLY8kelVFncdF9lUw6B9rThsjZUJKirH4myFyipdSwv
9tGNJA4ETfiwAg855CwlK/ePQj/BCDvk/v55GsOr5qjB93zVw/wpQrAwT+mgocjHCIwEgAyQqBmg
I6DxQdU9+N72HSJgMcgv8L4P9Pa95q628Ql15lkEo9cJTnorQP8I+sNC0+KA8a4CGSkHIF85Jf1m
HsGk1JgW4q3THXyuSlDGWI/b9iCT0UA5r/jJu42ySUvHBL4Jud8cQSDcOYqSzVP4fXsd9b1UPjry
O4r9XHgzSxHS3ogesuS9unvXzdtBWKaMJBQgydwHxYYkaQmLVR0KoesB1yzjqU5TfV8gWyo5PqOw
cAvqDwCGDPIEjA3b0J/dIMGnhV5MYHQ4hR7Q+RIThOid6WbH4jNhFLyxylPwcLS2UBfVAH0NziTh
aWqzvQ5qQVoGWPJYUVDNYUwuvwlkFkNQXq8kQC5XVYLBg5v9bSTJSAxFpUa7wbW0558PXSVU3wlH
YPSBUJgh3YZQ0Rs5GZeNT1y4IMl8QRCBCSG1BFUmWPCfB8sr5pnDdkaed4ZWDWknnIY72po2BkdE
nBctmmE6f0XNA7ht9w3r0EPXhnaR48bUbFpTH/wtzHyMcfE5WRjSiWCchXOw9cJcMvpqvydIlNew
pW3hrQM7cicb8OGWGpS1cbCGeiUVzEm/1gnEAMaOMYr4BNYS0IJnFCf0K16ovkcmDJvEQmU0bbhm
Tyw5Tp6bvw0Vnx00GhG93ySNrN96bUIMR/xxin8tXGnu8n1EiKwccGAuozRIFD/AnzGpAtCxxfgh
xZPnWTEX1OmCpfrwPNGIfM7pqoRtd6eMz3PeHQvfKnZS49J3PZyf5sRlwb/nGGmSXHg6hS4+GD4J
hSreZbpsXnIvPwarvW0mavxqHtT5Hhkhf4n/uPSAcXrUGVOr+eVZj4F7PMWus97BtTZ0cCgEONBY
J4BWOioLMjTni+sgIVQLs2fgI1mqS0dlfC9dQlvUGw66ddQamlNrlqVztBhxJ4ebSKsElblQBpP2
NGUyNe07lIFmoqOdwIOlqzURH7XYNoSvuHKuHRbL0986wEZN1u+5yk+dFCjdHrQyZ9hbOO4JbGIY
/6HUeSSD4laz5pKkLnOZizVcBz1UAC2iBrIhXkrhJpWE90oaFnn3MB7/JZbFaO78juWKEQjrTXQP
L95fGGfCvagsz7LIv+7M/gqQeNJ9Yz8mQjx4rGPZi0QiHI9XKZQLXhNpNQ7DwrfaGnxHHwAHvcnO
cPQ766Obigfg+4zAeTd+0rZwKI4jC87ObBymRpyVciv/TYXVaKkQvUsTEP18k6OxCpdCVOUNUo7r
wUaQgXUfTUJaF5dPpHDoOcD/Pq5cNt0ombXwDdI0wFQ7WFXKEDcJoPviIvoyuZQ0yCkuy+jqGyPt
UGaPwBIAkqoDGeYJHdWYzIkN0G8sCAcrGko59CFlszTA6aDWHqbuAnvGkeRZeZtsHqfnmSGONZ9M
NaacZMwbdQPpcXdN50KMmqHQdBZOe61TlXuMR/77ZuGgg7ol+mlDB5BbPle9aErtd0NDuz0ezknn
siwTcNC405c/c56Ko+Dd+dyFZrBqPmgquWVkC5uLUozB3baVYL65pp0QldBH3gMZEj+DeW/ktTZq
i1LG3j6q6VtJb6ErU5T/SQ+OhMCaVv+QMLGniWLKb0yxUKLJBpJd0LbC1jd8gLPdQNTQ2XVOKznl
gDD9yE1D6BWr8WNpn2QB/PcPDGrV0aExxL7+WSMSueD/3kRLToOKXHQZwvXTFxqmADfuL96RWeOj
ykGYhHjOcB44n0EKc1YD8V6qyvik/TLPQxT5PSWdigeanLJF8BM0oxi5KOmosQoSgkrgfTR91V0d
k3fSYAh6deKjYFCGOH9luutk2wi2hRpFf0+IoIcETrTft+HaNCj4io2GHl2ilt35ozYW7yf2Ghm0
3ypvhdLdJ2NnSrLhh0i1oWjLJnM2SfUmKScDxXTiy69H7B+FcwE+wiK8AT2nmc2K4wk7rTMdAlr1
jGkqoSXYVBLR64aeBiW6ML88/gbnpRZ+LDybfSZVsIaNLHhRibtmeHxWjFfvalmg8ww2B9Hl1iHp
+addfPNvxQFEyfcgRCmDfdvWg1NZDsFgs2dyd2YtyRBFVNcmwSzoA9lFuWTqRH6M4gHbUtNWMeNA
d/Vr+pIv2ds06nJYlBeOrS2NPlFsBQHewbQYmxRPlOFu+gi7SW7g29lFAgFqrLQp5rzT76Ep81c5
MGT1MuULqI9usu96vyf9ZFlWzTeYVzDCrCwqtfCvM7a26W3mipO5OjElxyOraHCHr+M9yI3enJte
MKBAW7k6lUVkVLlSRXDWMYoXv8zz21VSiBnv0jJm4e4Uhe2D4xHFIHnGBJCA44ubsSpOraZzYVzJ
9bIybg70/kSo1OzleTf9OKuPUkwHXIatk6OaKcujGQCYGKQ7dW+A1ooVKF6qmF9+Uc56KTke3QdX
PajtoxuxvuOodKbNRH23VBN/1kG4/Sl+xULm0f78mQQ622xkBqfYwbvlxeIdt9dHUUHjsQ+wqGyk
71eDce3bE9vBqtVgcsCOD/VxoIK9hXQxN3q0DT+6v95VBhQjq14+FcPmHHklBaoc3VNvvI8I19qP
7rvzaS74Rhpa5gFrJNeQGswYw2FSgufO1NlyByPBYB6LfSsgZhk4C0HgLdGJ3Z2sn9Nn8iwc4NdW
/HnfkGiFBc83Z1pAhQ0ajNXykv4o2Sd8dL4uM7sTAPVDoGalQo3PIxEuJl+NHA74YvNlRviqtICP
2J/qdqtxJ41avecHjKaC5cYU169ZWNfYL8pL2ubXPRm399PrpqhDI0tiHuQq75a2cnP4yhu+RSt2
QnnkrwO8Gwg761SohCsabTMzHmLnw8Wl3UzUDVWKKlHpU0lA11OWz2oMxaacKhnkF+k4HtVQuCrQ
/KtCFBljBwHZQY+stHBcedEtXUaNgFzp3VZRFk11fR47+LlZ6lMYi81VPH8WLkdFzCjD0k72AvkM
hAfKUMpwS+2lcmhrcFD9POCFHO1a/lLIlupa3erOZzL1Mg163O+3WFnp8lIykIWbwzApHHK2ATQ8
LkmFFoLNgvbvlBKYTgTCjGNLNgBJ1piqtQYLhUhyT9pOWxbJV1ek462cskiCZjvQKgqyIt9pxKu/
X24SyfSnbynH4FHSNMZT1wtNgt4PDjhbkfKUVKdbmgRYIRvHpHLjjnRsslUIHpj+eBrXBbrQ9GSP
MPi1exYYN0P3hnr1ScTtmGqAbC9JWN0ZBQt04e+fVyAK+IbyPzQ2bq84pKEQFq83V7ApXa82AYmL
dFRYX0llqW0A21llDl1ZAZ+hgu5JvfjZFT8vjgUQ1qxmQiAXEOKQ1WAo5YEHsAKNpDFk4U4NhWg8
KfQs5dVn02Y4+zLZsCFEVsCgH5GnUrh4Qtk8w0TI8oezJEhE2gTSCc+lr0gLxWIv7dF6kpdsBzLX
O2LJQfO0OAq5/QbAuJqgR0oP8LVEynNzRm5qsbnCyMYdPf8Aw3JroFfOvvPmDw8wv98RRBFW9/Qs
dEroMlqESpP57Ou4AaokviJW86rNPqrDnZ5XFvyWgwyP7lWq/htmfw+EtE7odWB8oZu0EaDrcMYR
2jS2nKULJxS6EArbgdAMDQqUSNbDDAdYuLdgk+Qad3FDF68UGoLtDzcJ6p0ozt5jR5WVbuGLZYIX
T8eEuG0uIuMgmjKAWM2jqSNpqPwNbnt1mjhEXlJvFxYT4Xo1QpJxs0Eavjzd6Q/EMQewuTmEwG6k
wBJLUytpN0w6aeX++TSr946THiMNlcbMeSuuXp1ZpDAjD2SQ5IFZGrBnOctg7ki30+KhPlDNwTQq
Ozte4vqMLw//CFHKTikSOsWRo8icW3PZuvAwNg7aaYQpLQ/Ji1W+5P4wbA7NHadQHcPFTmP7r5Qt
udQ7Oh81N1xaOtW01xWuiUcH6MG4r3zE6zrawg78Hx7uXXOI8IacmcBUydqOWe835TWJXTWeKFef
OHdxrNYeAaY61H3IHiSuG8ARUiZ+9uYSHNVFqJfGLpsy6qf7o2cfew8Y1KRJtqyTG3K/XolmiVCT
It95ZlPpUjkED1+TEiZCQK8Ft6YBRNq2gepERTST1Ro6paTfCCIyFtqtRY7NrVm1mjoTFCPLlAfV
7vYFOrnTb6Fmi2piAgoW3EhfELBzN12CLBsw1lXa9pmIT9KiBSdlq0e80dJrjNY0aYKARHti3fDa
GOcp/Hjfo+B50cSC7Fg/nLHevxHAtpEULGLtwEJPSwQwhJeX9F8sugzMjrl3/7vT+2DAEmMM/fUG
Bwe31EN9IK2z7qybXjVrSOBuqxl6R0jRHtRMmncMEfKCgFpyngnOTlMHeTdt98z42Irx32ZY5lzS
LgKoHahv+7iYE0Op0DBmFa8ZvjB09oOPaex29NwHlIeLRXjYZdjBQ1vDaG060VuXLHP7Ndfcswco
3boxUlqBtreEWkMrPZsrpu+ac/80vOAgaan4xv7tz5UPItqSbFbw7Dsz1rAxfr7hqrIS2R9769eW
ruTwPsiQvZ5sjDVQ+8pGq6QsyJtXgzJ7zOHNIBAG9REzyUYyFrrpIQZy4pYbWYbAhWQglstcSF6c
/dboVN+GGuqxe0yQFchnf7ZfzRp706m4iSlncZ7d9uspjeboF+wJHQQLzioghhOC66XNypPItROv
O8gtBO4GJh8dKPUy1XHubTCAgmN/bEKCv3k2Bk61a4KxyQZqJPf2q5NRMmsEPMkGqqhLDnv30Zdl
Zg6TJWJCJQpWmLBPYIKblQmcK31bqh3iANS0LZ/QryOdrbvPyiT3g1Z/zbTIg3PT4OmoGmMarjZk
i+mXR+Eer2+S3CUql1TUDAhFFTiw/PPs6F3iClcgjtQutC4DdjMfhPmMYyRRYieVuhTxduTpu2nR
JD3JOMNPkDFpTah2mFQP/MdA8tWbNpPPLKS5t8UlQWzdPvIr21AwGkUZL09LqVAdpExkt4NEgxdD
dDC6XngHFQJiyNjTlbpW3KzXy5YopMqEelcfGXbcdbLrvAWocucn6qQEjasmPnPWuBI3gygm9GIA
rpn9d5RdAovQZ8eRdLWSF98hIFUbX91MKuV+ZJPLIArPK7IFdM6/dq4J2/1nwH3BBxKIm7wU+2Vn
3twzHjTQUptmdJvrQt0AZQhqy03lOsEQtPCti7c9gGMghGK4GMM5wLoSUEbOyW2kmT/tg2++WZmK
IVQz7IhwYJrMwsQOH0bfBHc3b1izTUjzgxvcjqVn0+IbesmHu8sDW2wkz901QQsuesCgI0ZItcwW
8KRMDRuaF8OlEEImErvk0UGaJ/rdvfJtbDQFUOm9Kn7Q+VlTDvT8fq7P8PrT+kYU1HRvx1JlPkKL
z4QlAWzbmFwr7GD/f9tmMJLN+7/hetaMPNsv10KRWvPf7XcbNH5PYZA62RXyJXqAzBMe2YlJBLCH
9C325ce21/SnzIM3laOpdNGVcQyBm43pd5nG+Em/K94/2SfyyxZmUBrjOJRklGHZyJQtjtFSVWa+
8rRnfOYquZea4sWRt3kJo+Q0wykcOtE3lRLl3cXT2bnYBCg7f6ij1RCPnpcebBHpJA97WnHsHrMf
aPjTq0OjiDhQyr5zLCFOXCV+KQwr4n8jp94fyVAGwnere69aGXm+zzjpoPufCWIRREvG8oiZARtR
HAVi8TRmxEyncrN/pgJXMX+T8mqgbjcOTiR3gIDzemAHmeqXwwRPQws8+sjuQTckmEPbQ5/wE0dU
2Itp3yX5kGzRzkICsYVJVRq4f5+8AsnTjupaq1LCya8saYLha4BJ+gAozOS9zygtXw3XNrnKui++
vXug9ziuiP8D2no0RJe1Niy51fuehZYrX/wYcY5APXI1JXqBHcsRtzCBT78RebQGiuikcePZp/Ad
Tptyl6kbo1UHvBMfB9w8U9wALn6amYzAM/0dw2RyGNoVd47G2Ns+XKejroR8A/32I7XpkRphqj0d
BzZqhdm3sVP8gnVjtTjDy1BxLDadjEFWyNPKcAV369fylW9mSmEncc4CI4rvGydO2PoUnMRosfle
25KraJkrP4vUSYZKAwB6jZxgNift/DjarY8rda3k0jjp4owWTNo2oTEd250/QL9rYOZF0B1amZaw
D2ZzMrXwHiXXjHCRJHLNKcD4Mc6q1dMklK1LRH0nuIXQPtB++wCP6druq9SoQIqRLvXmV77b+ybY
FtLMBXpzGAzE3jRLrz3DALHInt1kGW84LRrzRjQikTQCiOp7HXA9HPEnZhycijFV5R5r7Lf7EYsR
meaRziNp5xkjtN0GhFhoQaBpr6hYRhoT555eb7uEKlpERWWv0/DiYdTeyyLcrDdIci8naSPWxpgV
36quahnA3gGO5Vf3LU/QpOtvJXFPEgR1jpERxJdf3SsfMENr120uVrIGRm3t6gaISbUfXTf/D9JO
Lv/yezsfH0GQ3Ed2TuYHEXYzpX8iGbOEmT8cYLa9n5JM8mgY3mBvFaM6lq295kzKw9dVibUyLY5i
1gN6MQVk//puKcVF9OyibsEJjC0jb9S3tyMJ+bPIFDvILgD0a49vhTfYyRjokO2+J3CxAjvHOKXU
R5UZsgDkv6urVn00EkxkhlOENwdzA4UtZX09rdOTlQe3j9hKxIPd/T+lLwHWSPOLXBse+rvCyheA
FX9l/ZWY8rrvH81Qkwvo0agBBgpaKtsYT4EoMJKTxoRD2BhWpKuML3c7YB/lOXnDiuoHWVwwypMv
on0Zg343HHCvGkrKH7yKK0ncAQM0h+5rDA+NwNB4xMzh3HgJ5DoYLyWdbp5pezfY8Hi2gITPlYcH
NsUAjseJTq7hsW/YvppYSZxacH03pnahjDiPUVnLBzRHYz5jJykhIMOk2sI7QiWTxi2C7MVTwjg5
mDKTAq7vPw4bf7kuyRw1R5Y0XOXJtSUeQJPpUK+Zna1J+tFh6Tt6SYa3pElLpxlTrKl3Fx7K6qlg
VFwoxzNzOnqgSs/mw66T+hne5kQkwPY4wQvGBWpIoeGNbHJ/56eAXj8qzUuoojavhJ/D8xsofDmb
yko+Y2YjijUZ8g342549iNc28UKM4GEtjmkdklwwzzTOuCLoTklUlNcPUP0GTR7SUHzBkD6OJabp
gKyAH0FO3VTynKuLaWnj75vUX9uiSRoF1wIVjkGgXjMEfH1jn1U2yu4OOoTuz1XJE3Wu6ZOAVXOf
jffGXRSQ/NUnMRvFZTruaqhBiOBN5QsTQx37scR1zeDAb3jxGtpjGkvM83enyDfpT1D2HaCE0aEC
g2zxx33FD5+DX6O24YdLDKWO4JN85yxkhxd1SrwcG/Y4fIzbkRmHbL4/U5t00ymQw7QZSfnswf9L
VN/ws9cRW5U2DAWdIX8KxdkE0NbOlYrIoHPftWRVRijoOpR1ENQbLMCDcLxE/u5EEkJJRQ1qumy8
bWhPNCIHgI0yHkjYutDCITxumUdPiYlLYglCPdHSK5UQGxBEk+k1axQT5xIhzWU9eJQbyEEsn3ca
afmahk6ON3xE6CcByh9jAlNjJAI9BcCkq0AF1tHqnnTHVwBD668H2GKqjHvcL+iWOfmmeeFBiUl5
ilzxSTPg0A9S0PAUG5ppYXEL9irjisVdFJt65PXGLO6tWYTsQ7CAoQQHcQlVNwZRuHM0LM9V46i5
2QwmqIsnQmPMHAypa1FMw4wAKoCwa6V6HpoI6Y1rNIBsTyFmCUwkTujZQFDKuf8pzdfdTyKKgWql
9M2AsumBHs85PH4oz/XbFyPxfIdz71Y36MtRrAiG/6pNjTn+1waDchJzZcYEUXelU0gJaWyHyrO2
GGOhKYQkH32uyxjvdWM7QJILHfYII1gm0AKR6emSQpXUfJ14iAuCoydE8HSMiaKWNsdqA70y30in
BkI6/A6tvBZgrUpQoSrpfXFciD+GBPCrWREPpuWFzRyuhp6yv0rgv7tYQpaODaNk84kspGjhKZak
gdjiGuxT6S41hwQ7TJHuPDluDM5hEibLXVk/yk4UmSK9wliB2kXrdGgNTS+lYZYvR09eztvSS8/M
DtZYpy4m0iCsfH3XEn+BYjUMg517mT81saqpgeRJ/lz8td1gFtyRDLJLPBtRtKmRQ58Pvr6v0Ri9
uwS0hDRZxjn2Z9P4mGcbyWKx3QsuG93RY8d0Z+iigzJFY/urtmG6EDJF9RHto5extuw87PqWZqtg
RoUQJI7xC2L8vfmgsuyengB4hyJxw4rcT+QfyTLSAEd0X8YAzgr0LgdD2p0LnP7EdI4xOsjc1v3k
wIhqkGVhIvC2JjGi/yQn2UFQ15e0T2hJkVutx13BaiGn6D9l56joTJ2veU/dp0e9ekZM1t6xWo0w
dUdowi+eIOSTHfmmo5YAL3yKCY6BcMy2EdV7pTbfsPbW8R1HQQnf7umNgWlscMsFVPyid/EYIShT
7kh07gBxOAoenaM6ACIvHTeqaNOLx0IFKAq0XcK/duLUWvPv9stDaMlo9/ZYPYE3lPdesqeeVm0F
OS0nXu0vuYg+YqGeHugDlW29bb4pFJ5HMLiykEoGb/zl2CNbmjqWARGmO9oJ4iZ19Axuux8UHqiN
2PB+n2rQV3cyE1naYXkTLVWWIZyBmX2ftjAuUzSIC5IMqPQfp3VuUqj8m7OFUfkUqjM8JXh+AHvI
RoQyuidGxfGL6gbEYHHyZSdGnsGtefkULfYj9TzelRPwJv+iyx5Dej/Mv2XjHFgJUOa/6HC6FfzD
EmHIc4dWkf6kpunkHsoO6f+40+iWqjD3fQJssmX+rUUGd+bwBH6xM8fvlF8gT/0W+2d+YvX4UmBx
oRxSSGhWvSvVtdw7CEOTN8S1gUMab17QDuIK5chK/s6T8ub7NLnKgoWFrL91EdPTMZuTyw+1svld
tx+9EqVjRgoLoGsdfemQFMygNP0UtQUL8oS0QqUP46LlYxpeYAJMtJP2/1XZS7lrRPUbcoRl835z
e13L2KGOaJxqkLRRgSbewLXicYV3QGqLRSj8z7XJAfwWE54mHERrjTg1ysZ1i9Y+wbUEeTo2dIlR
KB5yHH9oiiB9Ru2LZMlBDMZ+GZs2bTPRFrPX/rHTPbT88e6x4XdTjIDchFF/tYrHCMGGc+sWQ1Fm
RzxZac+C58sVhWJVYffjFO9ekFa9eeYMUZbVdisbavYzSxxXqqwCToBmTmiEkGq31Kp0TOSHX/YW
8j6WYyTnAVd+YOP0w+kwvTzpZXYItD4P+W/9srR4i+ZpNPGD9VJlMlpNsj+2xX8OQL8xdyL0RHiE
S3/SxC5CElGXEJ9lyncYMndXn2Y+ymshSt9bTnHk2AdkjQ6sbRi8qt7RV2Zd1Li6nUg4R3zxJyfX
sM9EJiiev4jxDnQ01TzzsOjzUdZNYfOBe5suEGOSLjJg+olhuiVtqUjrJ78JStpkAdDlvfPbtvBS
2GqqfMSNKIQAg/OFAMCSrug8m/93gVqvnMT0aA+HGBHPOjqHGg6E0aNFQyZrL47ErKqJmaV4Ad7+
+fwlnVV6kinlGvdhKCNkva3ihpMKlMyBtCoc0RHgDSzgubTtHiqBer5YfziKbcqFKDAEZivNAjMg
RpLZb0+L3OCpZv/ql1KKQ/VFKSrxqNfC0Z0WSF2+4PBtM8WzrCwkXtsVx1/WJtBhgdEph/u0Uy3G
WAcAqpmSUnj4lQsxGm4aF2gsuB24rmk7Tac2zIjFO4vMkpkIjZkx8BACQfbGDL2DyqXQB5os3RlN
zTxNTJ3YEsesNCGZd/q4kU4ErKVpJoI52UtGmfVdQyG91k2TFY0L5Opgr5SaTe2Li7g0WH1b6Eny
sbkZNWDa+4/nbhmI0jjT97+NF/uPLg4HyiQWdsGjmwpXeU1vcpRRC3MlH6bCs3ruKahRetYfOnEs
GKk6Ms/AmmIAti3jrrLIzuWb3Lf92SFTN7ZwON7ewDjVR3C5ktDBKRfeM/V94sJ8hnDCMrdo+9BB
C2d5D77ltZtvt2xNplkDZ0qcYSQPAzcF1owFX8DsO8ZKiAnwHOkfAhivLmwYMDjfLcZoy3hIXS/g
P5Dr/DYo87JAiwyY5XiNG1a1RK44YwA7xtqgaAIrIfyN/MkR6E7kYqq6b8p7SjqGIi1SBvJfvv1K
0QbrIdWRjVIZXEpi7e5M9OFm/q5a6iwviNBXnlxK2e1JDdEqyOGa3dB6T7xlZQVh4GFFFCegQaRE
XaFuoS7wCKEmTeMlJmstm8sxf7SGxm1oX3FQc/1mXm8TRUK8cPwsaxm9nXv9XRfSqCAgyX0MaXjb
3ZkUKUTbrZknoOL4vo0owHJGPS6p+i+rCXnuNL0s3wqNTB22znSOeSUAkIKy9RPvLhe2zQP3V8wh
oY8hsYuzPeR/p8ukAdbp2se9P1X2Dk2jQI3zRnavGYxSMsG1NYRay+2eMS8MMmkDJgUcDcwskHW0
Y5ex/55+PWTWBuGHgl/8uprr3ccCRtzzDfoA/jLlXxBaKWu3VfOqGoM90BWqRhkFAZ/8DPQaVn/y
LtbH9wlTrtGdQwaZPF3HWStImBPMLiRv93K3AhYFFeRMeaqeiLYCwbUipzMrTHC/wSOztzUAvqJY
MtF8qswlGvT95nPRf2U0Sh5k2eGWVK4xs4ZYfXfh7vYA4tHqJ0VnLfJ+seuRGVGPJXCYUDPCFY2l
i/jqXMRKyMIjrbB8Rpcxwguv2G4LtwxjHZkroRXThvRKCR8iZLepHNCQCjPYmFq2j3mKblfymfDj
roxrvawHydfH369c+UrS3yPn02S2XY0v+ghN/4GB/wgb+kzTXWqQoyDATDQsc3YXXbbiqyIsHZLb
F2cc9yoa5aT8SetrdacLQbwpyR0oBvQliejcX4QWAXrUXY4SEtUzeB3ywotPNHDbLRa8L5Jj6kFJ
vvkWT2FsQPcKzrJzBnZZKmrDoiCDilfxiZF7d4b3iUS5Vmdf0/eyEu7pdGkj1DSM1uwzNuiBOUTX
QzxTnU7Ve9A30EGwFqOXMxsdNJUpkZMWdUUjEn3joKqA8xie5hWm0vu6+Icxj/qVawL11YMjHugn
L/WnggrWWj4PgbOMP4aFYhQdG8SeadfK1+BPQHobDhYvQ965EQON7liBtNfuiJwmWTt6hg3SiHLS
MmVWsrpaNzmmYDVQLMFg8HetJLIXA3aLiJ4FatNrhYaZvLeSgecXgmz5S7PynGucUp00C9P5YTn2
hm36QTGW3vjTVwD3OE+xyXv0ydlyLOsyWCbk4YS+9e23vxRm0R9eR50eGpD0I3PKEyw+1oomftOc
GupycRvQo/WHDif914MKkfqGc18pduNyS0+qwstdaNII7n3fkcFubNc6PxNTI7WhgxeIjD+PeKz/
5tiXmJLIgxA4/tAkTuFBJKTrrEv14ax0TN0517cZIAyOojHzNRn4a18Rvsg09GNj4Vf1F0dfmhfA
pqj3zl1VEPUjLGoM8k/ozHRcQd2M8cQDCH/6yLmnJJjsmlPMAgDvB4didjk44OhrgF4jwefumf3C
THTh2m37Ey1AGoLnJVtdomrp8eZnYTdrWbpxh5UUBw5Nup3XWND6TQ0k5Yj8WRxxJANi8cPcMxRi
epL3KUc+HQkxhGus6iXkFu7wr/vgwJWdQEv3Q7LFLbjCH27ZxzpznmfW8XLnZko/0JQSJUbU2+ZA
AOZYFpfdXAscD+DyWj6NAn3Nw3OSoCbfBIvzm+7IVR+vVWfQmBNMPU/Hr1dTBt7J8gGV4YWjFVt4
ByLx56s2SwNMI0U5LDMZcP/3mcC7kxMo43MCNHQx7rezF1bms8ywac/lP/2q+s3hdBRETncAAM+f
bnxu/z8FOKdv+A5cNHmcikKVdaitQz/oXcihnJ5pLs1tzJsqvIkXttzj8ZwDVMCXbIvj+udiJ+R1
YairC46auFWarZ/eXb/J08VCy+HeR0Q89KPOZdiHdvvQrUBqSVdAc/73+hlxQPF4qUi85ayg4d0/
F4/0dVHk5iW5OdX3HeITlSzupId/TnPEDQowgpdFbIsd4pomHeixk/l+MzQm+j3f0s9mdnwwR1ni
WjqQhvIYV/YPeQTRzGP5BAK5mbXoj2S3T34cEImtZyvoG1JqZzsj78He8S9uwZmfJsbRBWFHe/rc
EDu63KtWE3Zw5w2197c/KdjFv2G9xOLGYRoGxrltuy6wvEkvL47u9zCuPZpcu7qfqpJiA2aH2O7D
jOGH4Ha/KGgEHfvFpAHMOzZ6HK0I47UmsHNIxT4yNDsy5vB56yd2K+ssLsf8P2vBjCL3G5QLYCUS
IcZ4uWcfeB2wdG0K8iH1fe8lm/VWJqdf6AxZlvH02QyuMP7Zi2t2beV9z6FZLT7gn8A41MTCabSQ
Ss7nWgtl9zgUmMbb9nwrfHfBrIOcoZtwkZhSuI9muToAt+oqGKU50t3xDIpXewfFCl5308Mp5JtE
95PwPK1hv4o+O2xIfMbOek3JTAScO7F9228YiFtN1yUj7R28V4onsov3+1nbqDRNeIELwgQPFmil
hhkl/Y7I+8m6bqM9vu9cjnL9Gy8MOd/FZsOdq64/o2vU7/k+56PBXR/gACUVvPHtBpZaHJyxkgx1
szdCITTiRVKgBPIedq039rjzfmcoElUao4mqv2ICnxYeGzESwB9N2pi3Hzqs/qelGnqr6fh2yEMw
bbZhH9eeShYqpuqwAXjsunpVMRsLuxGezVhw7dAYVo1l1eJLUhjh7gs4XSMy9ck0Bevglav06olr
ffZdKPvbY2kHpavaT6IzCNGPbboMzDwaxKZYx7D85LpU/4dIT+FNil4S6/L081wZHDotJGOyFrKH
mWME/05XL8NUDqdiRov4KjiOJe6OvyJVflANt9oCxEU1IeCYlKyMi+8Sc7vQL7XtGlwRF13c4GKP
/cnVYs/mNCY0jwO0YmEJLF4+pfEftgeaAksXxt26nJYWJuiArJv6AZETd29AMKN+ZSesIbRkMoPE
mJEBfXLnJ/xQjo+oxCFoGsvXOyW6+8uBqxg9GZO8G62VsMwdAMVb1OSTr1GlpJHkEIPrJCHB0fKi
/lV7sUBxj3eHOvo13+ZAW6mIpVMc4DpgWOqcYZCbVvZ4KJtm/Ta/+REp3RAN5w2Rxy3kczlDtDRb
yTMstbLz64yZ85xPAWhgyN7X2gMXDjgXmTOCspMWBvc8+is72d1tUkgY+bc8vSZSqXUqniGjIyzl
gwJ3canWkdn1DcoWiE74sPG2gVpkVI1A5fgpqy0kq86gtAKl45yMtNMqp0VVSJhZrxh1jvqudjWi
x2PvEIXkhaAko32mjRWWJMnPK4TOpsPS9gZ3htNmDUihn1+zBEFRt9QIAJhE8y8A7agJUl4BoPDG
/mNbgQ30fkM6aO1cEeJv20kOa+5kq7yLR3YbnbGkGlFaBGi9nNV/gd2sggGGgesYQIH3NMq6g/6y
Z+34h3LaLMrrRvmjIIQTVsQL2FU47dABtBLXRkU4rExYSaUaeQiliBIxgH0vbTE+6gIm2P0pluB4
BPuzErSlEFDXJSsar+sklDh/clVknM3P48Suwh0r5vcYzYA6E8IVLLx8dpMPuDhR4AOulEUXKJ67
ynS93xORCUjNp/YKXuFx7gv0J+JyA1V7nBRQeDvg2Y/+12xIyNE2ETT5q7ToxXWcis426tANVTNk
Au1MS/CmrIEXSL+46tYh1s8VZ4IKctpUecCjTt4hjSFlkOURfMh7DnvS9ZJ7eM379RdsqyrFuwe1
4Bba1WS0QV7rB0GmI8FrE3RfRbr8l4jM3FptYrEwf0cLDi47GUFDXRx/qZfdvXxD9S6tB8qce3AT
HtDb1cifJ4Cd4iVXy/q79g6QzI+fXHP0+Gy9cGsgar7Pios1XmHdOS9Mtb3iWqzDweJFa5fWvOIG
JuSR4xw25zjTpFIO1K520zdvuIJy8GYqk6xzpE1hdMWgreyS4DRuH8VTesd6Tnc9a9ZSEIjFGHI8
URIAykoaYCu6oSc5CnoXFK4GTSfkbuZjn3BoxzFu4h16JsIrvspcmhcq5VVEarofzmGBWTmt60wU
wA/WqPzn/hhl44qpNo+raUWN5pPlSq0GfMC6coUY8nm6YK2qcAMaUFzy4tWf5bo/RNE063IjraXV
FEh/0HXz9yzeb1XFES7ZFmxqs8cvjx6VZ6805YQvLIsNNf5Vrzd6LALW3qE5xJ+ZpNfaP55bC4ER
Dz86ryRQe/fQT70a1b9pIX1cYTf0cnbNkpm+xcBQgRcUnE0/l2ZpULYcQtqRAsW86R5zGCOp55M4
lN6xkdFmQPxJzLi4ckBOo8UhFSS3JV8+pgXoUa9zBuiAAKWYrX/yuCBtyKNdeVu/ExnOfJvGpi/6
ha85qLObC7las1Zyuu9/Zd67Q1syRmA4+RTd0Ne7SY0F6+Rmm+EPoXythHO/sl+Hz+Hq0Ilhazas
48YOVtu3+e7jCCilebYFJVBGxNOlsqeCV9fmfEOADxSxZ5J6kbVLCiL3nujmBsRsQKeNYJf2fseG
BR0wFzkB5+OqftkSdd9e0Dj+JZQlvzi1VjFlkOyPWxMFlBKvnmxfmFCYINQzodRJNrpYW4tqlTb1
p6uM7/Pmn4DsMSh+UDVpKRWWwFnPiC7BQtycyvU12K1A5iCNpvjPsYy920p+ncvTB6UesKimQiGo
q85QhGCxVlNTik39xJY/0AFp9yv3O4uGcgk/ypYT3Hd8L+waMPitIi6DM1qIBI4ow7/V9ekaWQ7L
i9Bjr9EKSlmjodLogJjC+28hD1OGHjQ+nmt8hwKbRRCDKtVotdXB+gW/ktXfzwTkqWPdwnHmlmAg
Mv59aT9zYw5HkDU/crI3vW/wMlr/CyRxxbm8fyD4F5qdTk2MMLkP9xuzkjDRNF67NoWk8q0DI5Yf
sf+Warw+jRpw9ANluULX9pEjiN1eIcV+wySObsGGslalaWkvDhkOnkZ0smsmElEHpdGAd63n8c7G
H8J3fU2tl0pN/l/dSXgIr4cGo8SW099+L+XBfwK8sKJzxhg3+MJ6rhDePggjlI0cU9ZrPAuhdEVg
Nn36SfIhEwy2/9Z/R/l1qbWX3D4dn5klKUIUjgnz29JgZ76A89tGg0QnAvslGudPVxHMkwRN3/MY
kbQgXj84FMgop7iBVJIWkDEFd6+ggwBC54KF50zf6KFvFDFLhqclbPOctd30MIDDycBlg6HzWr0j
4zQzIvCKsRcHBdWeoalUPCnRTqRfHtu0+dzuX4x+4qYycRuadnm0apheoteLM6dEmERlKJ/SJo/a
jGNbZK1HixNoevj12d0RX3PPRgXzn77GONYghpisJVrsPEnW6s6A1G5WMZI8VOK6FFz4ibz48nmi
9zCpT8IVybras1oX79zG15FU/ptrY7R5+pfsfOZlQskJYD+CE/Ltx/dBA7GwjjpkQJTxv38kJuCc
YY+0RjazCq2XPM69uiki9EAqE19m1vq508C8ady3MBczK06EO8+0CgM1CiTydJH8Oswoob6f0IbE
4EImRFFXxgbd6i3ja0YLrf6tyPaNwszR/gockwx55OxgouAFSEoSzFeCGNXrrpirgGo+3uA8UzSk
ClKLSaDXdko2pxw3miB7Z5ym+GD331RgwfY/EjoDBz4rVviqci5zEBl00ieS6+ErNO497d6lJrZl
l1K26fH3tszYh3iHpsZCGleei+bCdBliSWlFYGvInsPjH01Eyy//VZpQo+BMkxTYw1zxFpsGiOL5
Wa7mALjwLLjxfq6A/9TJfdZyHTs94C5DC4efV8yswAr76Bpbo4A0CO1ka1bIbcL0ujiyDdmjyUGP
fgo5s/SO4hzdZ3JQN9pPsUa+eVoQqDtMV6B3FgkKVxBHjxD70GsgODxpJINvWjOp5O6L332zGvjU
4q7GS685ba9l3OJgNRQJ9kzXAHtv3KkwDo3//E9wNZHAqJlMm+SLXMpTvBJEHOdatFH5WaneyAgN
u23sxarZETEZfnIGKgymvnNX1/gdCrGehergTYFnVyHqK3+InSBQZYlwPl8T+E9pKB8oHGyYpvsC
6BK/McbEHIKpBXV16+C5CDagJQlUrMoqUlVj+o2A7OvCUDrOrv0N8RLol5zMJA748it3fd+xdV7Z
Ba9Sbkjx83rH0HM07faw+1849FYAu92eJduPh0GJJQ29q7cwbJrkTOwziZH10Tko5lhAtjwZpbpH
/+pdc1wvDM+qV77ySsBhwhdGNXFTT8cfwpUr+9E1CGsHmRXOr0eINMuN/VjH0LyeJkMms5zMarwX
T3dbl+3xuAmxJDh+6UlcPiF0cEmnKvFHkYNZs65tZyzUYTyXBtOhtT8qZsfzics/37OZaa1m3IEu
XTlh9pyZFjjoVN4WvNh2ggly9iA5YLobmoZHWxDxLWaPgxAis7Mtm+HJrBHUGoJTWOmIh42z7aKC
G8iLTHytDJGgCzn7hUtNxlNssbKiWtxIGqxvHjzdeIHTArB/1iRuw33t5pYZJK/Cr2qMpEqpVsxn
ehVblkeHF+vPuCHk1/9hR4jfAteqpjOZf5MBz/uQzMZ73V6EbSQnO9t44rC3MVL9scoPzoxBre1y
ZgBlwQhZkVtIbIeuWlT7qgrOzvCA7sR0QjflbIssSIjFvaLVNyGjeAL7+be7JS8KVnGvZF1dThQQ
adgy9Nmaq7KLstazDm5LnPnDs9DGMXVjG6W0/LmOcPK6Ykx4VsuG1tiSas1RF+saIc3VmkvbHjLt
B6hmoMFxyOw2Yoqrvk7KOwZX1+nLrNwdRjr0zH7xxYv+Xdyx6xg6M+nuUDyBzwgfqYHnW7H1qtFa
wl0G2ZTBPs5j42dh+QfuYQOkZgpGq3tjkhlABfzOp3QrHCheybwOkHl82Z+yJPMWY5BGH5Bwl92Y
8mCQIE+f4kNVAKcpA5GlNy1U35JP9XU2BEdh3tPHyfv/imlptTNFrmrwrAQgJom2nLsPL91nxmMD
xdloULQSlTB9QI3X25TGPiRRebUlEhx472rZKzkS+qtxaTrUwkFBSxTApw4+zpwc7lVKUU4LMmH7
6h/OHJJXyVJNaj/tgTBP6qx91rgoiQUlGw63IdNDrSpSmrvfswRpGQg/skoTmHDv+C9zw/+3UE+G
MiCDs8p07kp8zSCAj3GooLDv3wjPWV4r60EIyQng44n+kSJfFCWicX1VPt/jiwvHKdaA8iNm2xpc
5Yi71tirL4wS/tH0wnkwbLrIwW9fVFKpvqG8MUeUVpdhZ8IImzFtdH5SGqmdbjDkUuTm4ihvLcc4
k1OicNGa5EB8sb5jSilg7sK8RT6fgheDNJDwwKSMXq2jgBiP3tCRi8leVE6kNJeEkiKnWS0ks3hF
MCsCXzGETF0MhkfNCLf1/3BR8nwbyCMyJueSkZ+Y0uSd/tAZ2hwFMdcJaIk2Lr7ZF5O3nC8NJ9qr
CDSfqYuFnwLYGIuoudHexD2ynxkvHWEF2rrf11j/RUsQcMotvyoamsEKKL3xf/UQ+fIC4Fq1KUxI
JV+B+3CYKWwaR6utC0nr4beBVQcowPfcjTYvt+fHV09e78vZky0kt+1vP42bp58E5Usze6xEQ7PS
ejUkQ0/Wd/fhPlf6gLUNt+soQVAm8AHEDuNfmfOeGJYGqDjXzrMX7UmfahBkhxRR83J9KojJbK3d
yP4Bj/7p6UJbnL/IQvOsQHebvTWWqM5dY0TwtSkRxPupkyFnL+HijFeQNALAqvD6YdXnVOVaXE5d
WD4s53J+jEU75/Du5CIfFECUcTa96PHw8atk+lKCU7u5EzVGkCZBMGdnDlTbtoWIQgkya89FULSI
BTBLFMQcZlmLi6Ln5+i46KEc1y5ooQGjyqXipuL8c5yE3uB48omd09bu93rsCLwNRjN3iP1jsf31
DomvR2SbLYRhxPtJZLQ2UdnbQNrYN0Diah7Kq/C5m3YtSlhJNcwmdIeL8klg/BhXxD9iIwvIYqIB
PBGceqwX1aVszgtXzC8HKabnvIdvJF1jeheJqNLvGTyeh6twr9GYmNomuDWwysSGiL3VI9HWh2ss
cj6NlePn5quuz2qD14YFyfEqv+M0UR8bR45qQyp5IX6upbUisBKDmDpAe/26Z8IiwFn/YNDkTieL
v3A6NUSTXg53kCyKpS4DuJNseQbPOA77gqnEYQPBtpXJByB27N9iEpQuCMhPddn5yq1e9z7WjzI6
rSDQ338nf2HYm8ZQjs8sxJxd6/NGh4LZM0iQHQ8MvsZt/Y2drcJYQg0Qr1+a1ZRCWOWTLMoXGmKW
A+hkPovJmydR8gm57vGtTvzkvoQI8Lf2xGmzLtFAraiKYLcR18nea9NCHhcrhr/XQldaqVtIVYrt
lJuI8tlGIyne3otROGZH7ANfqUBpI6toD76wxWDDOnMWc9hasa8GQOMcfoHnSuSH8WrXVAucEh8o
C+QJ2adO7owIcQRXYnuEFGc4KU69KDVM/RzChvP1pqpZT9ELLv3fSyYN5K5841CdC9JHE3j90k1D
nP5IKpzwnjqSME24RQuX5tN7xIVBEb4pzu+TsKUzk53k8OqcuC8FubuVC4PZKPfStFxriGCbJoZ+
9fGfcxEGvoWPPcJhOAJba7B1wwX8NDxlX4DynwKr6N+Ppcoz5UXFgCYOp5ct6uixsgEgCzyZJt2M
H+QUYbtCYVJh54s4VdGoddKCo4VsJ9YHMEt6mnVfUjfgukPE+MPvT/FLQuA7tk1mQC4HvIb08zJs
ZwvQdTkOI25Fd52EPE/t5SDUV99AsogcswmgFlwVH4t3Ug8YKNubHrTAAYsf5cQZr6EOlyNYkErX
fiqgzaG+/Ak3vSO8NMI2Sd7ZSgKn4qkoPbPqJvvHeKwwR1qIHY0bR5wCZqB7v+h0du4fMApP20nU
18TiBFKZVEmDaL9bJmXZ58sMn+9mIKoOYPzz+Nx0gqLUhyvcVfLBuybfe2v1g3TBSDPhfxShDrsg
AXPJN8ethDrmXDq+zdxcQFgWeBxlJ0ZJ3UysoV+SVpM8ACj/SCUvvmQRThK4WXsuOoXUqa+g6KZ1
seAUzooOcM8t2qmIavBCU4eyIFuYFQ1OwxKxmsRZrE0x+e1GBP4h6jXuDNOkNViH8ucizzk+j2mT
7QaFM/HgdWUaHgyZb8AQuWcUGVDLHgGizIsdqbK/6qo+wsEDRkDJtKcwp+nlhqootcshmC9eWNuy
tfiqPy5krAXxsv6DDB6nyHIMmLyX0dtCxPhD6w57gplTMvjMxBTIkLMmaYg13xAMBdtiApay8NLA
Zy2L4MmSyj2M8fD9AKhOc5yA+Oi7Wpt7DHfyrq+/Zg6ll/2Us6Lg2SIewQANg76OTnI5eJAac9hE
sd2IRLVi5EK7CaRgXoc49gX0cFTRNgtINe+9/IA3VuirVMbdcBxWglpRr4AP6FzgPf83/i6Tq/RN
6hjkgtIyW2vBF1xGPUtwvU+zgaVmIegyjkl1lzhU3IQMwIE6Iu2ZTt8nWmtvTb0f0LDL8grmFmbS
euvDx4o1GY34euc17CwlRGSrN1APHakMG41bTXSQ8YRQRFggD9Xvq1nnX5997wrPM0KzRFqsPeDq
RKhShE1efsV+xfEMKfxXJX6OJfwvo0Vn2do06RHocms7uH8d2gYoAF2xuPMaiyL7sdydvq+N/vhW
JurqIik01NSJjohO7+0U1FzSqb7QYpAnkkCDE4gdjcdc8XA1sU/AfTSWAwtQkl3scIm8eBjrWnxN
5c5V4DOSIC/ViEm1H1KKQAJRYQ+M3pxtQJyQL+9Puena98eGYWSpw8q1ce2nBi10e0zu4NDBGUVM
9dkVIyA/8j5zNTrHxZWoQwegp1Ow5VupLKAWnbxxH/JHY2jKjlqzODeq+E4ALKtc0memgudT1Hlv
Nf8FP2gnwHqjCSZwW28/Nydd9BpTqGznv75tH7KUzlCCOwfXFA27/Ct4Ojb3fDHE/v9pn2i7hgH1
S+BsKd0D8f28S+VUdXMSVF28ANAIBNBfkQJF6YnJFqk6aQDWj5+/08O2XvbxCn7QLze0nIeyt43T
gN4qhJ6s6omeuqyJokK4yzGxUjxTrAGkt34wazE3q9H/PIzPuUZX5mKp2f3tFzkTCp8IKGSZpk0z
UUhyKc4yqDq1HE+voZSEr9KDFJGSb08XQlfn4dfnJfOU376XuAgFQwsfketAaVet5Noy45CEv+/U
D8bgghWfxhZTROxcFTaIRwFDvsXUOCpBZIHk7x39jXj0UcSfqaXtmckhuITmFjeIYxiAUFE3NwOD
R6o70IWiHi0FfLgMtaQLpPJSEtBPlEkzKkDmvxulveBAG3nIkugoxYpNGECO4yZ4kbLy/iHmCLwB
zE+krwMsTogukjLbJs6qQLO1xDIarWKfXw4HjN9M0hOKVZmV48jdBhx3CxTS3AVkeI+qpqJjZDyw
TSyK2mH7Gbsz/YqNlJAvZjgbXNqetfLUnINv5Ppy6p4ctD8Dj2iyopV8OGWAK7a9C51JPI3nwKmt
xsppB6DIAqXDXmQg+AbMH2v9QcNCNUG00gXQgXURzi/qed985LXsmXY6dvBjr8TCo3FPjir+J6Uf
dROMffYFB7+m+yGITi7+Pz5THxxhL5cfQhSYb7fyAkycuekCwSV7ziPhKbhqRioHzH9oPKkHv/MK
bgI/JDjX4+BRJeNUHiJ5Vm/5b4sDxnHO5AKphlTlPvsFis0GwIoNNVmOVuu1tpC+NgmD6t+Thyl0
9kEXWI+sT4UMlWlurTrv0wV+w3Sjdt3M7Jx8JNMMXE9iPZWQv/AC+gk/5Vc+cpEsz/9aCD2j227O
oDrEV8eCFwFUKlXNCzhbHWscGgWYq6pzz6ggGkRYXmIhi5SPuqtPDiBMfpd8MIhPuOSfKZuKgsrv
thwho8IAe/9SeR/I3lIxtpjNurxABfyUU1NI2tvNhK7E3XqCEa8v4PieP265JpBBL/LEcjD5v9mt
qQxZfkBsr5jOAiLVqJqFFsqIoI+4HiMjinJXEy46UOXThsFuRXSdPZClCMtk1yHyzSArpW1b4HK2
baFIxHZwUU8KPk5i+mkQ4CvlATygoPqfJa0O7Lx9m6eD8HQwawxdGalAOpBdEkrFrtcJStrl8WUM
JymubGOhNzEzq/iBw9i3mFRs6ViMsUoOmKNWte6IRWmMmeMVuxa7OOc7lMKVncdpoL4VkXUvPrL+
qK/WdiTCr8dMLfKLJhCAEPY5+oJpDLkjgMlY1FhRtJV3luryIlYZ40R2N9c2y6UTT7KmebS9gtM4
IR6xAHy1fHPA3VygChC6ftI7x3JyVKdNSRPpgOHoBahL6J5QnmpSfWs6577bexf0vhKzoi3OZeHA
YfSDEsM/DiHfwi0gzRnk/gL2fiRN8eoN55YXFaBnsmpW8thW2FM4eFFA86jnlX6iS5lvrNxbos87
16pwTC9tYYeQqoXorajDC4XFNNzSa4kytcXkicfkEnMVqtELVdGdrGaYtEYnzGPUOjyzoKb9Ljjy
htKb7kBAQZ4anQjpdl5eyRLiLSFdpZJc1pGBcuHuIUCS60S1nlABKz9Y5sUORzEEeXIztjkD03aA
iekIwEgLS6GnNvN2tzI8WDpDsZbK23GsWsrPBm27IS9T8ZZeIVQvnYvUv/HcJMWbcHvI/Xe6upAm
noxN+mM9hPYDBKl7JIBEJPhGDVSUo69BrzrrJSGTcwOEybSyPVqveVbiARAFe1UwbZCpd9R806Jz
DxmmlJUg4GxbvkHATwSAwqySfFtxVmpMs2qqjUcTZmTmpO8dw7yppqCeAf3DeJ/xwkWR+xh4X2dH
SZhd6yptVg8Quu6Q4QGk23oJ9iYUz0c0zE36+NhuhSH0YW9lTm1Bs1ZanT8ceVyZg4o/xMAp86F1
91XFwANox3+1v2nE0QyEBFLCfC7f8uWvZDb96oyuqE2b4ZeTm4ms+3UWZd9uaEhgm/aabG1tuqTF
iX1QjknPdv2CIXTad2ZWy1QhbtF/PE1t2WHv2bqKZQ+BRy3UvtsnC5GZIkrh6LZOc4QbD+lvNRGA
D5f3fKz/FqZl5NwOkY3WVKNXVCYlkuAkCY2/BBHKUp39973YdWfHWw/zJMEUehFkSfF67tWBZgls
CV7NwuH7/tR2HjOUed7rVNjdNGYvaKrM8HfH2Kde6lvvxfu8XYRssmonnu9py87ucxpyzXHJhOMB
DXaI/gTAZvod7wvXMD74gRAyRQjw3BkVlpQCqMHnnqztMSHIne9OkhE1KJKokdw+9liGzxwoSilh
t7TTruF/hAfAMkpdZHkEkk2FoCxUPf30GDzBN5TNU+Dj9KeOrmXjzjBlKSfwM3qWSBU5MdIuGGAZ
LeKLH/6hi4qpx4L7YYiDCDH065j1T9ShF9dBG+XHfWfz6kQtoLC7wmNToCCD/dEf63wNDOefjdCZ
nc0tuaf49BGc+51cpuPvWs6Fr4Wls3EcNMpjwg/svZnmMa48DkawezPJUPumpOacHDxZM4lMnjp5
Mo+3XZh3g3cbGAPg5SCJjiBu8oDymfjOdL0d9tcchAYFthit02oVbYZf/QXtlX1Sq5VQpVpSBBDh
xz+JR0qJKUzLkCXNlf4NLNmNvBXyGoJx+H9efxS3wdOJiheqNdrmcOy5Ibar9EP+VXpyWGeBHzYt
w7tyHi3/CrolqSJ3/dtfUXvBB2vzCmqUKeljWCOQuKPfeMI3ns+FluQGWUXu5RYH+BfbZCLrR3ps
pn0xUERaRF/btCIq3Nay+VIctOCU5XXXOsIil0qpxq06fhOM4zgHYwMb5sUkqUxQEdYaj6afblSa
05Ri1OVDp8ACoVxi7wYKX12IAdNGUSZWtq1lhDZtaipYNfjsirhe4KSNxKhMOaofQo2NocGCAoah
JxER9peominaMyhU2GNX16b1rpHBagyIO1MFFJ1kfJQj2YWEt0+fJnNVjX/23Ak/MviwAWOtOJkR
dnwoKxnQwU/pltUaF6WEQFzcPDU9Yx8APku9vk+yJaxtqhGT0uxh8ePjhTe7xgFqcGfVVdcONXvg
nUkrD2U2L2tvvkBKUQ7VISaY5wyzTzVlLfCO/DrlMJVBe8zbVgclkwcIyfjuRrrdM9Y3bwUYlIds
lrVJsnHwhqCKzyqiMJl/Fw553zk00ctfg/Gu3oeqdoFLrrIwMokmdMKTPPe2XYxad+asJgvu29Cp
gw8fsqOjMibsHC4WS9r60v49Q3e0KbfpkTaUw/rY9BifbQcRAzJCkTEvxXVbNkxNswE5KAzZHtRE
biMfagY1HStPpGgpUa/I9lHhAm/DkrsyM7oXIGO19l4/kklMIMmSVZCRS7maySvfCqTHeDVSmEHf
5ocZcTUFmnJNNaPI8tcZQ88QuPXcHp+yQl7SbICrt8Q9LB2+FJL2DwSQkkqQ6+HQ1EwRPb6LDtMp
GhUkwldppHVRxQnFActpfAMa2MBe0sHm9gd+/XES8iNqW3cN+9h24fLfM5PgjcsQPk+av4F1afjk
1Q7ci9ZjWbVq50R4X6p8lPE/BG1Adw6WvPWa3C8P3I0Gqk8xUVrmG+tpYfICvyKmfHMT7+wOM+DK
se1Oi5ehpGXfhcRprHcDTg2u2oYKsHR+6wqPQPKdQQ/EBfsJk0x9ma0TAtHeF7pCu4GuxY8oJ8XG
IOTie+4PGoq5HpgLVEIH2myOwg+8VciIMn/uSIsjEeA0u4KRn37vh4oTvuJFVYcuEgiIo4/RI67N
fJa6GqN7JGGXyVlxm7YNQ/4clNv5PbMNOrgopI4Zk/UL1Be8NkVxLLyKcHhCivhVh89hhUuuOIx7
KztZI3Kld3ICA82P+vdYdW+Hf4+dE/x7+h4ZhRq9E++3C9Jy4MEXfvmRPmNAq9HUFLu5nJx86MAn
u3mqx500OhD+iZz5aJejroDOen/gHdp7nIaRXmy1vmxToABZeVyW+3RoyxGq8hPp3QpMRLAynVal
HwU7hqxCwppFpcZqXxlajkJBHHrstAdw0b9j+Bjl4N2Q4sY2YEFoBk8UD5MCosBQ3V0EmG1U+yi7
alITROcN2cM9GvlIRaGU6klfPWWWrK+cYk3WtSdKYAvc9e+whrQxGE1TQf32H+mEhewF32pRpZcu
C5imXUTDH4oiTsj6WDfNoXre7ofiC7PekJOuicnzr+UJZQ8nWnqzWZGo2F1IC/MBHPL3MaByfJ59
/rDGBn8SvyOQh/OSg68453E8Q1Q9zVRmH4kl+ihUyQZGkYjZNp3e4tC/3MDwBON8PSubPI4FrM9l
J3pJKKBMRqhbMrU6qi4AUrTMYGDs8jC1/ebJZ6ldNWQFJhy8clUxfvQOKpJkfPVMebuV6wPxo2rZ
rOcCJmyNv5kurrbGnTSXKF/utzHcn3Kr8ELM3g5X1rT65MUH3WJt7PsmoSylYV67ejwLAk+QjJDV
IXkDG+rm47D6kMw/pDJcJ+5aQWrqBQZR8QzF8wfKAhayj5YL7mCYM9ziIohI20hCD0/HKwpr+y7A
o63Nhp4enV/1Szb7igv3GPoqAab/SGI+gWCO9yNEV+p2d8OxM6oLEHLQFkW3WyujnAOT5s50qXHh
8fF63W7LLAMqREm62qvMVYSxAwlxQji7vOM0UPUwwTd2iIcHKRn4ho2Wd+MEyZ4RfSzuObEJlRdE
GENtgJ+JJHB+buPc86AIJWW9USkSo2QNkXIsdef/54k4X7wOmHZpu2i6rZa2nz5n3dC+turOWuir
iOcU3IL0qtC0ZGBMCi8l4IWhXtM1tjbEtMdZxyins+NPeCz+E95XUISMc0C13J5vJ32OCp8PHKVZ
ophrU8d9Jt8nkozNA3cN5JJauINyHpn3lRBETIHhLYY5QD0VUzf6sjPEf1rRd7ncVhhkASt6Ec6j
inuLPwTGzUOrlpwl4lpPC27RKut3kaWtCrN+CEsK+l3gp9iCclVQM/DHCjqfgXRIYDL+ZS5nVULX
vycV3o5plpAm5x8cC4tUYwuSFddvsraTNsskqM3t2HQBbyodM/ZPfbi/SGEUNgrBYcscqSs2fQ0s
eZlMaFFt+/yaTrleqKC7+PstMp4k8swqi+kFR4BTKyruN9ByXtwgXWJQKteWFU2T/NicBix+zBHI
5/a049CCBQZ1hoHyeojPlQd5pqOsukulYaRPNYLEQdaqxOa9E+NLw+xaofy5QQrf5MsP2oNVMZ0R
N8UmeeRCAfffT2LU6c91xas+xwyskSjkJY7nvHeRzcyZhbex17KAgc4UqGA8OBWcJNnfnPRw+jK6
+BstUFZL7/q8882va0EvPTBADB5wWqlgDrz6W1AfKMW+pKuVwyErFxv9aU0uwn5+I0EpVTcfiZFd
JLoXlpej3MhWca+YvdX7DmiHJBai8+L5EYLjc0w6QPPz32CGL9dUJcMReeybWRfxd9zP4tpVSZEd
/a1+delKc3txFSNRBw72+Xa4vVT1mgqtHJkPp0TN8FsDEVAX4jwj5R+78pDjfyvw7JKcEc5lWFqZ
l4epMBGEdp53+IXGH1VGpMv4k9HnoQyLmCI+3pR79jg/3t/+4m9ayZjxsw8lLL0jbg6juW/0SeAE
BJ8C4Kkr9irDTyR0+b4Wj7XpYOTM22tz5F725TQ4vSKWSfX66sUIgogPkwgsdR9g3foaojNOGdWM
4fTz/iFFNdGBiTlWcsS7Vznn3HbIzCk2Z5YoZuVaO1X+wt3UOtGKkUg4PVL2xmjqqw1oOg2APn5+
dN6nqCnOPb50JH51pq0yu6G71/etyKPX8nkKOnF0MEA7QRamDkdJ2Md7V6SsNIM4MUVPJk6Au3vv
jRDbqc10EfriBO5Vwc7QeiJkwlZIwnBI2I202PNwAkLH3LDGSIJPAeiyv6+LhJ39gqtfNAe8wRJ/
JqT3w4wP5Fov/YHMItn19KZoog30ZNIYTPNuft4l+/l7YtIcrGYmQtcm4JeNySqhNxs8ETEHcmSY
kBNB1j6gliHXAAFMJE7UtGwZc5w5l0rSXg0UHb1PDFuYmwK8HmEQoKmJGi+E1YnV7bjLX9zvnrj9
UnJuJznXDdnf3Z7wUgbJjunhmjVz9pO4Avh4KL8RIwizmSBI25AOColL1ssEo1GHosExwBFosO10
0OtjRXIIKTWwpcQM1AVGpVY7hf3vQ6+ce8MJT0eB422QQvwefue5XK6+8Vso20RK7vBjUPYsMmTv
E10eYHN6Ne8rrg1MmXcKLMzz9Jl148Y1A5jajvE4eTBC7zmGBwsdPnRjPLh+tgYPG8ke84P2NoM/
eKZDGvRcK4wNCs3n7MZSnmAX2kZwpL4tkTaT6hUTNoR0Pze1AD6sxmFmQR4P30O2uOEtxB2io5Ft
e1RyW4y/HJvZJjP3oE3PkDvufcT04tZrwxhxQW85cq5b+7Ab/o+chtLmoUfYUIZbU8ODS2+676+z
Edy/Af9cn7vQvr6XozyFJnFvm2k99GZDm3JJhpuk8hXmzchN7VbXsJZxTZsIA9nNxX1HwVZXUScV
sCqe05nvtu3N3uewbfhUq2JcmQhf4nlzQb7xP8ayVr68KgnMIFLHuI91hnWyc3lJotTGsK/mmqFE
7nKlbNZWnMq7rXBbf/nGvhqYc333y+ALp8VCw8/cID7dicwuzWTr53pSpEQCe4qbrXXuaUha9/7A
S+Y5ypZzvg1IZom/LTMJ/jTT060p0+3x7Gh38G8G0V/gHsG3Nvu0aSSM8K3xpuirJF5+okgVZ5Gm
adG8w2HS9jFdPocGD/9l/DZPLo4p+bqgwrEuI0apTIvExAn8nNPii/Uy0NBY9qCdAoF5iHQ98TMq
3dpBQiKOuokncxqY+nMUmDxPI3CwtjR0q6KvnHhJaaqzBwzSuwR5QSCt8WsAwGJORw1SaGxwrWkS
zRHKUumBBB8TIOkMw5lCBleWBRuEu9eBuwmuuP5Hc5Xfz4iVRzhA825rgBUDLrGbWUiiaCYzsY0I
81r8pGVQ/UV48mzTyyOdgbfrW/LOMM31/94pBJ/yqfRZAwKgES8SMY3bgThupgbSDuimdvbziVIq
aWTUR99yzrb3yQuASWFFdVzuvBhyYjk52G2PDA1d5UZMd5BNUpNwZkvDeU1rkugt1zSvXR4Xrpz7
2IeG8RYt7fWDo/kgG3HGeCFCygczx8KEOFzREZxpNHHyV6+QI/0931+0lpljYpdR6LD9DF1tQJlO
qr2OM0+aJRwsDEmXyDab9cSnrqh5ukD3Jp+7cWFC/FfSkEhQ6VVBAvOslrGxDxN/ZrR4cx86cXpU
re39YVzcJKzCiCD35bRqytROR02ZoG5Y4zx2Ps+0tnZy9qslt0eygjBTb3hh2NhICmqW704P/U1P
U0r6aCYsqE2uBXwoVBj7+oEi16oxG0VcPUj51M5ALbEgVkT198RBzeHUJGLccscSjKLQ7QXnPEB5
KXx1UDFl64wkTMziJOyvFqs3xxt5peRQEnKG98KvFDw3iQyqgHQ/liuzDR5n3HLkrdKhJAnQjNac
qJua83lKeGJqIdNdRVODedyDF7q5CxR4XCtvrl7S7IdCvm9Oz1cmC1MU2B7rB91sCfE3h1qEUksG
zPoD5xCWA2odw749CvITwf2Fg7cnkZXMxREB1WnUskJSmgmp14L0I6Joi0LPyuW0nGRGql/QtJh4
vPysAadS8HDVd0wyRz/5UlpNjexz8iUlGhI/TcGZ4uQRoSSsjAygDYGDmgzkR02tFSEmzI6WU0Bw
1UIZ5HCrnDlFlk9uhgtGzB9BsJxqHKx0iTbcwH2et32aZoUdeT0d9gGPZhR/Ov6mjNt04LTglnTP
AOdPQyX4DRFR2vhkSo5bmE5xTQDpB8JvNbK8F4o/SiupGGJJktwz/mzdS42T0iJBlvMT3CZ31teS
wHNQ64jqV95asXpTlYVlaePItgC1/rDRMZWfxnmSEi6UcGblggfPdI7iGpb2Wp8NnI1L/ANTo5rY
kpDWmpv85pHyrTSF3bmRvJnlHsSCVQOLVdnZaaxi1L1gbIDgJDPM6D3t5wtR4WcSSDpJF2sHt+GF
ray2wCc3IPbFtKZdRhy4mMl4zy+b4E96E0ueWejbm9lNs0tUPbNEtnMwG5SfTqltSQuuEe74SExH
aT1wb9TIcKU70GcPgv2x3IPdasqgYVOkFUty+k3xEHpH9DNbWBN6BrdVW4z4+LX//8cTCCMBsASN
V2WCP5REvHkEwCfFHXJ8/Xy93vidicuxMH1e50xuGh36mtrqeZCXHlEsGagSV2d3anD0XyUagdzm
isqthxbtE66P3rG6srXO+hYecDwrovNXS/BNMVsIkbRrF9koI3fLreSfjyptFq9sHw0tkN6osx+6
+9ROzzjUoW4poZ5Z7gQL0izzBATM2Xom6lcieiP1sspPpVZfdWUKEa+rfzUq/IlGif/BLXPKjLJY
4iqzpxTZv/QnU4FOQXB6LJ21jRBhv0UeBwtnOtpSRtKjDGGUWNCg1GfqRhLmaB4x4eSokLNIE5b6
8esWwT5YKaxXF3I08HTsVN+wTbuEK0NFhBo/Bz8r7zhDJO8aWJGTgI2oFGqbc11FVrn36QPB6EHN
+yOd2e6d7G8f5UeqjgD8qEW4MGgyPEHAchb1uRvv6BT9YN3rQNJSef++E07nu0ZQBAq4o1eY8scM
VWZNr2PzxncKmIPAg0G0W2ONd65ZbxQq/ZLWlSBafrMQoLDDkACO7x/TwScLDCHmAydAHbDwoxII
NaI6yF/jVio8eSQIHkno++nWTl5pxrLHujAlgX7tDNBDrGbh+4JpODZ0amW55zWBI5aFnQSxvYKp
5rKyN0dGqUpKXVy36J6VRgo4fYRPPFsH4ev7IZwhnm1c0Du2XJi2XIp7ZDxwVxuEdui+ZLVmz/C9
ebwYQ0+jvZME8jl+KaXXMR0Vn3Uydph2NbM+PvDoLrSV6X2P++/0WWlcFFHt+87wiIeJg84Cy8AZ
zSIV9vFxnmDlecNYaSZ7+anVxu719Q07+6+7wSICsKwZSMZU+oh2fGrwQLc1FzkFAaUK9/2QkfHK
zJRDQoSdxxVJ1L/A6LqZ3O5zii6/QZJgEiz5LDBc+DTUztf9RSQGc03NCgP1XyWf9m4T+KCFUTaw
6jI4F2SPFxYmZrFWbyEzDzxhA1/X1F4gS2cln4JuEsLI2rvPzlOLgKd6TvMK0YibDIWEZqViziRP
zhIkFxGniMhhCURfG6PJwoH/BB8SvjBGxzqFDKiiWqqjzsEtbJ009KstxqY/QypwKyuT4uAzaPF1
4w65k3Vbl1vebdy+yhDHMm+Z5qG27lt/fE3yRSa1mvHVrJ5ke8AuK1LSFd+ZV425VqOnVrUL4zFD
7nz9SEukUiBZduA3sK0UKLKbjSS0GARDd0Xl9c1PXTIkihT9MOewKYrWp6j0unTnwwcTMPM2JNTX
FsgM+DRC3Q/ykLOJd/p519ExDSEzuDNQtQjUo2AjNMUWV2+4fR3FQrPVKXXdtReXDy5n+F4MMStD
Ihl+m9mQL/GBGrN6NcNXAeT8fNEOVviZgCHRtCQewbHcQlhn1Gke27pNSllhdAbXbvOETFjwANr5
dxlITQxEqLrwr3OJDhbyfEDk79xOPDO7sVqxtfGFzgkADb6vvxHUmP0mppNJ3pSW9nI9GHr56k+Q
fozQ2A9ejkD/ke0zCHWvhKcMHTCjYvTryJaOnq3KcutzkG/+ncD2zB8t7+lC6x7v2EBU8vK+7O7P
Bj6n6CDb7NTN8bpvk5G0KU4/oy9dDvczpEOdI6d/ilHMrI4SNUuBipAi1ZlVRSR96kpsYHsnzSQ/
HKDF1j4b4In1enjRhmUrTFIGePxOcGBUUfcVqqCF2pGry1t68X15X7aWsKVUbJx7IMMuCzmOGbTk
1AsdNkhvS/AwNh7DJ7KSjdiUp8l4Y8aRAfLZCv86HJJFKeZOp5j0l3CgdDcuNMUY3Fb84926sbKf
XIul+GZVPN8nQldAPO53+BbuhYVGdD3NTupJrJ29N3JTe2YxZmz+WniUSChf22SZh+d6IlnAdMQn
pJoTF6dtTyl1WoQJqa06X6JQ73Z00OLyCB2thUqmnWrq8+D1GMRaAGlMGSg4qeK0PyQHf5cUbhC8
Z/OxBVdHWaRGlMcZGEh/YcmRABT7OdUNP6qZAbsUg1Vn9mqFbCdCakrQw61C7oVN0FvhLpsIO+yv
JxuG39nf7tdJlKO06IYLcgwDBfj3OTJoIBFbq4tHCpCbAb5ngHVZYN5LbhBYu7Z/T4+xXZwE6EeE
7goXZCCVVzFodc67m5DIFqJArw4JC3NcvoCMxDnSG+c45UdD06VLbC2InqD411qiJH9rbxFLk954
ow4rSEpuWQTp73JOXzFVQFJiEktSB1i/YnC/GRb6ugj7zKUSNcfWgrLXMldQ73wz9sXRkW5Bpmry
PQjoQKQJ75oOjbvls3t+fhBTxHj3526OygtzlnZ0bIz3PS77ipBV8gAW1sE2JK71M1Sf44hCkhko
+F2jlA/Xon00K/a+U/l6FGXHKOIzRkSV59t8AttMN7xfyE8CoohTiwheEL/iR3UnrN1+tN62tusH
YFWrIoG32JmMlFiAUuCnT9VT+r/gVQlOlANVPFX9ml9ytF6M+QZSSZPswfT1KnRGfYgXYmAWkzVh
Sq++/8VNL+DTXHZS25yJ9Q0Kjx2EtPFirtvF3Tn4/jukRLpHMZFEzBnsoLqICCwfCQrvzzWgHg46
BUooFfjq72YlK4l2MhQVYTL4WVbxRmchX27ypJd+3wxc8SSwMpjyOkfUVAQDRnZEXPbvAeMo3IJE
Bi8NbUJZ2sAEVigKmaCE+uAtkay47rcPuWXcSBokoGyhyH2H33vnneqjdHkntARMOGeUuCPNzYkV
P7OWCiHL1KKB/63fbcRxWuJmmf+6NvaNCALOol3nf+9AwbEF4p2ug0Ewi8xzR2P8BoZ2Z0NdcpVX
lB4daHpVAeqctEa78COC/9TFomHTM77vCMd/3+l/WucsucVM5ONZgKZpwY5sdqCQCkqaiwr5kN/h
cIdzk/NEKZwzDQw7iXT/k/9gEkXicAUDviUxzzIYMPgGe1cl+6y4wL+iHN0gGeC/8O4tamF0xsnP
qv7RbXFMao7654r8RF9oi/uLMlyUUiuvT2DUjlATd8KNILEBwT3ZfwVK3qP4DDKKaYgBdxxawHuR
espktUoJjqAZFYAvgtYesuYjJFv5LctdJiTHK0B8zVegECtOx7l9zBSym38N6rKbVORZZcyxt+qT
rSwG/u/5pHaMO9qId/waLBvhVtzPz47zoybPBUassuCEGPsUs2vjwsnGRBSp7ZIorq0/QzGvWs2M
1+k1PvuB9zl7JCYii4otA1SHA/0BjG6fiTQzdPNL3JgtsOSZrmi3ftxzXdJD7aUwxebEHVaY+r0C
xjAlKQn4jNH1iYII8fjL7vGMeNkoKXl/4PTVBx1ZrciW+G7jdIXZ5je7SEmgEjGTTqCF8v9UrwV6
hWpPjj+dBOB6kaascnInavfGjT4oqL/ePeW+icHYQlu8Wg0CYbPX9pZe0gI77J+n9BfMIeGPYxI3
F/g1Hgo3KOptRqkQezzKPJE14WgF3usLixtLxi/QrSMMJxj84WZFvBEO3MH7YntBELe32t2VXBDn
uqTYPHfhfjBynaAQKw076CLsrWM1EBhALmGjRoLe0KZK+I+nyM5IV3VL886szo+YF9JCc5lTOXYq
UYxhwcn9pvG3fngHhQhvnnhDo5If+1ETkEOEHzJKnj6OF7tzsS7jTR9u+N9e6mYzK+7AenpBoQz9
NFW2GaFaZj9THhUaIgItbSbh5X4lEuyg5Z4SO/tYI6htzYUCX+oLaRku9LWOgzk87FZdWBTOYzc2
OzHbTejEvYabwLT9OAuird6l4Qi6wvqFnDfM8zQerih1ba3rHHt4puUK3FNWwp4e+hucW2rqDlat
GmrlfvIBDn9icUZYsEVNhxBro7Jca2tRsp/wi8YyRfq2Zz7pvS50Ejgt1zQSdhgGVy4Mi7UJ3F2g
x5RxhXgp+iyQi5CKHYG73NymhQ1QJp5R3S4cDtBe9vNHE4sZajciVss/7MZpiOpC+VYl8npJNfH/
aq1hFNp7Z6rcwLbRxjkrOXpqvfVqQSKTIAwgEAJ8HYLwGFxpreGw4CB6lPLIR7i8ejqI1T52K8bs
/cUYEWfGbws099DyBhsk5Nyne4eR4DA/rLwgmn2VB7elOScr/tw+nXoKNNUTOHle2BrImFAPvrfy
stos5VdrlUDKogPUh4nRPOTAjS6geF2RWTF0LqYJx9Y1tKI1D+yitCQiXLuOV27ETLYkllkNIM2o
orO2m7ymHW0M6aQ5pzIbpjJ/LVVH4fXv1GcX4RNOsy91GoH7PQoVhw9U4dAMSH77BBAbRUWPzE/s
BflLO/CQyHZMK7mKtVO+NtFbxEtOyffHcsopCmY4Nwkux7TsVOCYdBPWEb2AFzFRLmlyvgZtspDr
90mFFMwH8xcvSHxgEdsX8D1fmdFsq4QqyQVnaU9lPMTr5TGCfSmb3ed+G/wV0UvflWOuqpoY3B4g
OyDa0JtuXKhDYzkuMhYny3Inxna1LvlDJ7QKvdl/EzDjjyWeixgDVn2aEDs26Z+Ln3aIiaAmTLkj
824W6vB2WxSy/oNC1XjZZG+kcsI2j3ppw9EyZKvfMJNcYhGejMZoiXVWGuAmurmEfbxhafbyctk3
qfADQZeGWXYFD5UrhLH+mQ4/GddhJntbDc8iTWvGx5SkgIEa2/r0PDKkQPKS22Ut6MDQ69B20bkG
ujCXM4YlZNuok0Vdup4wqJMiGF6UZW5FU8wzT/PRAZKjSnr4DU+druA1pu7YqWqL+fVZTn2Cl89c
kRXbzm4k5vie0zQJ3c7HG3vR6KZBT9OM7d7fCGPKhCNKxlO1oeqjBcQ2vPmA9l6sAYmkYGHjy1MK
jmhDWfgczzyHyhi+im0pvNFGNTo+04+rBAd0E/D+Fy8R7Twzvy9SxV7xsw9tuTWnAaENSNI5Q2xP
PkOcPec+qcbChuGq6WpnJ/zzkKtpACw0Fj1qYbzL4Z1fhGln/l8w6TOYwjgL+61Kgszr1MuulSw7
n0cX20TliPU2vV03Mrv9VMC8kvuLg/sn9Zsim7LcNnDLP9fhaV/ur9dYU4bG7QWknkpaLdWkWquI
UedtoWb29GZQgTGroSlEXZPHDS3akgsHhgm647b3/JOLh6Fv6+cfWrXUDX3DUOVDQ+D0ddbMQl4w
wHVpS3qEfcqHPqXElXjux1vizMb1H3oVXa+9toJNVfBNCPcrrsq5KkOPyU6kgBKzzOt/w8LpVeQ5
S/utN2RlvZAO93PGtB2xlLkYUGBiA9x78/sGmaG49b4ERAvWmcM7xPVWZrZcY9Imb3MySWDZqvag
24dtC8ab+6OiUaJYf6FzjfENELA8c2p1l/xXzKe9h65+QW6L88NJeS1nnUanrd433nkSz2L0VIMS
GGQ6aWmCbsyr9oJ9a6wtOdAnIe/cXtxmWr/gGmgpf6XusauCBPB6cSVVrXGLCm0+r7EjxLoHdZmU
UWVdsnwYsuIibXBclD02suAXS4+7T3XTsR5ks6UsdYo+QLqsCZ1JxZXfRhg9BJ4OBmTpMI+geKBB
MaFC5ethCgS3N+G0HKdo5Fqr8yg7hPzLG0vifMORoJhsRCNkI7sZOezirL92GnUbDyNjbrEht11Q
p+gBf/s4cgDJswB5DySxAG8kW7tGhqkOvEmsd2s0lqedMdv1Itxi+qLC54Qe7wDtZ+dn7CrRL/Ip
JDp4IlvNIfcN9W/oGbwlMjtUxCixrApnn7uiM5XHtzl4QQ5NDsvVJVAYoFm3axbaO6VBDLf2qI4O
Hbh0AonGsQEnhMhC0WgGVLk69WcbRq2O9IFespM+yjonFMTqTTr5W74CN/+saUv4/kFkSwlDQid2
m21Oj5TsHtZVoh+0ZaQbbwL6FdP4a+VdM36kB4itisE2mGMb8Z9IbB8OKXSr8Ga+71Aicwrvg1fp
iDfznm5XU2BJOuBgP16tARDwsPe4K51j4JVDecoTPAp2CPEVJJ+G6exiYqWXsHpYTiQDpDmJLEfo
TvNlQnvpfh4RqLejNRyzvkoC5tm+3+rKccWZivo0ElH/IRbx4H6ohTn9t8ezUQ+Av5HwH0Byj8hP
qRvbtgyXi2zzGtuIRty+M6GDjCK9iZU5bggA5D1F6yLF0BpLay6GDQyZQ7nstmFNuS0g05hXBefL
027yIXF/aHM42mAQW42bO7Cpl9gMXTyHHQzrKgVEHs4DU1VLWXqxXyWKKhZHho11fsVCCyin48vy
jT9JnxqeoSj/btKwj8GGgGIhzppVwkr0rGW5pgngz4kaxo8Fv0ZTw+U2GFUVSkLvf8PTjcIJVqx4
nflbWmmVtccPZHcx9fqSiKXKnnZJewXcJdi7v1eYTrtwiDCm1JghEZDlFmo2jXPulTjOUIPdnw2g
V450WaFtjAwIwXmNQtDb697HxX+Ajq6gcNLkDEqTlv8dej3NcxOw1fWOUXS3SjwRQ9XqXiSa1swA
9thcro66sBfxte2g5sddA/Z0CRg+CD9pV9so5ysY7LjrzdgELQnQ0GsLA369zRWDnqb1ZsxG2Rwy
gduvtR6P9pm67hI5SjGN3+Y9cSezpANkww39a4tnijV9eFKfkKyxItgIdqTQZKtlX0scCmuqQhtU
61yM/Qm2RJZFeicZ5djTpKqoL1OMIVGfute1lTdmQ7SEhAEU35ICvGlJVMDIbZEYBams2nqdYnhD
4fSSULhk3H9Ene8q8YXoVDgfoubGI8eeZvGj29Wb37dOOWT6Y2C0/EhOYJvudHJVnGeY6ZrNwMxw
fDMIEQZjzESMVtiVmopu1FJhAB5epHbrxNMoZFn3LyGdkXu6PtwbA0zS5o1V/9ovENtZOLje4HCq
BVViSDym0N23QLsUHlR8xXVe2+wErEWNdbY5oi202PFp+z247NWOqB7ns39Xv/wjL6eqJgtE+fQM
/YLY774jmGuaTbgoBNhMucweqga2lcgSvWKasXoVXZudHCHWV0M3Oby70UdurDvW2JBOLONC23Yg
hi948DaMWcEhkaL0M+1dYCH1LmXyDsh9vGZpo9Hp3p7Vz1gsXr3hzCX3YGS2qab+c4PBmfGxSnzl
ly9FYh6TILYS0ME4IXs7ld87u+5d7difdqW56+rp3m8I2BRhHaoE92Nvb57l5sTORlTiIGpdJwQu
euV8HqbQx8uWjKwXz+cDB+Z5tBRo357ph5hPAt7AH5cR6mgC5eZX2Rfn/OMXtcIRFwJA4O7Ylnzn
6WCGCzk3sj5kkPpjyIuisny9LKKZTIwneswiqg/Jy7ZxLv2rg/ljUk6juQ6GPbGkcWYwvHegfMIh
KAW2Wqd4MvYxmYFgWVFMiYtSkaAn9aMIGQDfYeyTdGW/gpjE3Ato0d+S15Af/yPS8POreAkCkpQy
uQeq170MlF69yYkkSsoxGjLCeIj5bQjwSTgjWzUdlbbO8zSS2wg36ruM5YznHf9D88jHUOu6t8t3
B1rezhKM2qU5Lt9j9OliR2LA1RtVYj0Ls2SK4/dsWvFJSlVJJ63UiIBcpLgUrEqfVL8x9fnMvBDP
MWs64WR9hJlj8WerADLX/WRmf1tSMixnoCXuuQ21Tc3vzam/9b3BAiRVQGFnrJdE15CIlY/aiOfg
CqlCSH0UyAGReXHqOdmwv0pZtLPIsnHHDlE07hxqvWC2Un5glO39ngOcZpiMPOXgymbz0Co8FWX1
f2KDe9cr6qWpkidGGSZAjufKQWUwgG9InKcM8FiDEJAkqfls2Pu0C8hZhHp+Pp2K3cIeiYjU6dXc
cKDc4qt8iRqvxFJqipA4s6tEMUVvmOZZLZsD1vgBY/7DI5SiAnfuA+UW7lxtewX060pnsLLYD7t9
Pr/2UlvZToOGJBvbRXbq6M5fH91hD5p3ryiHkF8hwtAmpiv7+olzFxQsvFxIjr9VrmX95r6Cg5Yi
OcGAEjbgjwZCCAmLF3ES92ELRPJ0fX8H/RQx3RgCZQGD8u1UQo3TcyoQGWwvTJJeggO+Wmmy4e+E
Fmy/oy3F4+Tb8HiS3cWEfJC6V4UXi6LD2AsynWTQ/i3J3kxd76YS3deZ6Qyeew7XPmxVq0ROmLWL
r6tkZ94F/pdKyJBcqUu5p1vhSj+Kzj6x7Gci0efWRxxOrUVX7vOYbdmp8P953fBmP8RdC0AuAbKN
THAAqWRIu4VJ6SkyO9PtqXk82t4SKew0FHhRYZ58vQUB7WhrNnRIi/22Wzr9HncLMiCMmH+FpRvU
V/CfKIaYvNqzbSnvTOw45JTX5Y2f+YxwHzlZyX3PtkMgOzo+/JQVo8jRhXOBl0iwbaNBxcbdorwQ
DmKZZk2pL7T8/xGx0/6T9pdTMn8ToTYBcoQVFvRoI13j6tfiSvvDbacUUMMajumU08Vq3CDPdOrE
aEbC0qgu6lLjlMVbU69Zt2UaIfcjx2mauMgBVMkEcfP99F9nMr1/QOcX8Az+254DR6rq/derAX9t
A0kRdRNCAI2wX0SnPm5jWOeFKiBCBZ5czdl1YKKvLjgtZTwEuol0vRZGzrDAQIltuxtY31b6cOak
nu0JRXrrEhYullyGapBMt8C89lsLLYLUE1J99zKKoD4pZkCFvXEzMxj0fuYR/AWW53dqdpDgDs5Y
T9Dhv+VeQNdxIvc0MR4z7h+cVqhA92eJkvRScI2g18k9+R8XgBLzKqLNZtuz/PweVRqmvf28RGcH
Omxw2alAuYoWIv8BYX1MZ9ozZ9T93MRuehcTEunqEyB+g5AQxJFT8HwtJrEoODfVFTtKCTCFdRgT
1Cm1wSjhkH21iTvF9n/4StB8jtaX4/hi+0Go4XIpkjQsH/4JDriNa/cpIm5MlmKkUP48BrVgqyHo
V0MdrVJbkSRTUpXiCEQVZstG1SH7gPVXn5qxfU20puPGyQg4B3M9nZ+YQOpSG6HUE5mRBfJc2kMM
91EQxyL00eKLNfThLgL+detIaVUD/k9BP375XwSR0Fy2dfs+NqrsFd9AMGbgF/PxriiXHoRogmif
IksrIe7SSC9Nlcv+7wYXLcWxKz1BxCCkg+f7fh71xfV9YW650iK7qcQLlAuPa3lmkA+GMnZoOYG4
C8O8Wz+kY6F5VskJFNzAQFVXdRac909+ly/dFPkdAujyQMuLX/BLwkNBnaY+nsIYkY5k9xv5Wcng
yDSJOaq+4ZW3e5ybbwjbxohADbXW511wsF3KtQsblKkdkL0G9qOdxpwXB1AeE61qk2WRIdZM4rM0
7T2tj2Ofus15f888Uw8eriGswJWHvhvwgfhs5PL4t+FZNRFlbvlYRo1jSTOOq5oMBfY4f7AKFtis
wqtisHwmM8aKHD0jKbNFz5axsmsUfu5oKqTwFAKK0ceQ4P5CQ5dUrWr5+rot1UBaAh6SC2jeTi34
np4QQq6gst2nHPedUjEyngVl4bwsTVDyHp6xKXm/qWoCTQ8PpJE+d2MkpDjGzOV8/KTSavt+qSj+
xkjR6M0C57307iiK1PQSGMsF5OBQ6uX71SXxDNg6hfgHOpqy5FUvVaR3uop0YO9chzxYfyiQhMbf
NWIUyiwf6bOQb5MjLkJVfj/zNgKdOzVyR74ZLc0e/qVadNZ9vzMHcGdatq9c1HIYL14s+xeBlxZ+
7kPzbC4EYwDICODlo4zd5NAqZLl5Ecie2+C7ZECGZZGXKi90prPWhM9wnRYCnavI6dL2sVASjvPU
5t09VPdKrriTbwHPZPd76xvhNp1llaqTW/GFajL99E1kA5hkWqgR4HBiO9F4n24XclAgtH7QSlvW
VA/nIfHOH3xUO7ZXfU6HNX8XpjdaydnKZ8XbaJOBoenkvITJLrZTvhSakKLHf4IsZCmY1T7mdlGd
REFPjhLTFxdcBcH6X5jhP5F7Q1IYLpPTThFUlHP/MAzOYOCccHpRN/vEKgnc2/bjBPZgnzPJZvqW
QCigrRNg8Vt7h5GWRNRaRZDPD+57Qmuwasg5hcv8zNnQnoUAWAzei4fe5KIQU3dh9M4JgWdNcHuP
pfDJ7u3IahWlMSm/4i2Hh8xdMZbs4tF+A3vrKvTRaT/HOSB3797UkCkDeK/XuPFbi8ccTBUNeoXi
n3BYku1HB+y91/5/Tn4pMGNzwTJZQG7SnYkVGnNnaiTnnhgNneIr5O9GdQIBm1duhDcKl4bmlFiL
EfYsm2j5ro1dHaF8Pn1LD+S+RF9wX2e6XAtqJ2R999zEeJrJkbkYpba2YKlObjeH9KzWFgBG5Ytk
E6UmC4rgyA0IlnNoaAvo5nB6JyWVsAizbZcxn81do8PFu4wadUo2LvFXRn/0kEuqfDP1YwfxJ3Ug
yC29p2iU82v4jVECyG+DXwm8eTaxPvssBCUfTt7hngf6OMqzUKcM+KcNZWsrTzv56NxojpR+llWp
NbURdRX9++JwskRWGFzDu2UasDhNxh9evskJVHc1Db0oY3nhe2opH2yvk8dqkrgBVnvYUTcRNufm
OpxA4u4ShoKfCbBgWv01X0tpeAPHq99nKLYPcNuQW3M6PP01pRltLVrrmBnI0jS+nMCqT/VuII0d
niPVeYLhh44OD741bvC9U2Ak2MSxMr5tZcCeuEHd9TcOUDrZ1MgVbdoKcUrQkiUFhnT9NjfM70hD
c9m4Kb81aTKm1lkOQeBn5hGeIhI0nXj8TA4R7TBt2o2l0gcMgDwegefKrPgnKC5se3B3Cp1Y00F5
tPt5fFH2d87ifwCErZFCEyrLIJK6DHhvYgbRsy7ua7VPDLh0qrHpxLC0T6IzuM0gxpMG3vCGzC0u
WkLTPTLUX/j6aiV7UDYw9C3AlXlE2+sQeWpfJCwhySWe+Hrd5yC+xGsNkf8uHp9EYwWhllhqNvY9
F+reXYzyDUqbxXe43eCP8P/BaEKgZDwbU1K9+d/VWweNk4UINaPfr53WZec/db0UpwDenAXQ5tkr
kfMcJYFbMkNRbsdlk+HnDTZ+L+wPrzS/5C2LTMGXer8eulhn1dmOXu3xxkvFkJYTbmyZAwZuJ4Wa
54e33s1L7Ra5QQU6Cgk3zjJ4xZppGWOPomv3eUo72Iw9m6mtAtzILAaAbGxMYyDdj00diBjU6tpN
/eeKXkyr0GPb/AKeBfuOw/rA5kmDw7KfaelXJvIvLP/muUzX0EZoWo2VVaPh1QNbOPJqlMGO8Te+
pNYDunWXMGb1lnKrt8uMl7PW3FC7un9mFQ5vbJSt5IqjtRic+tdjsHK+SkY7ZtfGxMixcskJOice
ZoEUFHNdLx8j5xlnR091dEnSc//gGKK08RQuL/08vwjRo3XR6+pr1XqN9Qsuhb5l4EgoLGC/vnWU
Z9b6YpnbabHr+bdRnSQwOmV7z67t1etmgl7BHmobW8frgNy0E5ggzWUh7GiD1sPqRFvZHQjIigrM
d1mTEEXZPX30uMeVBjsUjoz0cMkbrChZJCL/LwY60NBg29pX0w+ONyxZ13kYQNn901+AA8E6LfJM
Ik+QLi1Cep+gK3qYw6p7Fy35Mea9OrkjtajItEKRcjV3Q3FjrGbHpk+PCppvQH5ajOUt0V8N4z1/
mhR4wKJz2rbIpeliufuhh1G6PLHPceotjJ7LXSyf6xTLsoHBdg0TF3MDw25A+Ixd01Qrk6sONE1W
apszts2K80V0UFIUwtD02QlpJa9gvQNSEYqWb/k2E8c+vnKZ1aGdebi9dthh5RpDJts5nvWGUNsr
MgrkUPBwbH5Yuv+ideT4e/cg9QQVWF/9qtCqTUKWVaXLu1jMr6e1AsYmK7hdh24X3dqx1n6d52yQ
Q3eaEksAsyG29iDEYRPmMzZ8s+KHNQ4o8wjdenHmKazj1dh/FgteAUnVQYPTvZPeQej/qNRe/WHV
Bfb35EP+CazSt2DZgqeG6T15PbHqn5qg7VqEaPhUXwl5ihzlSnxg7jw82g7l0jyyV2fIkXc+W4Gr
xcUKwoet8/59nBF1ARbDNWLNYDWMafmuFFeKMeu5wKWSzQ4HYR4/1Zubumz/lTHbQy+e5fBzsl11
RCOlKY5x6RXn0jfLwYb8QK67xEBnTw/uY+4OChe74RmaUMuczHFhGBzByPWIlCTsnwIDvijqEKmz
Ji4e1EG6K7QmwfEJYReviKs7Yf+Mnp/AQmh6joL2bWjy7UXA3CUcvL/b6jp2vhlO1Fm/YM6rWEdY
41xZXAbfo+gyJCSiHOJK6YvPkupRQrOC1G/kQWMzY58IA81G5vBMfBVymVmZ+zVwWc5Z4B9vrYcZ
Eii6H7WqMaCagBEnc2CochsSIAO701BelGD4s82UNM3UMTjF6spUE9rf8ojb193bQTfOuT5UZ7Eb
0NvxKNTg9rSMHDR782oM/a2Ap4Mi4PzI+l/cnaPZO7/e3mEKGrIKr5n9v1S8rmIp5IjFYIiS2/zx
+r021XR4DzAYIp567+86xv+JjGCmcMpLvV+90omXtxdTLrGZ95/RvHk6xulXjlHZ4xsPfquMrGBF
FL2xeC8X0TdvP6pQLaesjifbNfu/KFq2Teb7EYEQs6+WyhnnhegEI2xnqEbOt7PW5sfYWEp4N1cm
cyx5FahH9TC97cHXG8DxXAozpDfjkr3spZ3HsdwVTVDGs7pmLkz66aKAeJpTXcgRvubFJnQ9CLKt
QvJL6p1FjQMfZDdDcKtpGbbm4Vq5jhduSKkMbTwjTfj+G/gw8v4UPq2odzpeskgpIR2NWsRHoZWR
bY7sd0lSyUkM0LJgMG7deEgktj3gj84PF3xI1VJFUoQCLEjygUauduxdul2/u+liYnhfbMBM2F8n
6eYq1wcojrD9AVwKVMKffP5aP4LC6ucY299qD5Hr4/RqilprUGBYhz1iE+cLYNG/53yivI3LMrAO
FVbyC/YJnR/eQtKljiZZNshEjO3tcq/kmYMjNVnOS8Ov2NJOVV0vqcIrtJ2gUFMQtZ7k23UtQF+x
fWYtNNVPrlesDhSB4RAmDb9YcS5H8l/DeUwzhkRZVAdUjEjo7b5tRzUt7D7I1zsB7CfXpFC4TWhc
GROOH+sJyoHQZGjbm/NmK63kcCNVeoBz1FYsDIXvVprkv8bsLjfHoDotYr6mpUtGvpH+ADJmBJ94
aWNJYYuEbDblwlk0wNrEz24HerMww5axh3QwKF2TLYNXcVzlRXg+SYXFdB8bmbHP2g6A4je3+bpW
a69iuApDi9sHacKbi9B0CTn/aENkYQlDNvAsZqMHG29/bMPkgLp1jwZYxmlUmDvm6UqS496uE9Fn
8l5kcBjXcuuGUBskI5FiXgGAmlEy8P4TfH0CO7scxxK10CmY50TeEVwmo9K4DuDFfrbBp2q72wR+
G8nLM9BRW5muUOmat/jGHnyxDVKg03qH7SmWgPC8WKjJ4SoXUtAIWqwMorA7KTIsCvCwQmLWBEVT
ycWkXlXdS/kKfy9sPdmt++mYi3/px2Wn3NT6rCEfjWjLYMCfw51sn2jYBSp/O9R+I/vjnvn6jR/h
X0ZpzrMj+GdEFSZTT8qxm4hI/0qv3UMJ8r+hHd1S6zirMca/Etyyy6WcIhoQ22OT/Oavs4CucfYm
6HE//PT7C0FSnXkLmrYOTHKsLmKuYmlo55uUPPYwsIJJwJlygbKHHY3Ycx9AGCxKRxh3O8FgtaiB
tXdOrJS3Hi7v+dXtyRFys+jrDgp5afaC6oFAVPKne0DX8Cp5UyNWKAjjXjUiwmwwxGirwbSghc/f
b5Gf+K5CpXYet4ImIBPK/9vyNecr3+9Ab6PBkXFbVbwy++AsQSiIa0gPfYIo3StLTfq78VRhZnAE
rHkQILgaBaqQl4YDrTLF+EnbBqikphpmGPP6Q6tlT9+S6HWdw83oQzjWsJUNyIEpIc+CdaPWF4q1
p8yjKHgvmy7Jd64HCAF1dVNXb8M8+vb8vXxIw/ybzWZYEzpiPhJg4MQOw+V3KURsAYoFkuIVcWgU
Eu8qHMHJ8eNQP+AaD7HunFu9lE8dHHvNj6+MVxe6Pk8/SOE3uO1uCrhjMwnUzV7uOogwxV8bNC/p
lbGN0bcEJhnSF6g4PwWAxYdUExeaGHACh+FnqzkTttUPz9Zw2GPbpbMF1HB4s8aCVyTLOUMtg5dv
ifU9ZXR7dBra7tv/CB6UV/xCkvtpd+qaYEbdSwUYGXs9CXGF3knzfVRyMv7Z4XYbzvyb7y4Dc9nG
DNrgJ4yAqdYOpb32wJw1/9vwMccev+n6ShLX2bLd+0nb5UhjLJssUSGl2ySd+oObfz7HH4PpU5xq
qRA3N3bxPMWu6Rl3Eq0UHC/kWr34MbIgLjj5nPlLZBXB9CcbU33vV9mlyHapEtbuqxhFbVyQMA3g
Ehe+CEpQcsPVNJEwO+9C4jB95mOOC0W+rC7toHxCHAsVdrFj90lUayQmMj/oTFB8VKpY4doz0NCN
K8baXieuz5+2L/OqSn820Z7JgE7P6gPgWbfp95vrKWixyTmAanYdY3nvpxUkWfNaCr2af+iYiNlE
04oWRLbLb5mCrV4DEGAE45w+pISSsz2fzonnDWFAD3l2xSW/nWZFSQ2+GsKjJZUWIfTGNZ5sAHFf
kcghGxp0C+YMx7R59g3EznZa5OrtXS8q/GZkMZQPB1hOGnhFh5MCH8iiE4lbO2Xn9zUFJ1wkTc9s
FwYjs+5G5+4ZKLuWnBSURu/dlNd66CvPhWdqRZKJjFc1RTVbQ9L/zw7FnXHjFi5DFmNYW5IaltXN
JN41SNGjxElTKxn8CByjMiBZwXaaCYMAXDUQJkWgb+yEHkTAKecD3T1X/ra06jXy+rZmtKRxgwlr
GFxm/5SZzk7uhSPvKUHe68v4wwJxX7MNlg+TtmRfIEbe0GbICPEu9OiQ7Hke+eunED10a5/TqkqJ
PnFbh/LRmcJhBWAPW/Cd829pHRzECcIHrdR9BiDtxtLzqo6HAD1Wy1JQml/DgEqXHiTVGcLiy68C
C5pY2egm6AnDVRbmzeq3CizFslL8l5vNLgFC9Kqjszb1OQtNNh+A5yshJV8b8vx+GOPk1l1+UGL8
/xHLyWdi541Y2Dq6wH0A2XofJIsPP2W3+eDIRuUuvJk/1SlYrW+YxUzs4fPE/RYyCOMCOSDbLy70
j1QXoAwntZLaeATfCQAOb0Ri5Z7GsjV0DVZKAisHUW+XMOGVt+2Jc+4gtAGsMurKViPEc2m8i4Ll
jUs6l4nBA0U/4LiwGtO9BcdI/XeBFDDx0YRZkf/P0j/5hOTGFPHllPacAWzLJTfYT5+UcBGGauQo
qT6Sx0Eqk5hS0RgZl7FaSoVL1OINxhCBodibthSzlEE/8FVbXVzhqeD5Lt/Sy6ibfAdcWMW1e2Oh
2doPhWujriMDuxY2B7z6x/lmbOojJVtyHRn+JUtn5piiaj3ixdtoASk9BsVvf0P4n0tGARpcNVbX
85fiFA0U8rXgmD5N7SkOjZML2pxeklEy0joDIPWloQcLTHHUeUAB/aEv0hG2zCkdVqfbY/fPToTQ
Pg4KQ0+UdlDNcYhAdpMs9W9FOCXgUQ917cyaPx1AoOtRTTfDM0BYxblPyUvxENfHAcFGYJtjsEmg
YnTuIk9rrG/BGdCDZyPE0yggpJAeq8P7J9VbW6jyvP9vMOHRVeV5O5BoOfJShROeaGIawT6kYrtP
Q/2qvI7iBajAtcgfGX5/fi/AM3yBtLELSBOiOXkrGnxVClXnF/ihn0fq3Gl44Z2EVgiPCDs7mljE
z8uTNoI9AeQ0SeYi3D2P2I4W+klh5PsLKQdbkDpq3vkmJ75CgG3ci72tBfsA1eZR/Q/RM2C+0flI
fX49IGPrj83Tn7bKCy4jjmVrYjzeBmtWIwnhIkMSbrKTIhtsgnSIUbssPqQNWzzMNBUMIVlSMfHc
KgvIAJIyHeLm2baR8dJCo3lDIE+dIo+VRuYV+8el6AiImgkrkHMy9OFqEEQteV2NfcReFge0o7DY
iffPAvpD9n0/qorxiPlSqQJo2Lfr/dTie4qukyoNZGGcfNMoZy7BbnSp25FEBugyJ2cc1Q8GR+Xk
JEApZtFRKwNR0fD3L/VHHAg7VZ/nJVLfOMNDorAHjnF4d3pq0sCFm2G0gwqDgN0fFnQ2S9z5lipO
zVZdaFaItnEgc36pCBhz02rGJuN9/qXjZdimCg0aTIeADjSDarJ9BdfAVJ3P7jlCeOSZPXRa8eLF
OgUr3U5l5bCJzLY8e8sKCcJgNHBnEIwMcnPPhJrcxIOSvUlFKx+FMFNDkn/xQTmWDbTp3b2bXAtV
qB4SL/UtzreX75KmiaiQF4OU5CcH3Yz++BWWF0kmzuGwDsVmkRy+GCIiNRx2Wd4XDKMGz8tBFVBz
rwnnqTgvKQ6Qu/iPUsi64I1bWegdDzLrZaDV/d4G0Sod/Y76e0lwpsbs7Y6COydrSJmqnY9CLS4V
8AqYltGJcAY8lVhmqU/JjvcaehYYWl2tAruFcOC0YV02ZTvWPojFyCrrhb9WRBxrkeIUh6uuZa/k
hIYcDGlTzgP82iYUAWGYTMsAbR0qvaLWL/5k/OhMAFCKoXkdhT6CXgLrooLbrtBobNgdmjn2chqQ
+dOk3l/Z+HBeQBXdwyUZMMVSvtLKw5ifsZtRgJiYdy8T4afyHzZc9jD9g8hqjVo8HeALjhF54UUa
bXDuKcscCMU0PreiGcqeRASgS4yUrbfcGpIoJ5L5JwTYspIfoXNdxD83F/8ZcJe9ojWvVO72hkVv
4l6z/QSSCGfu5M7qCnnaGtZpjqmOgkReEpmA1RtN1ZpwHtCJIYxqTK7k71v7MHGp2QwYgibHrRHp
19wVq4vDakMx7agSHDoT1C3P+wbyXOwOeVle2Yy+QYW63Nqa5ZT/cNmreqXgozyr5KzOaQPOSNpb
L2XRbIMlGTD0n8lIGDsSLldDYq4yZ+pvYGI1BnKiB7wNt3l8QjDp+TId6e5sqpsuDZUEbec1ZKh2
h6pT8U3UVE6GALZnZWn8ynpXsaS3AYLHVFHpYc0qqFvEfncXW4qfoanFpsMavGQO4xTog5gMLaJA
Z3h1nksm0bKd+eLu0Uf5jw5C33W5KcPsnyI7mRDr15ZQ+YjBaNcli5Gh7gyvXiOEx5h5cVrJ9vKN
HBIhHNnitDH3iwvC3vOb2k3H05/ie+bMG5akiemWMRwWqgde4lAr9XnozvIRtAMGAnjRVemsAoz7
ipwjHrziJrBE52KB8IgV6bW8z5LmQAr2tnI9+bD6aZ0oU6wJOBUwuA3nVlmvb8brWb4dso3Ah8q2
6p9MuHDXRDIOaajBRE9pRxMly4I96XM+PoCcZ7Txcl0HRv2EktMatAkkL3Xmdut+OazOUi5HfDYF
ngIwxtMU7cGThQzQEy0GRPCFDCDiOT6FkzgvVx2e2ZLhMDOiAGal1ijOB8hLPypL9NNEZRzl9WEC
tpNp8En0W2eDBxnYdV+avmnMlC1aNL42fbMyZhRL+yACx5YRhyqbtxt6ca7fB1j/mEeLkqa0hS+Q
eFl7ymQjIHLJeo4pDA8tLCrlHCO4kojmu6LkaZvVxMK4vBgPTxp7IlsglNIN3xwHbiD1cmDZuwZr
vR2bHf8H2Qa465bKpGZb5HlYJewSIBmh7XySEBuJvEJ66k3h0bt2wYBfF4KlntO2SXw3P35RLjU3
11gJJCP6284lfgzdE/95nV8eZnLCWNNp9B2QnDF+XayN6b/3jlxVHDbe4qg3EidyvWrhQRW/AWo3
mrW5aIsH65TAdTAI4gJLga02izybZlAmAJZ9yWgJO7VtttJO0KPokaxWxdvZ2Zi2qvVgvSo7BDMX
tGkVmwG2N397QtgEF31uCuYojoJhjE96WsCLYywz7sPUmrekVsr0evEOdsiac/ZI9DsrzHQouNY5
T/0eWnpKbdkeTYeUL/4cT9pS+sKslcVKjLRS0g/BO1LuZ//261aaW97iK5L/XQWDJtvxtuPMCNyo
ok6OmnHYyK6sBY7sWjoYXlOl6YiJehGWpwzWQGlld6c4ys9yEbRDZWEidwBDUvFGqkeIqyvU6Nth
ZRgKi39imfPKaZ6+PwWPPgX2MUuTeDCCfJ8OkONweaAaCzPKZ/kwK8/N+ILJ979aBuCW3Be4PSZp
A5UEDPOKUBgmMsymoh+JbVagHT6AHumDCafX4/vWP/ZVIM0DCEK1SbOtjgDnfV1AS/FahzAcmKe0
KgOrhOCKEAis+tUGRk8ONKFv/ozk7l0f284m9acqaX0FfZSzXsqGTtKKXQWrQYLhJeqtbbqHn0Lc
43T2zDgsU4cgs94G8pyZhOgc3OqbiEgEX3mJi9uK98Zok2Fe9x1zxKCYb3VZBHmfAbwKomCYva8Z
FXlV/MWsSghPW9rcrpnl4pbbXRwrn2DeofQ94G+jFLlmqFMj7oKeMEif+/C497LiuUtVa1MkXBzr
a2nSopIeqwvuBpw1T2Xx13BMJ3ZiP6+A6k4s8qxZK8xHb4yCQjtw8+Y1xB4iBsCs4f7lCwF25ghp
pHgwR6hKzibmOmxhjDuImMcNWD6yBqwMp6hJb1/Vl7f9u/ccPc7HUn9ClDxmPJS48TmmeijHqg6U
XP63TtosejyIFnIcmG2LVJoFf1lh9W25k6pj7Vdn7A43BycjFQUyc/nbqLkvgZB+jXXbhbon2IQy
PWIjVa4Dhj41I0tOqOKZ0nU+sayg7nd5ivobx+kfuOO0ED1acIH/jUYL+Iin1i7VNWyYg2UMIh/+
oGBbP9lL8fAsTVBC07l2GiAq1kxmFZLC0Igrf8q0N/e1PbV8Fkpaykkr3N/zl0XvPzUztVy1Eq2L
A7RUOTeFW3zseE97tLQbRiQnfy5amisTjJIeBG65dq3iDGQCii3OHz7fEQjH9DsQKUp1NIIczlsK
5uK7OM74QoIP4W2a45y/3ZVFbX92gB/oTxffiBR7ZNDDOVppQyZjJs5/JGU5KORIzaXUmkTzkQjY
ljNmBCRlT8AaQFWRcexU0FmW2exFcUlKnbuNrJaxnn6i65dPl1+NZ86UaJjcxrPVQLTo1Svyel3j
28AiIiRQLfyU2hPXmJs85kbwI/2G2pL9GYqwoIqtsYwLzDhD8f3/gwrQ9RkzVbe3j3bWjvVX1mz4
hvNMoSmoxqQjqgHUnuqA8m+ly9SJ5SxFmED4H52hnpS78xjlTCgrAw+QemQQTVmqIHod+E4Jqrsu
yxkHmeUBUxqdMzfCFJNXj/VxRqiTH8Hb8ftapLH0JuKve5SjXRg2LVml505u5OVhOATTckC5lEPd
OYud17PzqgdiKGtruUZlfDozeXZ2QtzHiZotp5lo1JqiNji9GhIjvpZv8E0b89sxl6i5eNZjbduE
B8s8iqwUgBI2LIzkpK3gUz3b1ZjYCl7vp0BAlLWzqNI/7xF7yjjki71r7rPAhh3w5b/K5LTlBVd1
/TAWmnwXSYSDewvc+FQTxqlt/xM4SjdCm4gYILvBNgqrlJVI9xNFASeqj8zS+rCc3gIHidqwsJS/
zrkM+BXwXVI6kDQ3ZnYlGsOj8B46aX1dYLzsO4XI1GtEzPz5saw3zlCekSBtHebm7z26BQn1aCjh
i5goa9asrO06qiZ4aT4L5xYDsVtfuJmrrFpTK1rNV+/9V3893EdHta3oqb+yAT/OHw0SjrfK06mV
8SSA9GNy+uXKyuYpwO0eMUdndVnmrgwahlqJEKtqk2wH3gnAexRqGW+rtoKdJcqszAUIQFWmcXej
iCd1X1TJrsN5Ia2Y/bY+LvD4NSU+DeGahH+jFAiJ4cQ983qYfi8b0pH2pm/CRnBkmt/+wWKlYPco
ToLvFZYmNImR1xTmblr9KVi2VzEH2oFN9+Htw58ICnHKrY8msQ6hI2rqjDURxbBcUF3fxEW/bKEH
NfOF3RSR1n7Ns/RIAj513fMwNoP2iqnuMj8s/P7TGNfI8f3tfN4UT81J+pv66dkPUYTj22CiKb6Z
30i2li6ne6DBebJJUkW51QOqsf0isdx3yFUW5EBJgETgrI1fCy+mU7vmXBWv4tuB3dyJH/Z0dL6u
I2KvL8cPZgvhvufaZHgiY27xy9nUVbwOULF/hs8+JwIH6bHjRZSPXD4QXYnvGO1FjfClc5CqNEi3
bYYztvGQHTWQfVqD4MmFIVnVzRdR7NYy/viaVp8ztbeFA9Aqfy1i7ErG9uMVe8cBUNAigacJ2OFl
4d92hsR/77uphRCLuIJY1eFOltTq/KUSpe2wMzxXjA/wSsyQBcos3SM3sdqJvhbIdVA3txtZ7kB5
FMfHQ8yngZ/wuhdbo4KrYiCrgwXsn2weyP3bTAa2qsMyHqgR2Yw/2U9eZVSPYtjwskPPmxmDv+WF
yWrOFDri77DYN05F5OfE1ttLIossCVUnfiostGrAk/H95AOo5alpVdVkpAxS3RDICRZm6Zxqfts8
edbMMBiQ32rKgcDY8g0cIGOyW6Ob1zWKsZCujhdmr1GIy0HiGHpIH2UAWVMpBz6I2Al0g01DalfL
TKs3my0wJVT6THbejt1ovMJjU5cVJhGFhr5PYkIFVtK12fw2uasNly4srRey3vjOTGmVvqf6UglR
0hNpkLX0i7UEIk/6QClJrYA7LMQJnJQlv3mB9RYkjYDsqCM5hY+eb64puSu8YEesLMW4LL1AgOBy
t7Q6RMcXoP3PHVJllp1Zc16g4eRNJ+TnD8PFuIvZICKeCTGPzxZ7agsKpVe/5OIUuDYfEEEtBePz
K99hrDY8z/iFullJTj+2GZqKXu1nR9/99lZ5rdHB41MvL19udn6b5f2CQr+53sglzuG3GpyzyTQH
ZkglyFUtcds61RHqzCWifMDiZxXQgij4kNz182vfpxJTNt/jYJDfLbYR/1RGTe/PHzhCDXgdFIqJ
/SvUGv/pIjW7zMhwWh/TezeQKXOiZ/ssJvTO8Ec0Q1sWNUvu78hOAPKcZ3dMFP8BmVAw7MFhXzVZ
V24Xav9rysoXAkVxowDBY3raeqPUsYdHHGLoC8J+lXYIiShETHkvSistGZbV1jqwKmT0hgx4FB4V
WYSFQ3y8hZikiUBJTJaFDUoeRXDimNvzcW+b+ArTh9VcfU3IH1Oq0JJJKioqwNROPLbCYRMgcylw
Vmhsl3KPZADrvppAKniY8440s6GAUt80tzVHDTXw3uFaiFNO6VKG5n0s15kb6uy0bz57mUDYHNZt
nOvhxkUs7n6622JS3lK4Jfy1FhSnP/19/Ro1jyRgt6OYYmPckF2QGHv/NA6dYZ6FR0/UyXgMPqEz
M+fNwHDt+ABZxn3uWXetlIJBkxs94Y/FngHyM669upcozbuyeZrpHVa6RrF9WtzACkfclmlTYiT0
ZONTKcODt92kcuYyfBmt2Q7UjuPdxNFaC+frNeMEEqnWPd5/RAPADkClGQCf4F/1PdJQygBgQCgB
2rnfJKnJgyrA9mD5Rymk6k6KndgUUtfetCP2+q0mj8xNBWZVWFcAcBoVJeJyhJH866qUJt33jSqY
9jpzJ1j0y2UaXEV3wdIDg8/zmG03Gby1KRcxXvSficVdyVBpBdwkL1VVOCSb+rBASuJSp2lx0NAg
+yBUneDNcHjScny8JYYF6az/YDGXKIv1sSHzrv1I1v0v+zAwofmc9SEQA4tpp5/S8Sd9j2z29due
Q6F8Lw3IOMd2edlJKJwj1PNHDqtWZhG6bZZVNAFUBfQ7QsM5IskoUMBTK1DqVa0jJw7rVxQBB4KZ
0MnMwjiDKjfsWBZlYb1XfbyNKSzYaZ0wq76qsNea+fCMZhxazVuyq8J5Cc/TwD+3LEI9RaAxhig0
Tzedl8AE/xVABOUYXKyHd7/L87UhIKbq40HxQZAu2OzCF7UKcP20yx2cz9HG48zXGmXeUvx+lm+b
G1o/xOVRaTibL7P0EYx7xQcxXy1/3pyyqw0NnQlhrgWCIcWCTzd8OvAqhaJ5fYtoLhEfAWY122Cy
h2OfbEjxK5PiVyKgLkyBeDvk0P+IVom3XF+36PbvcfWIuZZHPqMfgxgHeVnl4HQqNvebINUEzhI3
IDvrmREJDGscCNJEKN2JMlDsfbtt4vv+rejEEG5KYE7MJOM+cTpNXDZxGl2vtupue+hnUqqdU6Na
fDRv0umO8lWG1b4vUzWOaVrxigckD8VBJKTYWTuO+L42eIl5D01QIsowIhvbUwGy+ThWFVVpLodH
KuQJ+LmtlTg1DmvjGAZ4AVAWwmoyU/LkYYW1uPDGWTQ0yoS3H8T0Z0jbNpSqPapDCI8m14jryzJ5
wptww3dhhPHpyITIT3LoCjlEHdEjP4j/jZgmB2m3Zjf4AxhBJ4PRGoCFMk+a2bKf3ylVDMl0RByZ
RsqTRwAG4EqYK5LjlKHg7QLgDxmBaBTKLLCLa4qfBcoc5QRMIpivklaw0XUFujQQch2V7l6pWAkp
aM/jxZ8F1bvmz3ivq+NizF/AiBM799aql4n7rC2m874VoxSrAVy5QzmnxgIugP2AtJ9K5HCl2Clq
GV2ZxJk9zvfF7nx4PJ/60vn4a3hpRNL21vpeYMVKMWBe9mFgm0J2is0byNw/++ZGWUNo4wKcznTQ
l3PG9TqnRL4XDuRvTmB+OhYRU3fpWfhI7tr2qh4rAd1UedGPIRnzglP6f1TlHCAC4AkThD0PorDe
u2bMl2gKgQ7tY2cVqXYBNsHWdhQ+6tbFrn1CFU3nlBV4cxEBbrsYE2oALIKGjD+0JqMn+3KK1EyW
gtqX+5evKem1IUp3Rd3q9mTL4dOjBH0VBc2+nkH1wRU2/izXiis+z97PasdCEy7GYn3U1/aV916f
aLQ5z/LMXb0vqudX+/A8LB+CAht4jinvwYY3wpjA14FwMkKIH2r+upfGuHbgc8/58FFfZRI5IqiY
v+Ay2HIpbD1YXWQD8F7CPqQYn4u71Y+VId14rOzGRoI5mfQD5B8BKSMPNqATl9V4H/Pu4F8spnGy
9OmlrGFLSeIS/hixoZsF+SlollZQYjOVJNd2le2zlMNUKgaTCyO/tEZux8pwKOfRouJvmAnM0cSU
wT2mNGeFV0ok6suW4S5NnoJxB96XcVwOSwphLP/bM07pX3JJHDuder+F8YzSPp92g3zakFWcTJEl
A4n1NlR4igWGyE+SCUGZtfXplkl4SdKXgNNH9J7opMuTiSqKTQeVlpPZjWzB8ZXGqvy+Fr2pn5s4
iEMn+qno5KC3grZjxcRygwaQABM0iIX2NOWQJq9M5/9JBZleNBaJ8cWvbvswmC45Bge518mxcYXs
Llmj8deZbFlz4uNMDiNkCXHseTgKPgv6/pYBg+RPIqOfiskJV+HrW82VXo1OYMGGSdp2FRv4HxgW
PSLt9JL2J6AQbBRHAxW9rBAIxMpd/dXw8r64lXsWDpSXWr5w6+sxfNTIIsMh4FQ0MX6i1zOg2BWE
bm81Bh+V8dPF7E0pIfV2NXOe+9GwFwvrYQnwslz07dk8oUwh3ZSu5HXEZzNDRidkE1ZtiNsI9R6v
vxFRZrT551tqjGME1YvWb3HCjA5uickIdFwnj4d2+d09Sivnumwo0bxOe13A4/ZCnOG216z6ZiOR
QsEWh+mX5bUtj9KL99xsUOX/cLkce4F+w8gVY3X/EENmfJCW7f7Qr9xk9kedeYVRt17MycG/xIxn
dvNEc6Z1I4XJZEWT8M/NdeG4xRQr6E2bgxPVQ+1ih3vwoheMehmzh9Tzzoi2kxLc1iIangPWVkJe
Cu2NW/BlyErk96wpLVnS9JQqZ4NCR/JDu+W0/Toi6588R100NnXNDnW7peFhWVpM8go7ZoRakxQ0
8u8lK4dKEIdEBghdh8gCT7aX/sv5k8DP9zCkLpKamjiw4FIVj7FGBxoWWgA47oL2lCmY9N5SrDd/
4QEKjhspCPg5EgFIinyEac6jhmLmwbQN+Deo+UjAMYTWCmBXRdR2DthZPg2EL/XU+rfpVzl3OdA8
GOaQkiJ3esTbipvWCbqbdM7yUQ3Yhq1Y0ktfq4WKXCuDEM2QAkzff3U63lFfwB17lisj5l/lBNpn
7et9XoL05qsb++nAFhR0suBfQkIEAPXKO9hfmHwbkpw3q8C8ktM4J9c1GqKaJ3s++er4Y2pCDCy6
7wfzVF0woVcsonV4LJLhI9Dy4yw79QocBBdKBL0HE/oTxv7xmX5U8FJsycoEK9fTHjlJWpEULGf1
vDzCtiTjslrn4dtjjhtFQgYEnWf4LS1aIT9P90jGCu1RXiTM1jk9hRdGIYSy3Z+JG05BtjG28tcC
l79Oc64B7pUkzsiobIsKvoj0RmqM5YiaR5ioc0hinEFQR9vbCXmvhLgx+c8aVS0lcB9pixhE8ukI
/6ni/exgJ19/ZtQWoITHLS51w9ODtIwOkK2B2+do2xloW8PhaimH9zClMmmBiSU5H3AKB1wQOMpp
/pXg/uSbwMn6yPkt8m7GiT3KGqwUbaSbsh+OhI8RKaAUQ6XncyY6BMlvCCsu71WU2qN0udlXRS8d
Kqwy2t97FlsJrkK7Vya8Kr5tixv0MIQ6ofcopnMmaDrs2UQxDok701W7dmNjw6azKOOrl1SkP6jx
Jm8vUB3AWjHK7+dENceJJ6d4WlrGXDg1QzHDV4s7TL92EdUeyMBV6+K8n3WwqrmTmW9lwaBmKJKR
0QkdgHOKGpgUvKRNs4TiUOCzMZaofmRzTqWj36l/RVjeaUS6Eyzxu9sNZC6gtvgC0VGKaLvsMw4O
+/6o/2stDA96Tfyi1WcR23jR4DPBcAOlyPRMbJdr7rohS7Uwy7ON7LM7j1o4VpQVo2RZQcUXFBPX
cU8asa2mj5Ip/ImSutfddcaZlWYG3W+tDMHoZlr5CCyv/W+pqRvpQoO8BRmd23D+fEL/Qvt69j3P
ubidbyAy6KNoB01uCklnf80tmwBXDoK0xhb+DpyWOcDqhTXapmHMbHoWVrwrM9mc6a4mtlQGp5u1
XLB6kuAWd/PrZ/rV5HtHTHAYfxyTT7z2AJWtMSfzdK2cS8+cwcNVui/RA1mm5vCGbP2OqrGKzx4u
9NIoj38010KHJD/Zf1asKDm5uZrl33d/JsbykyS1K1boEAzBYlXZb29w0bzckNBC2xqGvxMZs3/X
+KGNgBrx75SVJTZROrQ9RM+ZE0ORq7uF/KhQW/p5kP0TZX47su8ntcGCKX+ROzUOKpn8zM97DNyx
MDatLuxs9/Mm28ghly3ByZT+nvp0wfhynnJioOCQfdHdyqFW0350xfWyPTiWdG3j8iGBvpOmJiO4
Dv0xRaIEGxLaXh3iceqgIioIGAA9J9Mv8DlobiZSmLYWntZzKmMrkUTThwIrgqR7aMUOjTItrWQM
LbdXkIL7ew9M7OaXi0qARaxSgNll7k4y8oDCmGXmak582BasJzWKNP4/MSBOS5eDaX7uIbWEfNAD
ARNb7zBCE/i+pl04BqgwsMl0J0QalajYzGWDSpADb36XbR/ceVrmO02WTJ5D0/r79WpHOwYSz+o1
6oNZIvOjf3Ai9gcZHTJ8YIontoDM8olxY+7McP/LbrwohQqhx9xlf+/Cv9VKzZ06dQx9gUnl305Q
ro3DEtoRYZwpbtYztcSNkH1WRU3HHEqaQuIX13GHdkhs2V0+QgXRWUKwA+bW7spZOrs5UNuQFPYk
Szec2IfbfP1HrjJYJWAG3KaqC1mV335lgSI3H7Rc/0zn4e2LHsJ5C1KWzxA+23HMldWUcUxW9Dsl
uoCbwcVlRTFuUAAdxtDimWFGSRPGSsV7vrCnQZJD/VLVI9DQJyaJp55kvA32yFmztpUWdZO0qyRP
t1u6Xh5UsXeeTe0n6F7r4oT2uA8lXG56EDmdjGGBn3VHSxdvVRt4uPRLORPwXZLQ14VlkU3SIi9O
k/1+LvtfmsbpaAbmosfjAUAoJqHtZE2kV54X/aAdQbnkKWJf4vRnKc/XxSBIf2y8lvPQENnQsqnY
weVfIDnTE8ecKM22HKtXq6KbT6U8GDRBCNNIDOv6HxI9tXHH6vSEaUp8I688VGyYH7RBz6mf28u6
i6PqGWW1ZCB8P23ZOiulI2wasyPTYVCtZ/W64CKQA+e5zEpOcbY4rKetKDjjwctojooTWlc2jw9Y
WMDIVNDWGC9gGdPseJNg64mTOao14pugvqXznyhjH13kaarGyse6ZxUs2TZSoq3Wd0t7lFUj5yp+
xr/5JGKkACLAv6vaAcRvcrXh6/q9l/EzQduTardKT1ODk2T1kqBNciHIOucv2uvK2uvxrZ5vDNDL
NVzJ4oyWNZrtEy2eXRYlqJRzq3qu64wTdW4XY65NfXanNmZNKIsUgh6AsUH2+GP8qIsiO8YQTOxa
CzJqFl+l/wYktzW+XKi+wA93TU8d/lEj+cZsz7UBuCF7lBuv0N2AE4Gm4XSJK2l0hkDQIkUSsqKM
WO4tnxyGrN0u2SV2p5YYd4bEeYMcQBLaGq2kpBvTbEeThRtEsFoXu7oUQ53TACoybwFUxDHynJrs
SpdjjhhWYhsq6rjSz5VFzaBobw2YAkfze9INKFYJ0kTBjVd85gnXswbQJT99O2wAYeJzJM70Yb+n
EQhqL3uIyPmlytLWzE1H9gUFnzYH1PB/pf2jOZl+TpSQ+/6R59n8qdLMsBNpjxh1WukUneGs8UtE
eDN4Jo/5F2cvg/t5lN+MR39ljRzLNYJjMQ3WTa3h/nBc5MUoIda3Bk1YGiMKW6ReaWkWbbHNcGOd
4j8oCauo3wEOeT5ddpF55doK4FpsERMt5wxIdHzZ+h91OmWVYovauHhHUcxM0+RWogVv84gmjf86
rz3jluuKQxOb64q3yHB96b2hm9eR2K8O4zuUEb4c4DwWKPQ8Xu3XXx9H10p+r6Ja/vbX3EhhLGvK
LRKI8OdSVBLlsrddVnqlBY+vJHmWzx+z5JwpEraKCv27NTYloUg/A4fClR6h8LjKTzYtWwFOjFK3
j2UbMcC9LaoKKbOJ0+/ejIDdvpXZdnPWD35MIcwDAnSSPXiM4frqSXvojA4+ZLOD3PpMQmXG9oJn
YPNbEKYqHFPO44O+8OxEhSTQOnP5aOoCnQk7J9kdLVwb+L5daoccWqqEF/1XolwnWQcCJ2dE3SOJ
aqkE7CuA54Jky9Lnh0gKOhgJiIfLt+hTFWGSGHuWUjxlwYFTkt3aJt4+tXGWnELUn97iNaFYeofz
PLaPbK1UABg1EDcUdBXwb/kT4O1039BDke9Xe1vLMRlI7E0lh0WDP+kyKOWfZkUDZyH8HyoBGNR1
quvxACoVwE+237hmw6RfKCefQ4/9DZaj0ARsLW6ATIdDPehfmLeNmwsrroR7ryaHbFIC+fM1Qk8r
BxCZd3ro6jSKWiCo4cR7XEo85QtNQDiN4O1KZmsK5e1zFYqTG8TzEIWUh+WJXqmGFJGjdpfrgB8X
3dZPpeLy/spAgHJow/VYOMd+AoxRHi3QhW+8/jI7ToL/PZR73bNiHHGABxYWmwNFrCyH2Kwlqtfm
+3pR9KA/sX0etyPOYmWlTTRaMx6H498aJa3bI3ujhRNCdG0srtkqGE7FJbQsP/vuHEDr6BFw1em3
gqMPcqMdaP2NRMB3z5266cLCzHPV9ct/KmFYbfBYYXVwW4bCgGGV3i5VpdODGF27OV5llgWuaHMp
OSjvLOodaYSEEW9WPVK5yD6KpeAqaFg6M36yr0bskvAQqBifXyEL6htsaRe7Tf+TZLI7DlQOsxnu
UTPEVgM2SVIJACialnEI0YwrcyH+Zwd2y3tfRSzqh5+Vcoe2ofpY7RVdu5FfiTOJDCkWS/q2UAdA
JzlCqSxHyWCkGNe7J3lQpMaKPoh3Yixq45KW4OSsqyvWarLXlSF1Fcg4h3YOzYkBqCE0Vu9jYsjS
Hf135DrtaYSr7quPMra6EUurqLoVnMeYpshMCBhuMVv+bAiz3Gl3T282N6Zqq/BjaWGpCZIRWS6k
R6nkFKDyhl3oEhMNTz7wS/h3hQ56lO5x+7cthBN44dcsJ9zT0jYMFqcN5cNM48kwX5RDmVSug88v
g62BNmkv83y+0yS5GlfglpOHnJQqIsnCIf8K6CAgKdKmc2VJkpetMYp5l3TaUEnRVwXyWTHTA0iK
qqn7db4v/lp6WkDAMiVIUi8UQjkE2thWz1gL3AuJ0LlI6v5rFkPFN9W9YUGs32Fiej1TciqTwkne
cfEeFcycWVEgY7K1gQ0+JzwkCefFg0Q/s3h0umTWo+cBheW28gON8roTr2wN0S25RqPC4DCAMHgs
cqNpoNz/1laNe6BFArMwhK/W6IHlXcLgcLwrVEHINBrnoB6MODf0hQTpHsM2bIg9J3ITpuUhgmGr
xpM+zCZq55CwDwwpM/5fg/G+hvAki2wqKKkFPk8DzWmpPy4P3HyyH/q8LiiAKQYtTnyOHYTjFs38
1ZUggx24MeiTSf2XdNQle8KV9xxCasKre+heXnM8uyXAI93xl7H7PeVwpNalardAK15tcTap+hHO
Tkp2czuEUcA2P/UqDOsMvCcNNge2kPaKBF8q2g/ft3GnCsNgBsX5/NLXFzZY4VaZYMN4VljoN4TR
9zUuklqRuzFrGsyKKPBBNi40pb44UwJmD8y36sBFueXY4NwPXaIycnyRLle38xqoNWB8JKfwvQW8
yXrJ7vq36TrHeZq7Zc9BD7xsucNAZ41EKzksbFxrD/vAPHbTibqrteys0a9THqL0nDf8ixorScob
Pg+hThM17Is0NhJVGYUdy4B7nxzS6HUR5weCZ9Ie/6JVH5+5H+hi2YmQxdYufDoggV85JkzbxnOh
kiBYhVgFBRDJDaG4s1ESCPz1msjIujM5SAf+/OPoRE9DD6bcOBDVhlDnLihMcP48iytnzWU9fckV
vAc+pD3BK6BixpjQXs0VoVCvSfqG/BNI/j7+p1Hw83QemA8C3xM4cq51al5Fv3CYzaXbO6an76ZJ
X1lDPQ/R65flTTHO9+tYNaBwPwa/td0IdNPBX8lVw83RQCilobZafQfRr6nsQbI9iNar4r/iV7Dk
Uq5l5t30/YF/fdIpM8aWZVIbTv/J2abjWqCKCSRs1+ssTGW1E3BlB+xMXCK9jghSfhlU/Ceflky/
K5ght16BnV2fXiTO8BLqliUMwaoi+Y+CfrgnzAttM0z8cmP9cfN81f58lkrdC/GOWjAQ+NqN3A1R
6cDkTqP9EZlOi+ShLkJYpldQSwD9k3f6uhwp0OwuxsH8VlsgfGGTPQ2mS2y6C29k1Ar+AS0Jhn19
l2+uYnDXNLQMgkTw1MA0//akjfIe8LUn3EOFkcUm4X88D/X5XjMUU1gBdE2x+5MgRKOU6smnLCCb
qSbkyI4Fn+w+8hWdbJkekSF1KzW4z3M4eNLdkbc9/3HP/jYSjF1neS1HSmCDyThgtfEJTpvSDIg8
6hrbp0cVvp0cUt1hcEhoacoY6n8xsSY1+ZKXxQPv2Zrb4krtj4IsQedPYs6YnLXCbWig6OsXUVbY
vB+sxB/1teU17QnaywnHYtPABs3kzERhRk5pt8CovDEbSXR0Tpn8i7uaJlOz90/EwDph2ASK2RYm
+foL8+PFljm7XzpAt2cOCTKOzi3wXiU+rASzFSMjknU9m/yzVbREGvkg3IYku2vQs1ydmeWyvGWP
QL51tST4jcP6vFpRx43vp48O89VlxivTaEGarU8NbdBNXqwtxCRNSo+MbBHuzN3VMkIivVWSKqb2
0Sx3lXM9gAwhdVEbwKcFg/o0mZVEAPSMem2cPhaAN8XCuMw0gX1P2uFDIP2j0DfzApdZAueKrdRt
MeljgV0WHb2qBCBdr7AT70Wa24Gr6pXQDvExngbZx6T9k4ZGKlESm+Bib9bLlzibHT6CP4pCLYWH
zpGSLaNk8zS/EhG+ZMJlybqDx8B4es7nG8Z0Ehn7tsvhr4S2aCMNRW2O6mTlx7l/oS8AuAaoYQIt
jXqRiOuQLva5vFnOtYyrjvqobFBi5kR+Wtki4bs9L+gFfn4Fp2gSSOm6x3Jn3k8c0vbVqZNlXtR1
Wqt4khK8sMwvn5hD5NOMlEhCuDEcPbHQd+n9iuLUkg1sj6tn299MqXaO3CKso4aOuS6LLeLrs59s
83hBLb3PBLI4LENsv/H2IHFhtNKJGvfcnY0aN678OpUEp4pNR946V/FQ2/dbF0QENCaVPyv3NGGg
RdHpMWmaPZV66uFfXm2zi/9B6PwIojzggpfVjBpG/fq/Re7suQvBCctptxpk2n8fpxmepPudJFpg
xZjL5B0/IYRhvnLQcM2euvk7zVWrHSz2L6JBF6tqod9C5QX3uhhbozIm3D1GGMpmtXg25hNeIHTC
fy+p4blKwwknuCJy77S5Z61u5Yk6UU6QVM6XVuhHpndYbwfd//rSu9sSL5qjZLzfEKsJmMVfBh68
eIyw3f859okXuXnd9Ux/Yx0lPtocFUlbAcxUV6bwGbyy0XFzKOVHjYhDMLQsXWp8HN8v0KhjJZYh
gwJR2ZF7uJBa+PebWWI/zKDFvQfqfolENfRanreUcnoHfGyFZKTnNJMQE0AWFKWxIGXc4zvX4h47
D09CpBslBV9D8KZXy9z5nrOwpeHzrBxrFsewNmNu8joOqNFN+Vqk9akWp65t1hOSnOVw4NZejY8+
Iuo35Vm9fi59pooGHp+mH7sY4tJFo3gLyjCWj86vl8CbDF3OoP15qUmj0Xtu/RLTi/+N5FcnC4k4
pcCPmxkKja23BKtmPmoSZZQ7ktQcvMnRRoihMsxSFGQiIlOYeBiJ0oa4U8V4fY6pflnJszINx14n
nUjl3LC344ueB6S2VAFeErNiE2bh9iX6CinSa0llE0OUdpLeh1APZHKJqjty7RgOuGbVU31WSO+w
M2QezbJIvUQVxOmUhyiZkXEC89vFSMFTjwk/LgUliYmDuNgy4ovPBw9poJz/iiNwIiRKq0dr4FlJ
KyjpgXYxeU2jGJq5LrBk4BzBg4TM/5axQWVxN13p+N1KGOi+w9vFCV5HRTWOo0lvkKBYxrqOdPzO
hT2UhIGA+jsIZOxrHr2XP/UcZimRTK7HvLezlzXsMERxOWMvn+Ix/p2Z2Y+TyaroZyfFKGvjwSzd
dsZ4Qj6oZZaSzTvemT0ylowv87cE/UpAVbk0GtXQpby46aOQRdIbrYXXFs2pikTxqOg1uo5tBduY
0r+6Vlhaigx8GMZn/N/oekye2ZomQIhgKJg6URBK6fr20vIFrpXiql0/J1czMu5IG7108cx92DUM
tpP1ZHPx9Ctep+oykQAX59/LYMb0SZQSuH0MahMM705sRH1Yt8xuVm3Z0VlPkwt43Mj8Tna2yyNA
mZxAjzwrIvyW/7fMJpmgEgPzdyau74KjlyIGyIhH4OjpSgzp/t2tpkjO+fySEtnCvAel57ylAYm1
AuaDTaU11/OpaWoNXl53Re/4AJU+iLCx2g02MB9VeRqtNSgWhqbEJBV9PhW0IbwYUgsqRCv+7oiG
+mBVfcDBY82rHXFA7WKcSwwlIuVMZtOPtH1aO5N0eFiGGhRKidkaX5kYUBpjn/w4dEwCuoBNpotU
cZiOUdsFF0JXjRvMa4LdWwqQl93YeVuSPJEVHRVZOA20MEF2OA07eb+zmpveRvww5O7/5g7CtfVq
D4qRaa/c6OOf1tRqyvYh+C6TnTcMma8nPGCaz3x5Djz0frWS0bSmvxvDb7Qu2oA7LIhTKGpbF63u
JyhYvh2hRNk57ciwUvnceza/XUGkX8H0dTqnrUns0IgyToTTpb0fQK5pXsId+C7jKdSv/B6IDyQ+
amLrIr7nibLvkiIHCdoSprcJHZ3B1s0Mq5r/PBv2dKmUtA8hl/Lpx+w+3cF+FoV6IH4FmoUtrhn1
PCtJKMQQjQq1YBApFKHM6aTHR6oWcjZHI+mX61f1HT2ljF+3hKKsqD07WTsMFz268krDJYKRx0/1
YTIaz90P+aujgBR55lCXmaZouU+526IeRRh/TzI367h0cHyTYoYXZUt+TAAewRskiIPHjJT4pUlF
ASKhMEl3O00fo+bVTMkn88CoXMdiFNDj00PxnJYeLnX1+JpK0vJTtzzOfgWyJct4rdLWPn22nLV8
8Qj30tzvmjzlWG2Rx4hQF1RetTq+gpCTgVP0YjBeWu3F/Bl9AmV3+Xjq2Y0ba/x/CXRdjpEnQRq7
IkHqgPIhPrE5DSWEcig0GtotdXIyIsD6gAgH3mo7cpkkN5lYPMtg15M+TCZlc+o9syjLbYKCbTVo
D/nrDfAZB+j5IFBfPPyD0mSexvl1+xbYXdpF4HKakDFKbEBMJT0nsKV6qIpXx23u81C6MxkyqNWK
H/68dHAS+3gm+GXQ3m2hXN00gSRQgQ22/kbim0evxtPFIIIjUazPNrxOHM+AJ3kCVdzsV8FE/ET8
s4jwPfaA6A3gl0NOcJP+TvFIspetenROXCB5EpiFwnx++rOvsnD2WSyg8GbI5LJ2Kp/6LXzc1mYh
baXEgW+fmrLcQoWVL0CMkvCv/15PjitJcaPhV0iUpx2pvIDjqm3sJ26/fEJUym6cwFdHKy4svb7g
D6PSS7AYqpZY/zbsmAFKIYGPpOjUVNcjDbanswWSCNqJlYg5cdzFM9TLecJKsg9qDJpcIWvygLGV
AWV3ynAQZ7WeVDaLss10xFepq/x7BKjQDn5oH9f1EsvxcG20wVq8i5OYq03TTQZHPG0G8y+kIOwy
YEKoqVB6JboF5HnyhgQiuYFAP6IqDETkhgGI8GX1Aqp+9GqQM1gZp5kcHCmJOdTH5GQJcrzQCchk
YHJU7Tmpw+bF9WSOqrPrY6ZHqsH4kILEYQDZsjJjQWJV5GhsWDlFPX3Lc5jl1c12MoJZ+J1ezbJH
himEcq9D+UYJ64ySxkBcoB7nBPe3cGSlQKa60heHLJvukiKW/7nH7DMzsxbQwf+6a8FK2w7xVPKX
koHilAIsU51OM5KxynQYVtW/0jhnProKO0mlm9a0TrjPOu5by/AJTgUQMpsjZg6cYzu3rkNxuZrX
KmNougUL/H2sOPpcj7iAqSpqMiayT03xO4M8n4nEQO+rbFdRr+DxenyJOQ+4PgXPfb5UX3Nof7hs
UUEtsoMYDnAbhobEA6j2O7V/uCzvSi3FU3zVhfaGZ8Tibk2OAJShp9lPUaFSVtXLNxNJHXA3C1RG
SlodfJCtDKxkhIPj4p4b9gGcLLdB8p9pm2LCOZWZrJGcoDjv9yGNSym3GxarnqjDXzbPCxL17vrX
wy99eJvc60QABQS5EyWxRYPO0hVd1BKF0efg/ef7Q50XkhdhtZ4ZQruX8eHiMh6CPEwp2a1Yxk1S
GXkA8tcfxKBMoBGvNaWEOigoRk1QY+09+L7aAKx+Kls7JeQq4JLcyA+sZ3ia42zNVvVPw7UJz4MT
hS4RHVAAM4yb8BHZa+CVdSeIXT06gqeXZRu/R0kcuJPjmAF5KS2B/B5MmG/eoGV4L8wC8vPIPbm+
1CsKPpmtwzhtQ3vl2++HlxhAw1P8pRJXwKSPWdDmeHOa4rAghNEFnHuFTjabfTZOBvaBSQcYztzK
0BXKu+Md8LU9me4mZCLsALQA16fisZmUHY77YCS6Zoi1zc5QGFEVQcQZ6/pm7L2R8ziQclgLWisy
XhS/lapKM17YuR+ezyziQGWJqxw829TjSEqxkL6l5Wwipx4chk/J3zrMgojA299WNlE13GvSFbxS
oEs0QDVxFBM6csnoZz6TaLJo9BM2H6qzXqQnZot4xV48NgEg6CgrAs3Pe0vVEPwqL11im57Bx/Ru
O62z9qstfD8eMrfjdllaj77Ss6SKgy/hYgXQh/3RIzMILAUUnnVK3vSr9v8ToB+o2nVvDq+Ulzmm
2trp3amvZMvlSTvXj9KAogzBGClUS5Qm+MdF/87MjsiTDu+ZGIranQB2oVD0K4wALKcP9oQB4zo+
pDG3BPAcfy0jw/c0zbjyWEdeUGKyoKdFpGaVjHI+w9GDpj7NEfQHgopId+0oK2goC5JmYkB5lqv1
mZGBuwgxzynwEBwpyxGsE8dM8BOT7tqS3bj8hM2csGLPqXO2YS8OzlGNAUzlS9K0ktqCtzRnfJ1Z
Ojj8MXSPZkZji5vzj1pvsHorKWeteoriMjOiQMTTsBMbl9vVbXxpIlouhp79AF/sMWra8FJ5hxRj
QvEVQtUOMbClfo3TsXap5Wrwiljlh4+XXf9RUIifeH1y9dGFTT+6Eyt/e+cI/v2qvh6AsZfeZA+R
uw9tRz0tm7JeADsneh+4IWxzF6jY5yHfH3Xh4sVsudDlFN7El3mFitHj9liKiSvgiErmg4d5T8T4
fBw7cWSvM8kV4RSb6H1d2NCvnPe1sbBJAMuFQs5V3yKgXpNXFC1qORJVW+JuGIKCKR/nwxT8YsHJ
pdy7ZqIpmCdWGJfXhuN7fpAm3incb7t1nKAf21kPlm3Duf9dJPp3rHI+rVvyTj5c3gxdSdKaJopF
Ux5y3lbvHNmbVN4wlO/IOfi1ceSMFmJ5TEK0pNi5lgMbS3YLSqxNTp7RdfQbEDhrZFVKS5Zv4DwG
0clG96lRtBkX8CmKLx71bKDXihfSvxdarLwJibR8DuKkQn53Ho4j0GPTNVGrqTzybNivc1CCJr/4
2WOqt+ouZDOVVwHwCo5YWLlt2B243z3eitp79G6JiRT14T9YlebZtYhzH90set5qC9Mur+LStOed
zFMvQcXmNhBUukJGg881rDGgw7sbYGIXiuBSHvxA4bqX02MAw/+soGl6MXxNKJk105FHwC/aa01n
3qSDm0LVu1h5EAbBZj8y/Q0S3h08OlEnQUS3ONwkbQ7QO/RkXOUHWB7M9BNA2kWjOZxWvwcXjY0t
HaWS/IqHKeBxXcskDJAErb/JgiI+hVbZaJrQsnYSEhbvnzBlgaRdD6EMYInq2ks5QlRD3QWfki/f
582LL54PipbOv5v0VbI6d+TpZyWeKYxekg/15BCSr0yzavXWWDOv5+nilYDdUHY1voTRCGU5z+ER
M8qkC1WnuZEHlpHvYE7tZpGcF7T338wSTrekg8H582TrEnBaOg9+dEDcUOPqWS/J++yCJ7uyKtMs
DnXp4gMQHDTdtQjsjl0Mn1AueEpUVuCqxPVpJ9SnI/MBc/BD8VaqXyhL/sU1/2QJlIwfJD6EOMBY
uKJBFmT7tNc7yvrHn6mowpyV6f/1KL3yS6xIclfHmeCbpnlAhfqibbV2s4uaZ7ve4/19r1ud4AQn
paJtfoTdgosl3vkfKK3a64IfwPqYXXIoIjnOJcEuYN0hH1j1aUDndL1pQFrdPaJ2+UGuW1ZQ8nfF
sM6t7ZyhPXegyC3MCSbxOQH/0tnutbUNGg7EptDRZbypy+dTucM6GbCPs+/m9Zn3NS9AYTCTTnGW
dcWdW5QkCWx5SefhFJPrBJQJnDV9zG2yoaiisIEki/fKlIKNuIrmmQS3a9njUdb6xsw6zRRkdi+F
fum0gjLrgzZdIS9VFLj1hhqq8HiEw1x7KFOrVBTAQq1e51Y/CZ0Tng14Y6BVkuGbhmcTKjAzK7HX
13vMS9gSp/8jrRELuxl2k7id3wE+av/61ZrvigM1UofrJwX9UupELJ0cKFDKbHkl5lu7jnX3DcJh
2cffVjvH/CVyP4EWmf/OXHn/qZ1HC0xGOVo3ysRUwYcT+vVJjmal7wsU0CBF2TzbJCWKX6bVzsq7
MyKBLOC2V11CEaDZVOeqQJEy0QfJ5q+2cTWtyMy+5X7SbTPtTDHDx/fT/BT3Cw4TQv4uX9mnxgbO
X5Is/0fM14uifYHh275kek89AbQLh8saMelRskrBVievAeM+4LpIRxy4kIotlKj7s7o4Y98LyjcT
oYE7ssvzCrAvQ+QhfeiH5NJek8rYo+Q3YRebMIYzYTWveJ0c3ZXHm/F3GxZgQ5dbDDM9l/xtiXC+
aakoR6xjb1kU7naPSowV3ZSQvbaYkfPeV1boa/y9HEVbLCLzNOZowwYrjE57Ef8D9cb+vNzbsNas
AtV/FvDIld7nRIB7d+ITrdTWgeHrvM3uVM9osrsbXJThKKz7ifpkbr/uURVthMgOhi2nhnMERvCK
rd8mgn8XoyTbuc0EfWhPDeyTwoSYNKvkNFAz9b2Nm+oo9VghmzsllvSNTqh6td5s90YwB+MmieKe
HhhzY61VeZn8sl7UbNw52acEZZi0hkIZdj/QEJyuQcQkhXT1/BXMPQAG/fGgCzgubmKXdFhPmKP1
dH9f5EvBgG1aPgPBEhqcPWU+JU/JFfYm23UWyxxmOHvOht9QwUhoUKQzS0rTC2aYdBZmVzXhK/k7
sMuocTWHHGH/hGr8ocVq3BTloFUKuAYCwJgdKxbKKQCw3hBH1wIGStTzNMySM2PAp7uTjmH1sF3k
zeIK8XjSJ3rEWenQVw50g/G+ppdVnngQcXkwY0+zjjeYy9uUNHeQHIrc3BqMiuqO2Wvc5c40U6vW
LMNmpKI6gRwGi+TLPOjqhekqPlZVD2GSNUG1iNrcuuRgZUmbCATxwcwIPJCw+jNXdMnhuGQUmrcR
FjOdxlaZXAKdW92QY22Xfig4HwsLe6W1qLtBPD15Sv+DGKTd79e4sPLicoRUkUem0rRwETOdSaRr
ysHhbtEntMpT9D4XicAsRdmvCTOqWTf1oJOf3VLDMYVfZdCGHFgagXOoJ/TKZ9R+1wBqcbVDGgU1
mlyDkhmvNkx7wFB/6H3RVbX1o3y7uj7lA8NNt/KOH2cd/0lYguc7HxoURIcf5frbX/ZBC3ZjE3qt
tX98TLNUEfKFxZemX/gFiEJhzOh7njZZqgYhZm5ZaFhiArvT+X5eoxxIf3RYtMYGhTcmp06OdM1H
eduvFHj30tJagZ9EpTGVzejKP431wsd00xunn/W8vd4mbJBuIF8TMSdEYXtl+/AwbNl6nz/zeBbg
wb0QNghxKbEOWgzSONqZ389Jn2HZV+WTjdJhwLCyR/nJCFQYO7TXJ3PcNZkhoE5Wzr5261LN8rro
El9P1PqKOXM+N2n0DOL9lnU/Vx9VOXFjZ2TOw3r5xLASCAJaWQ8yfOjbEa2iyRWjKxORrqTRGOw8
2svnyH0cocUIdddmBOix5tr72NZ5HgitJ+Bamg+nJjDXR8wzLUyW12Dz5RiwxvCuxRBvWTZQAVgM
8wkco1lhLBAKogu1GlqrIfrj0LoRhvRHWYVI2XXQPjT2qQUrUj5KcHVY77U2QlE15nAl63r9LxBi
uaioR090gBKykcK1SknTRiikTbpWeqbHgQrcT/5aPr3eSsgMGl7i+YCY/T8Y1AyltVToVlXnkHLh
h+RA4BzpX/9kputaT+YCxDWL9KG7bAB0OBocI3eWecnGvBkJV/a0LdKuH/Z0DkVavR3PKarYktl/
4s5cNtopoSCmo/I2iYIdc/PjoERCW7xCTiLDdDthuGahPzO5X98zSd/mnDqpF8tDfWMqh76Qhm2d
h0fggPCSQOIboeZferxYEblAl2dgxEe2HGZvysyqdlIMBkYKXPFRN6lWKC9YlOM73TYVcrGscAdJ
j77nDqRr2YpT6r71/NkuPH+b5g6l59EATVlxFZlgdHCNKYLKiFi5UMMhiSSVFSWu44YxUgdfV/mH
gQ+1L5e+vCJZe5jhQwXoM8ulF3bz9Jid86QaSwwVXco8yvBANPaXBFBpPYrgzSfSDHSRcisBZ+Ov
9uTxKl8lLZ1K9ETKgqv0RbuI4Bzi/fufiwyUCvQVL7G8neQikIuY1NIgW3tozIBln3d0PnYj60Ed
pMq5McDUGvCMLWI2Ecq2YSBjIU1cAH7u5gFTYeMt8/ymqIsSrkAQXCI7aHLjeYBthwl/cF2GBEuG
YrWWT3xnJYPW3HoMv191XImymcZTGzkGM1Jc7UzMA9ZiPK6b+DHMhDVumf9BEhvcADccVYRgAo0q
EejLPEEfjoOpSJZPCrDTPflPEY3SfEjbAklFsCY0bSiw/Msl3eKoy3PudWN614PFpjZYaQp3vZw1
cxyelU8vrk/C/sNbdrZpn5DkCKL564zUnBk6y4KMRl6Li7+hTyYFGJaFKhplU3l13sJtRwQk+QTT
BYJZgdUwXp8XjowFKEU+g4KktpB3yoB+DMkPrLJpLAxOwITjA7Hmf5IvqikGMOP+JtIC+GYJTHIz
tdoenrCbSHUVOR010PMM2yrrBzZOIPN7WY7CPlEn2JqQy48Temhp4fW19rHGjIczCVf2bTAlnp58
imv/HVJPAOZYNxtipxMIqQQionCRxQZaxID8L1izgvnY7TVOyIDPEEik5RKz0e8gPQjIgvmnkB2i
qlYdgEDJzhmvjbUZEIvOjUkFYE5vv66thmYwdV/BALM/2ZkLabiIzWURf9qeSMzVXamp5fVevSEQ
bUj+gWul5ujYCAjPLcxGQ/YUXKsJsTm26yDhGVwGyGKvzn3e3cU25xXtghOb8cfqs0WVFO/wWuct
9YGXf4zM7brL7DIDAkyNdOS/27dT3r82Ihf0WEEiCN9P3j25QguuAbGsuyOqYURjsttJWjYzH80d
BPOUOJlES7k7a7RwT4uezgvnup7qx43gZ+6bqujhXwllyoYutCAg/9Nc56Yr6rGlLMAJ+L2qVp6t
jK2zHx6fqCqrEQrO8DnBA16DPYCZIqxTleFTy7qDo8RaNtERUuqkOOdep9g4DSgHXb6GIo86TjII
Lxv6QuHwxySFu5qzBhKsoVMm1iZsgAxSHYwn9C+hfgiLO9N8MDetsO1skVCLx6kNb3gXVc2M8+yy
nhYbKhDsvO4FrByZmoW/4yLv1TeVLx2pR1NyEkB0x5JXpRetG6afK565pb1TMi5bhzE2Jpd2N3ls
OoHUTXkOIf/PmwWTjJsGtjmv/4SUfICDpExBEr3B+mhM3eEFZ51pUIufB08xK6gKzlcDXc2EItMG
UF5O2Af77UoKJBvqqMc0VZ0B3eepf4E9KYUrAlnGLQfTeG62zdg37UfNuLpNdsbqpR+Y2/n7y32r
+tK+b1b2BJSm4LlpquObSU3pV9/V+oHrFBmw/oA3bjVaeBOpkepGkls5fq+6TDWb71AYUMHxyfIG
PBPIox0XidzA9RyOqxhpSWTes4Cie/VNccwjBFrMQhrx+HEEX/AlM+VW8aDBf8sKHQQ2SmjeAZNk
ZoYwNWIgkj/HpK+q9I2O6TeRjN/voLCoS+9hYlSowQXeJFKCxFefytcrY6WzacD2t+EXYedB0j1j
SLdZRqNqgCYMjVWVFg5HJ2SNcbgbIJI8Gk8eoWi9tJoA9b0ovMeGxOb2jIT8gSotfXbaYfrj6Rya
1ujVlHJA0ErYHwWjt5Cu+7gUpqlxCmXcBEYPoWb6xzd8hOCOkrC/eB0Gpu6+7agmmB256QUgq6c3
YlRlgPg9s+il0c7z2mKuQa9px9/nqABNlTvpQMnCfz4ELtMxg5KrhUgBpBsix7J7tfFbQRYtS9q5
e2AyCagP5yq3pg+UdWXUXtfxZva2rZeVj3GkdcnUTJfkBQOX09Vebp1/JE7rgaqos7a15pu7cVPt
/MJIAK5EHB4xqigJmi0H6z19m+4Y9BPDWI/6HmxZQhI2i+dyGRcntZMUVSZmylLQOBilQhbHK/e6
jA2E8/XH3a6tN8vRPl0ZiDbQ1jMLnDXZrWU1OyIN0FaWQmj6xzzd5QbiWVDA0z9C6QZsvr8f4ptS
fIcX2HOeWMRwxilq9t25N90PHX3BAmH/tvchH4qBH/hPa8XCjsSlLDPO00jkiZD2vU7f3E4855pD
ZTsTtGGwLoWlWYZfYOSaSkgbaVl3VJLs/BSbOWOfoNf6/g+tWZ9lUdqVOborN/jNS3VXee2pHMZF
LEFOWctDoui/eCDoAFokh8+QZmZb+Uafk/L/4vUPoVwFTZFnoouBPbTvdocZA599MCBceeo6/Zeg
jS57yJ/6JLkrcpyq+3Ntk9J9uHNDLPrvM8cZ9urTqIEr5jI23olANmord176GeiwvCwUk1hhlNxp
TnpRe+XSYvDYZLotbGFSX0VNEt9fc4Z9o0FUt7pIVmwFQ4XzDlr0QReSWrGqJxH1YnrcqTV0Cdsp
K+5k3hHJj7L92iA6D6ywvZNI2+WBUT63PXWC14hQ9SCZ73Gbsxch+wr3w4pdWjTrrkjbHdm+ZL0I
9KGqDRp6zOnx88E9qJF++FkOO67iNzFz0YQSKXeXmlbuCCXA5O3nMvylyglKmEGih3kKwnoIbSAu
5eMgtYBEsTSGF3NB/zn/16p3gRzesgIebqaImHQ/joSP/b7AZoCasK9DXIXx55ax8GDPdzPApNGv
kL/8zs+Zq1sfAEo/e7veXNB8pMiMSsxT0uDTnTri3T+ewtDBqyB6HwS5zYhb7Jm+aaHI9U1ETykK
ryiTIlKGSK9IX9etIw68rgLUeSnTXN8srVWh1x/Y54JbE3RpZNb5pTrmj+kKrA18y1UB76fFO5bC
G+akNqXxPuDXtoqiHMmUW+6rOXbQTn8fOeEpDQOFNJWqWC4R0kCE3ekVEGVmVX78tcUIJU9hLEqj
jIeP9b8shgoun30u7Tq8Oa4CFN5jdtZ4nTb2jQcciRUS54kq5Xlya2qB5CkyYkxywVKHEf77/P+I
UPTHdIlshbmPl3njdYiCAKgyU4hFMOLvCaGqiivWZqiNtdnx0tP9HNj003Cv56oz6W75Fg6JzaoV
V0vMdIEN9JikxsGxwE5PeWgVf4W5As0VKyEw9N9r7AucJ360dRpKRg4jNrXtm/pLP0rAviK9/6Fm
i7/JLaBt55CgNc45GfklwdDWFIXS9K63YU7OwpZoQ0vQJ7qii/tut2JK2urUru2HDQ+x65kUPMao
TWnl32YAe2AmSGiGbowsuDtlSNJk++DrntwV5OkMZ1GhiDLbOqqdFTY53sgwJAP+cHBmKmKM148l
X1DmM6dX5XAw1ETPaoF9vIvVizDF3BkzuUNmQb6f79r+Apmf/Ov4/R8OBNLlUvl7Bk8k7nXrGzxO
RtL1LHGiQPGRhiZFTn+qagKLv0u5BZdSNMEozQrl8vuaj8tOZrOY4rQGpc56A/mMCO4zTFnfleFj
launzvgQhTrdryBz1pzIX/Nmdou4P42JnRhzJoRg3B7qh2r3QN6X/VCQoizbTDlRLNx03i/G0ZuN
dJbRaci0ibAhp0/Pn44yEADcn0Q/0CnjGVNMq8JOYn4TdxMvbp/VDV5pIi2ls9mGEOrklOWV+Hhc
IbCcqZxHyRcapWZ/rkXlmpWGLnpHgJDXH+RSNFYOLPJqGtM8pmH+KDMP4r6zluf6LT9DMfrQ+LqJ
fg34yamwt7mworUUT7yrckdiUIhXjysh2i8c1+9+l9lVSf0l3ik6qqO2/f1xYwMfz930qwLs1BJb
wdnV5S+6Qj40k4nbEv9UisBpGEQdd4ilk5LAPVQ+MrFYfapDQrTOsvHMY2P5h/3CL9F2LG3JDA0I
IiLHY1LwJE+BrKdUtK88N/7KtzqEJvYbVgy35XQenbkgQTVF+cCXoOIjVxMbltodtThOnHmnAROM
EFzgXdspPQ1vYJhC+g57GqVuSx6pnBdC49Ywc4vgFUS7J9DPtGllx3leni5UTPRH47tKaheR0LpE
EmJjudM5tN2zyKturE0agEqTmddqWxlFHApryv+0YHGgLX/Lfnv8mMF8TZuYqt8SgaNIbPyTpini
aM+KiPJld+sckClrGdCpcx73JTEYH6WiBVCvJi2qe3bTsy1Eht9B22jTFmnxEjvejHeBPh9LLHCN
Taxibta2+bhjniLwn+qHMt58UZddjFmJyWblG4GY2JldlZJJnjPxzelb+mytIGCKIOjOk7IEFQpI
/Bf/S4gkb6kCpCqKi82ujUvRj1Fm7RexYOniJOcnDxAi8Fk+7g2OLLdWY+QQrvmYktaevOADYxmB
5+0rCD4IilXh4Zkd4rWpbUrINufQDKdSeWxA6IXVN6wCYp8HXDN3tZzL1WFDAtjQWkMpfJapVghC
84rKol77RHeHz2n8XgecDMfnFjv5v//yWLMAyfJqULx3DGi6DfiydP1wGkNNooOiN9+TiZxe7Wkj
g7+s/lcoQafn7Ijo+qr4WrfL9m6+XTBTfBikNEHL9FrFw0P4jn3P12wKuj4/aKUR8RZ3o8zQMEM5
SB3qtKp5cT9qzFrIq5HuaPDa730IZbUTRhV37CyuTLDfFwQF1EaeLGpDwLtIEgEFIkAIP1DTo5so
gOzEzIIZRB8PI5FcQ9OE5F6bw+CjlB0lnZmU7comZMFhTkj1tNS/zEWjOIfBshGgfEjfotKDp1S6
hLybZL4LhRYrKgxpfs4RsENLmfkWwBTmK13l06oHwsmYSj/sFPCvGTYRFaF43au5UF0DKWG7eSYJ
c7+05Ed/zchcWV+53KxXN4ZkIcdZdHLJOS/DmlAQhvLo+GwvP6c29mAdnWzxWuHeKTHhVqZtfXUd
x/S0HfpnKXb9l9yc8kxdF8NsGB8SzoUhH03KndBdqrIZCy3GgkTXHz/F/zwXZ1ZYr6Wcb9OMsAM2
X6qhHamd6Yb85OWU6zvljGO6CFohDSVUrCx4uS2HiMWG3aXsVtyPRfBDgNyYw9BUj0xAtj25tnoV
FjyTTLwfFaP2lJAuOGp8JKQain0b13V5HeU9p2j0vHmoBlpCylJjApF+AUw9lZp0Q+d4EHdngtx3
k/UGipTyqLIETyM9jhpipRu00nr4MtKujjq2QUm4HlXb3ZbpzdqLcy7hjqsEngnMifCxy0xLTARP
xrl9qb8KYKrfyDJNsmYu3OUtp7BFhNz3JIQZ7xxYo9CwMK+Ihe8Tjzq5LUWo8mADWqI+34y4KVnH
7p8d1XWv/D8v/jFim5dMoQkD85MMP6/xlWLIqrh3pPCmMDTbZ4OZNGhOHQphgKP1YcPjMwjiupDj
Ybb6B/iA+Icm6DatK3j3/dWc3ervwzYHeVTFhzmtAG53z7oK+5FKvb7lw2lItN7+AK3Y9IYnCp87
+jfx4LX7c8A1ignbnpqRmmKcJgzZPXjJO709BZJFUDpO7YCJTkJZPW4eR8YNQdWDCg5qtCxwFTXt
a9RxZSrBsZ70EWqACVSwmFyRnBKZXpu+WJr76nkrlMuf3fLGAiLv9BGrxH/TvcdGnrrefm00TnVR
6p7IqVugYelv3/YZ6buk8uO4Fl+lzUXS2Uy44IImcioEw7868OdTvpPpP21C1ZvzC01L5Zh6HqeB
56nRQQhuAbgm1namXPboANKhIrlDa3mbnfIdE3GEZ9lA/hfYPGLCDy3gsAeBIJEw00uf6+q2yls4
etBmPASlhmbBZdyYHAz87/GDEDjSduGESSUj1kThb2/TULBOz8FTsJdnBoIy9Xfzf2iQUoPVe/zH
XoazkcSEWHnQNAbDNP6j1eMEpwQInUqsVRREDTE1UVYjcvGwYBGjdwzSgZfVxUkJ+3qJFL35Lk3y
CO8qMbCrufAApcZeV1f+L65L6RIlIUau5C1rjHYDTR3UCM63bcmRVMdznatEZG/ju8mSHDZbtCuu
l/r7LynzpCzsILxnG2FxVohBm3k2MGeL57vtcBPE3iTd/E1EODFXrPlOCJor/HXKmuMQ/9hRxkTB
m4IzoXIk+sfKSim4A+9Hkg5qXt7/+bfrvA8cXmS9iVWhQGP3A6moSnrM1dmZDhfFAg+wuYtejIeL
37cImCDe4Ie7GjAhwmJoosaADNRiyhtG0Ne7a5vL9y/R13dRIQ0Sd+duq4lL0vTsan7H07f5OGdX
yH/lJeMnO9KzmUJlSdEpQp8KDS5UPdp3twxy6FRCYAs7MqDpL8bVU0saOiZayYbQ2YJZxR6QFVu1
0vRwAlg2XpuBPuIdAwzXfILIDhoQtv0Ae7ojY993xqfGpe5K45ZocYGGQslAt4jOly3lUv+oIfQN
HvxS1I2jmwOvmNm+bK1gSRiezeY1qGSKAKnNecXcwAFBU+KnNGgHoAMhKpZjbg3ly+kyA0i3lexP
KMlRhhDwQaeyZ0qjZH4VxjQ7sNJParJtM8mW5Nfso+TLu2GhCTfsJeDesAO/MeLSqA9P6MmpvtTJ
x3A5XxI1PHgjwH486/wcugVQ7KqHhEcNj5CpbY6cXS3xJjudauSrV81PtmtsPoGMrPE0vGQCOK52
SQcsseXPttbc11ypWJpos2zHIo20YnClluGdLPNwu9MFxuqtD5HBOXUKKTTo19BxZKeA4txhtIR+
rfJ2UpYd59apwcOus/rYeBzBfIkBi9ruRFB/6ei/OQoDURFhWolp2GYfFj07NW2P0dMkSq/lGEbw
tXj2hb3sfF7nA/Ty0hR7Pur+sI4lV7xCPuzOtuuvVzM4x74iDk5iCIVbWb3LZbwwV7+7vkNtUovf
zuA8HJCEyah1ZGxpjkupSTcWptTIkyOiVJqlqtFWRtHL7jozzuPOhHvBnLxLrhq/ixIdWHVv83rF
KsL5Dov19Zzy5XN87x5x0gOYL6Rj9+WDipW2Svk2tGFO3vY7JUH561ezFQNmXyYmPCAgTzYmaOHR
ZCcRvG7JT8oII58EPla764Fv6uid1fC30lvWaNZbj3QXAT7CSW1KWwylIyRNnBWpUkoLucDtre7V
PvN2WaTn0y+5dp1piQPrUVFx0mwlhj9E3lXpLuyvYpp1wF697+9G+TavBq8xVcFkKiggupzqnd40
IvdN2hs0izb5OMvgTuIgd6ZL0qhD7elA+aEWiocll9Cf+x+8/LKcyC86muRFktxfk8pF7rIviucS
T7W+7qFaxkyMNhB97wbVr0QBX6kpb6ubyN6xcv7zYza1SQlzZnDKhf07s4iU5snOGj/9ZIOXteu9
Tdf1ocXGC2azviSo55nB05bZlmhBcWmJx9mvCMukOe/DzW/mGnmj+olzaSldYddpbNimUdRksCPq
4YcdBCIhPJZF+44kBaeyyDzq8MI8/XN3LN/DLKe/dHRJ9hlYkvVa6gsQr/EEwdY/tgxFslnZqWNI
1eQxH0XllRxZRJltvmHvSQyz/kCL5MjvyUge1kwCO/dhOGoxNy3J48PPu4xkOHau1kD3m6bujfKV
q7Tnunv289PVGSGsRKaTbb9Z9C+DBkvJcssfqED6i4VO4XnlJPWZXDdQ330whgOzzkilcCuJ7FM0
bK2bfsOV6gS7Lc2GdkWSL0T6sJT4V7fYkdBWqq+8aZPByiYN2rklxPAzsIFjAyf92UfhIa68Toce
9FJkXq2VYzjIgSNMATo4nwhC1FRP6AKkX9/WuqHqfjVgXX+pJ7SYOO7AzGtbBuqEvVCiNEPuqV/h
xRmSm3TJJ/gpzb/sRJL93TciwpAt1XzVbZCa+itNYnEKj/rHf/t+GfK9LNUp7F4ZUwKQaK1skH+/
kUKUgsZuIPUDr7ofYr8vyXw9QvzaR+mB7aUZijf+8J5WSJwil80jZkILGali/8h7+IraAom3e41I
fY9XskVjA1FtcLUENApJc4tCWTzg1vBOSFPePXmd2CrOAniB1SXY94ksupKgqZIzfQQJTkl0Jq2B
QVW2mqmT950wZnaO3C+578GnbHQm3ugYaDc1AIu8A4u60pCabHhpjei+XcNMo8dIEooUqry9+yl4
5wYYsY0QEIMOKZ+ctOpxy76S7x2SjdH50IuHAhuCP/MzRVqOUbLQInKGspEQGj3DoYbcAj1djXBh
0ntpW3K8mNIHx7YDWc0NtHNPaC91MRNYXPPgTzGZub9an+qew9VE1OlAVQs6wPhYGC9k1QvdSiEL
JCSyrqJdhMVwX1Q+3jL42qNuITTcSgQ0XEfyKVCGcWcITQoxfdoxwtxZ2tlWZZFnN+E57pi/yd6F
BxS45P+QJJWHG27eSRqh9AhuE2pfDrh3kqFmNQ2E1bn1LONhh/G4HWGviMqPQ/ADlv0kzheiVU2L
rUremE6UdGwm78D46fJyRYoBUhwQ6TrziIikFeGAbTWh0wq6kMT3uw+hMoFP7dabudKHbr+UDjjT
UMIPFueZSxo5cM5hOOXer19EReVUWSsa83O9CsRsm8KnOzc64j9EFKFS8uET902eHxFsZQR7xsFw
hf4UDZU5hvcs61z4/ZIUsb1F/g/J9c5kZt/1slxrx2XVOOeiLAj4Vqu8aLRP+pyLU9NS5teTnmro
dWEjFqJLJkSDXKrO+3k7Vsb0ybbKxTN2OTPssO2thVXVb6AKiLM3In580hNMn3K3ZPG+lMcpua/8
JE1MmEU1+sgtZWGxCCpPSz2NixUx2PRLfDpEomxaRvuOOiFo6It825mU7TypiOB73MOHPRRlarQd
c8eE8YyisNJYcr0sVTIoWZ/39IVAapeDu3aBspwokKBhpqHS4vzXS/x59KnHWFjd9wmcfU/zhsSz
+BfmKvypzQJd3BoDjrY2ElPK+4MmpCP9tiwgZrBU0M4dWmUm0+29fd9vI/Y11D2q5g9WSp78wKKP
VoDCaFKjU7q/UePURCxkrirhvTcRla93J26MMrPvtb0ZV7zIlfPWo1GNwwQS+5JFKbWU8bIz7vnK
TYoX3p/WraK2BruLtC7G8vr55KdJkX5UMKZRe1x3m3t9IZMLCJIre2YhU7sPZoGO7RcrZVOK5moF
ineil9GAlZdnpITKszrSMTSEH45z91CwKTgK0Ztm7lT/l+MMpuyPJR6F/6NDHBroDWd8nZ6E/RXm
dtU2YzbvXc147s0SWOttfGZt8/lBeidXtoQpZVQsurHCtZAv/dGb49MHTpWlcKY4ouiv1dEpdL2j
GRFm6WZ1H/ZTbYXGzniDdkhGjdHX9jwHF6D8DQ6z9AqY9dCROm5gDwurBGk/QcXSPgttluR4Bnjr
oemJi1Kfnr/famWRICfHAmLkqVhmTjrdEBYA1jDsJfFzcdv/gJTfXGO3eEUkJgsAPyLliBUi4s7l
kS/qHCMzkJFsXI73/rCFG92Nhcrtptkhp6OpBtnN10BZtyyIToIeSCgo4abok5ZGJ/7bat2LfVfK
cQzQP69VR+i6GU6Q6W7XgKfzMEtxZiHAUld5DACJvkPLZDof4MpNGThuhtYv3jkDMHOh2Sck/Hxf
dtkJeoFOtb4FcfKtLsDmOMjt87BT7T+mFrbJ8VHvjc3GnIu9tUjnMIDoD21uPR3Ifl12CJZ3aA3p
Xeh8xPT4MieWZAyldsBwFYJR6K+4IFv4N8lieUbwENv74o2wIUKcNqgzvuodtXTI8XyBj9OABw7x
CoaCu80VyDZS+z5eEMTA6Lzt0754uBzSfZrua8vm83n4V34Sab4KGdNRcuGTumEN5Mat1SGo9WTy
U3dNhKVvZt1BcHgRJ4zd0aSH4Gi/y4wA8s9xlSZ/WpV2Q51kJiYWsPKXJNQ+rTYPUa5Dv/fjNDRd
Uw8XVE90SelGATM2OS5qplNjWKx3QOo5HkpWnZCC95/jVlbNQ67IpKfrxEVnDvlHxjuQf+5mv37F
BaJf1wIPFfIeQ+9cVLNlgrTpAbf4B6UTv16pDI0EGK8MFbNyuShhKwClH9l49fdHzUvCL5bwVeRx
MvgxNzUrBlvPf0luEZeCkZCiRRSvYN5RWiEdd9o8CAYxNa/CYobm4qGyVtfYFUAVl9tBX6L9qbhQ
KAUsO6nqDRutYHP8Ht+CLq395z+PGiwpx5SH9kp9BQP4D2jB5aAwIpZPMFxvoskc494UqWdiBaGC
qeTGbvsjFCBw6ZVRe8CzqsIWB72emfCGi9W/sl1F2L9CXWKTuQQgmJHIrQfBSVM16VuTq0X+RijV
IP+14D+lAbB4KEfoeOkWKyWIUTTtLWryTV7sxxzytt3PjdYkcXJhof8TxmaV6W8A3tKE9bVmUQEZ
XaWrZdNsrQCTmndJCDxCa2eeQXgA7FREt4oguksOcKXvvLW8PglQM7PaLwPvJmZHJE0py4FQkCmm
uHMMr3Anw/H9RRzWXktmoddNDIPt2CxRAYxN0vfydOkjQo5ZVVtCTta6U/dlYdS1/y92sxAgOmOT
i3OTSmAmJs/iRZrVuqT4abmiqz3qxK0thW/aXR+nbdLOf7omgXjMGG6Gah648QGY1v68nzs3axeB
DNba711Jptr/4q/lwFlik+9NOjQpOLzi1l7FYmiRxyh7g9apYJda0PZsXJpZyZal5pBBxXEt5r4F
W+emuHrMK9YsyjLZSrXsW8+9uoSW/Dcxetr7yy+cy0+6rt2oPaO1sAxDDkYkctnjf4CsZgTGWPT0
ycc9Ct3Ra3HqKIbm5Prlhet1W55rbe3ckq1HSQhNsCKGBMIzZ+mKk8hqgCH0O8N6jkRkoRAv6SER
Bdkls6FDraloM+uRf6JDXi7Ijs7iq2pxXm5IbEyFd3P/ptJ7YnjRN+k8t17XAPyuK/uDZXfZAh4v
nPg9kzh8QrmbJ4Sn9QhfBP4rNe1VPX/n6uZzl/LzUHUxqU2u7yQ1YSJJX2hVeVjHPlFDX31L5RMy
EEoutbqZl3UBFtnc1GuHr2i++eVhh4CB9D3g5L7OakGyMqMXRFe5r+kR0aJuAhKwFkeQXJLg2yau
xNKCM/f+/YO/zamEt8SGlWZ+KreHib6HKf3RSv/PE/ARH+H9TOK6NPiDs1bD4cPfgmI3DBOGCAtS
Vcf1DHkDf6DU/ySqvn70TfVd96mXpUXEpymRAqSqoOF60mKNXvmEyvKp9aE0sw2nyEkbx6VwtXII
/1+VZJ5okVNfgFX2Jxy2sS3i0+b88NzfbSEhGI2NuCQ2QxH9sWWfkDmGA5B2QVTJBM/xDtUh+GcJ
xuxITvjh+GLXnopvXp3p5bkejngS/JDeA9Skys98Sy+eEdb8xK8ho/QSyasWncF9l3qBLt9F/DTt
GTgOGOspSZKItk84FoQE0M0Stowe7tOGdDXBO1fNjnz/OzddgPEJ5Czo8mte2Ymz64q/vK5LLq8G
YNJxTFK8RNbELSllENo0IkwgVE5uvKat4oZJPItuo6w9mIba9CgKnGAv2bXAlny0YXA0+etxhOW2
UQgVS0FRXkQGXvuYCUOa2kVMMb67uAvfX9rTkLFNLpgXPqXo63/b6AKQoPsbQg1bySoSr1Bz/ldW
VZdNM2QoZfSXYryTj6klRyUtI5Jch6Xujevjvh8m2K0QbKeShW0vi04NzDw0hEtIBceH2fVyd3TY
Dij2S7Sci6cr3uFRfuq2BbLLPbcV/yQZfp5Q058qndc7VzFmxx/lXuL6FyjWLnwOSums7gO7T9lF
xYwDOmUs1p2+AYc0daic+R2nWMinIBQyFqK8/elsadz09VTDBy1Qy+tt3i5cJGeImq2JN0sFaNh9
lttNhIi0o9CljCutkv1xM/XLsXzkGokjHIw4uI9QgeUViBronQgwIG0u0gUOIuhMVxDgkAJriz1x
mykrQvcE2NZkIpwb109Jnq672bmRSyX78AJDGqv/wMT13Jld4FjEWrwsZhDPNR71lSZo5qLUbDEP
OmYh0ohtr0EzCJZfjiI+24masNrH6ZDRDxEfhLZ2jeWDCwBZf1VNF19baPdyEuI2VPsgVeFxyAlK
dbMN1ScvRNghiUEl6gxSSZ0zw1psJWmG8bs/SPdLRzDrMMyYNBmCpfsRwCv/i3KnqvkIlQuXJWkL
OAe98JUyHjRSY0NmQS2cbQjTe+RstOb0Lx6mEatv2wfCXrc3XnZyZUsREmkTWlcdaDKgcrlZtD6Q
NIUjZ2YeKrwZGkYFx8GTfjLQ9lmy+OgRqFrWoHRNRWDqzWkEbIcUJ/QYNld1h5UsFNzSa+KZQe8L
p/2+FRWgSg5ww1S+pbOnTmQdFPlEdYI31oOU73K9Afb5uw95vQMS/S6+BkVqWROKfYOP6iI3SOik
vPr13rwNOdx+ODh5XqUYZEIeXLXd5FE3EcnJrt86uITeL545jRTaVSGPhP/qip2wddzFlfViEpVj
0ToHEPT14zsmhcQFcklHH3ET9biQh/SQOkeXocCvdk7gEi4Ani/a6RB47f4ezrjtkSTZbXFPmoRF
5edQ+I9ziul1eiZjy29nVyS3ESmuCSMDqEWXb0jn6eyK1zBBL+U/8di+bAV9E6dNJh4PK2dxpPDB
4pW0zRSDaivXXswGtfoXkJVzxulsELPYFjLLHRWW0MyN40QufdK3hoEsKJkmnNX+u6QNPLe3yyd6
YUhSri0lfEqvl+wPwqDcaDt4JOOo45TfkLLq+yW5xFVnf8NBw5D9MCZTOJ8kLCxotno1lkwo3fT0
yoyMaqqk2DIBVcCm5xpSxIEkdaEe6Aoq89OUO0ZyGP7no8IgVHHBlBl6sLsJU5vL7RViX6i72GDE
M6F3QhecA3rWs7v1aJ8WXgSIz7Ryh7cMKdt7jZVX61OejMj7DUqVsmRU2oG3QJXZaTpMToVGzvkn
PPYqs5BwbXm3d6nsj+83/OWMXcr1MF6JBA45Vyx5zEv76G9SCsPPf/qN2sw0Hz0cmO+dqq84eA5y
wJu3bib1SQpA9dEj9fx2aStnvqDrGkjP357hlWQUeYBpwi5H5aVVp7gur9lIMU7/eKGjYnkNPnos
l7SaLBkzOsLLOq8TyzFR5BKQasNz+1F8cW7Yf0wLty/fg0jnMBsgCA5fni4v7LooQTxJYGk60i+N
cpyR6+4qAeZmr17XIk419r8uaQmqKT8NERQkP7ErBGSujqwN3eVVczYubo41S+qO7M9gFLn18O3Z
NpliAGn+ZCxNItl2I7xDS1kvgAbrfSrKpf0odqrD+PQA6Y1VVXIl6uSWAfQKJziRUBCO1/kU+Ca3
yRRNxOshwy7y3lNcZLDdY+wyOnJz9TI7JUVQxLGAB+e1CE2zyazuiYL3XaXf7UlprRKflbpuHJ6z
RXo03ecSPxOZG5HUet5owCEQXXKRqXePicVLOgF8hUnURmsJPN24gUve2ZQi8ijOuk+qjSQGfF81
dvyh1/kTKWEzHquB2C+4fceSt9gpxQG1dEkd/DjjtKkDqERhVwuThLKvwFw+npk6JUb4ss2rbAdt
BADwenqgEYmAkWs0q4N7mt/ECIDW3raNFVGp3LzXPM9F41UuhIiNBg3AeKz5h66VlTVCLf5PtFn/
Jccdfx9WJyyWEU4sorwaITG68Ym1JNQRgRLE59w0cTk89Hc2gCNM4tgw/VpscbJ4MKElN2lSudud
26UeljVtNRsYM/wV+BW7dQlnnxBb370NIh04CDG8Ip8/Oqc6Krulqaz63AZRBlGuSreuab5Egu1W
z+MHPKKtMrHpSgCmJ+r8kCgfyB4rxq9nrabym7T88f2YjylD/mnpCI+GtCIWuqU5qPTszDo7pg5q
/X1MjZTGpWbOkQU+c4lgt5oBWkWILt6iFIdW6PTidkwNMveg1k5aGZHVBi9ymgix/FzwlcYvEoze
7ixRNDEk4dSDhF/MlAUDJvC0O9SFnwgHxewOMb/rPaMRMkIW+rd51kTRz3zGW3PCgpuhMOhRohhE
6WoLN6ypnFFWL3Zwf269+76BKsGrHMou6xA+4ELq4k7vPboU5/dovq4q2hTgdERBw4mTnNcxo7Ts
ze9m/xqAdpKNKMQ3sLp6mkaToD5IYzmxl1ikgBhcuinnwl3X5VLl2gUChZlaQiVHX1g9lyxmDWuv
s4x44/zYBOddCa3mpWf6I3su5AJQAm93v73wIPO+lrhkudCDIi6aY1wZvXHgzoxwWuJreT9FNVWU
q5lPnJ6OepAjpRXnCL3Y1gv1jh2bssImuixK8TIUMAk3o/ZnXj3Rkue3cIGKhQY2eiKHWfBJem5H
h9o2eoCNTTRcoTHyJ4gXKeWPSqQLidLyljtrwriiLH3hUC5c+jozIina9W8okyeiO2lkOjY/HHcW
B2L8TJEzb7dowbTqVRUHp+oCrPu+AZ/xJuT91Pgr2wwpR4FHmHX+CqmB5DooOadaH0u45k9u7/FK
wi6uVtSf/vuX/4uoMV5RILcOc/St9K3BLJu+56WTO1/FkhwhEvoPs7fU6s4htxvTRLbXqIhKrJUJ
19n61E88+bVrTei5Z/q3mUZSLGrwAg7MLzli1OR/8igaRa36rkOZ4wWiZxZCiQSZhUpmd41GoVgy
z0ejL6aU0JCufiur31f5rsoLIY3TaQDcVsuI60gxu8PlNI22h4OGYgW3ltrSB6UCzciFvU0TBEuQ
QCzq5MnbpftnIYN6Tc8W88ojj51GhCH3UWpczsYS/44h0GRTLySG3jUDALADT6GEqxcxw/xSegzX
iZrdiHxUH97kOreaLuiBA+HL1gjs4CTSd+Jb1e+Ml0BS19stDO7dfBdwDj9IISFYv22G6TKAr5ND
OPlnWofuYwLyPdCaFi1gVpZX9+jNYfo/9fMTpJDnzE+utfUBIk23txKIDay3iwbYrZsCX++c5gLl
fYXcE/mKwOj0YfWh1p/bma57jYcaiG7m8gaKibFdF8/21Wf6aLtBK8C5lf8sgrvd87VkXZncD2C+
GAwIlp2sLeZycrYD8EHi+VPDueJBLWqVgXHu4KzwVQwpPmSTucB+99dSMG2BBGMc+WrCfoBMosWr
p68uF7w8CXr++37Zo+ujAjxJVGU1iOA3COj2mnJo7Osy5UsDIDnri6jqaHPIVkSlWsLhnyj7WC/7
yPZbW1NTEwyrEGJpQqo+CCQKqbiI8NYl+uWo1KUD6KI6NTulKoOG8+ljplmhj+D2YPEMWtSIvB87
olHAoB7xgEAszEXL/DKxXJgWndOjbSxL2jSBxLonh30NB9jKhCTa14bX/v2l5QpDVGwWkzQpanIp
KLvFn9Qs6ChyjrME6fOmqZ8/JAdKb7L6CxRvqPfb+OroN67l3kLo7PvfXGglsOw8m2w9NQ7JZOWe
JS+QSIRI8+rt6ang1bBWnWcZXyrLj+PfXTLeu4elwLVpguDUVbyxxoJ236lANoj8JzOF+twJXBPl
nAHVQDZBFlQHgpfiitm+EqWop23R50IbtWZn+2irYOfgH9veboo94wNjGH87j/8NunI4G4uuoOzG
xuCQf2pvEPJ+ReasKVfg1L/OuR+0kItEgNDoexEfJ4nM+ucf2/lTj70ppQdv8XCBUB1lQ7mmxzPi
GX6niUeq2OVGKuJSBjJ+R3lrirYvs3TZItOl7HXMB0XqQm0cNx0dJQ9NIi8tvYhad9Tlj0EO7o/B
+BeCOzpliy7aUDtwJcskDWhr30K6v3c2NYyRsoGMyFzTt9eqkSmXhgFXt36rd4Nx4LvoQ9cC2A4A
NcFjg8psQqhYfVNmz5U2qzlJyBWRsY5irHU+vFgoUtIgAayoBB88Iga3CPbXz3oJGq3tDVAZ31DA
PlWmqev2cvFKoTqy7/IzTYj3e1sVYdf6OWeMShbE9VaHIet37M4KqMWZsbcR0db90mty8N4N0Smr
KaZA42TU/t2zHJDoGHwmOtb2j0C4+rjmvFpd0sUNS1QmGBFJwxWyiqLUoIYm6mdQgdqDMkxGd2SP
aa7+6z3PfS2y0kDrvYMKnRY8b3kcjEWOT6hXrM1gn/vxcdC9Hpy0ckN/rfc71/ZfY/4fHOfMo3hq
a9gMHgjpgK3A+Kl/T1UIBeDZkKxynEAAk8qPT3cMrRtP8FNfzuoWD8Z+3qs4QU6wlUwQvVTrNk2w
cBlTy/sOj65Adpjivf4SACOd3rymqDKD9/IWrLLsq1N+bSbinSicU7ib8kJX4xXPsyyLuTEQ3PCu
U+h+i2QxeeaH3XKjg2vmwZyf0hCXuhM125wlA97hqvc2i3OHtClnNqPBKryNvI9rNgnlDBYaa7sS
6D0WbePqs5iHRb2uzBsEI/SJHYkGs0x8u3At+rPgWSKTJi75TrFfKv1Y0g4rD4VlxHq/Pbb0gD2U
/MVmi+hbrOOW/jfGwulDyaf6TUPt0SAwNOR63AW8Jvpn5ANY0hHgITZEa5pdb2uR+Mh98DaT/CmD
7G/FYbopvh7TFqCEhTIIczV+/Sj514EwDKzkLI8EXnQAM5zADW8a6hwTN+qrFO/9xEOd1utRD+yw
xOGNRIoa/JMRrEFtakfibIdyKUpYh6gRZ/5YU5VzQjdCGYcw/D4IUdGCkPGIYoCDd00J5Z/0lpy+
lbwWQd/DxRtP0EZ6Rnw5xgmeHggXXwL9btbys/w5sp532AgUnAS1vJHYET8AFIrnSuHoRgFHp8Ai
sXhCj7IQhB11Z/8/lbAcx8bDIAIDcuisRvnys6nPIb5OEpghdX4eV2BMwmMT7mbv0WRjskxJyBSB
BYr7Rm586wucu9m7v06jBCwcaT9R4lzKTMBXv0luAxsduKb/HwOqWQvghTLyN8+IZF5bM0B0Y1KX
+qHOa9zbiRCNz5wtD62EU8e8WA2eq5sDTVvhfN3N4ts/fyerpPbH6A6zGr4CMQtOK/Luvnihei75
E6xTNbDB3+ZH//9j1YhzlmYaUL+HDQbGm4AKGqK++wdQ9ANI5aIAkvG9vcfXzrlsVsis2tPhnpNT
eTlbiF6E3cmAJhcS79cZzrArtsG3qwg+ZzrqQEh2XO5GivvJQ6q7PAxy2LPchW7OMDEtmuNc5gCw
vDWqrPbA8T5Jl29OKy7WmgF2oCHr8+43Qt5v4IESW8u0Gsy/iC0zbIebeaCUAFBY7wizWIRqbOXJ
9X/bgNkwn0LxvqJ7fc/9iSS+YDnmC5DO9UKcUHHmooa65V9VJNaNacj7XqbPGbRA+DZjiSSTVJ4Q
sKZj06UD0xOYJX3nqvUmzl9Wk3RDwRrcuqIDZ7vKGbu5VD5ZECz05GQ/+Jx3AvijvjN4PhpSaxKv
3ersSWfwe2B/BiDua3D8ExlkPQD/8MaOhikBjj2hnI4fpcTKs2rWf5JcyvmvXmgU3BW65i1ZTvtF
mXyhSIo1FrWaNZrHDaiCdY/aMPJuKhH9N+kQD/vEURk1GVnHEmIiqMPz14NSX6n8AiJ+BRTT+I/J
XrvLRmrGmejBiP9KA7UlXmcz+f91UbpPNLRFAOG0JYfsFPoZ8x6KThJ88NdxAKE86kpOJlee6SOL
n1HFazBu9DURH3jplFzZ5AA7EDQGoO/oSWc7+M496i9lXlEsEvgyzUMJEa5wQT6AYixuMRU9FIOT
OKf80V/Ar+Q1SwSenY19AGIkUyL7yY/lnVab8ZMgElQnhwRuP4C7WpMIUYvbo07XIrMA6reo3H18
YMkqy+0XKC53ivA4Y8HVxyTjyuQYQUPaSYk4Gd/PYqgYS8Wbi6/KcoeS7HsNhpCh2jS9848I2A4T
ih+yjaHgSakmUDW9D7nQjwlTVLzPJ+yyo3nI3E7A+8QmkpZCuF+cWHAaiHswrPf12dIQjEqti0Hf
/3UOXk1EHuLR4/XOTnKXxNKUzZ//GrF5v9R9BqJfUnIvsoJlv3zy2xQsd+rV6hfZbrqIG2s1gRCU
+vEKKpq6n8/S9PUvRxJwHkHMSkeUdHd6cGL1kcLDTo6ZXffJWCfK2eDO4PJNZ6BqMgrncRLurpoY
yN0UIVep1NSyK3qYJVXi+vvEWxOk25aCoewu0hNUtUIUnqIqSYaztF8TRKpYXRGoiyOjBSnQvv6v
wcuEvdTFSiJ+arppYSzXvAw8FlPwBYCeRjeY62apXb2YtZjqb729ledKWaIdk9fDgN9fxOl+bAhF
yjSFAag+0qyNVumIvQADML1VOpVEpZh5W2WEmEEhRJCKWeoDbDFqz1uwR8dvsoA73Exs/WaN5HwK
y3DZSlRCmJqsLFFdjJEl0/pumqMQAc+hO1tDywm5vQupVvgv1BjAXnoggxy2wKfIj4qMyJGc/WG7
BZ4jKZKPoc4PBz4qf1iOiKs4/53O7Nc1WxK604bdhuDG2nmMaA+AmNTwPkT3IWFjPZw+2U6S328l
TZ2xkPPgn71514hsZ6XNota7RrzCOhOi7vwORAbkGtzJCbuvVLMeg2HWZN4vTvI0iPwe3Yi+juir
9D6Qju86TMuK9/yuplEmekgv7GnguNJE2oUV3+/hwNQWLV3GPoRXFLGdzY2DIdHxH5q4RgiNwY+v
RkBhYGevLwTAb8u5JDh19+Hb4r1HiR2mZ7Z8opLMjW/XE3/qt1YdKXzq3RW5GWcnwzVAFHEb3aXS
Bab2jCZzpEMQTmB5+sB3n/yg+CzevfUNn4aaBKHmILAe2Qzn+Xk6deCaOf6LSTihVkr1ssPn+u5V
k7pyNPD5o8fs62tzLiUWeCJTHShLKA7JFX8mwwP4bP5CDniRDFcg9jshPRQipyjo3uf4Vc78Zw4p
BqoaHeDYLXR7pnaGiX/v1BBcSTid71Znn2Fz6N7sD0rYZJzyG8wddmuZAdmyUO1/8H4upPha0oTH
zv2UBl30UVLeeKLfj1o0k8eHYJjemNEuumOO/kN1QeMOz9/Tcg/PxS1C3fpbH9Fsj+0jWWEoYWLy
dzi1p9lTv6CBDijQ46/mqsjCgI+Sq15si422T12DGXhT0Rv87cvsC3t0vn1MTOyYH4SHFb/u3jA/
wFbtXC1bJy6E4hbD+UfDEYsu897X/YlJURuqKlyZJu5xR0Zgw1APsnINBf1798zj8yOh1fEpOxkV
hPFbYcG7/9wdgykO2omVewth3RwN/t/gwxmtQI1tO1UPj3v5XUn/R3ular6KWqXcW7pOuZcliCLH
sP/lsY0VwHqPyti3qsDdLUiat8jHKLaBYKPirlf0JNNvPGv7g7POMau/Uy4ZLtBSXHO4AHzX7TbM
/o9eU6Lc/BVSgneIZNUXyXtLwc2osEw2I0NZEGGQPro4Xc0mM1TF1/hIZYbZF6HSPTnkbPRREwEf
ZLy81ddNvu6jlPz+wD4CXz3ume1puJAzBtHJodtVo35TjygEEdvfulIYeeVjdzaEuNtDGFazDgAr
syOiRPtzKApWIv02K8NXzLKSIbOpdBqIK0eV7zEaj7d6zAKu9aGyf1rWMF6LjiFXlPwy79BmSk1J
Jf01h+KwQWYWgAe/XjrZRxfK7wAfkoqWkNVLtFfmFvEX1GPsFSl7Otssb9DzIrwmUTfKzMqSDu6w
Ra0N0AbA2mzuVMnprPE2TAk1y5azPIZhmwGbVEApKdAEWOau38JHNvXz93U5XlMSeifGDIx+XJC0
4IO38W6RzKtJKbc9yYXS04jX4DZ9qq2akqK9W/wGZzZsghkaJGDnZjghQW7TEpgnl5ZXk6pwbUq6
KrAtN5jP2Q6sHT5zBf9uUVtAj1EFOVz4mHMzv1019y+TFtIUdETYZD84eNYZw92kco0nYKoiZ+VA
BW+20JY3CLzZ18Tm/JKGyrNtGaMgDq8MtpL7+ghL2LZDwsmuoskTUCm1kE1Gr6tkPKVQgmjNo3ta
tvo/TVjXSj3GH7vVdeNj/v/k0tQ6uiGzj2FBYsnpVR8bSTRDkMjV1Y3wBGM4kCgZG/s97d792OMS
G0BP89BzWa22Hph8TFXFXFmpr78yFFC28+jgG1MpWZ+SHHGnqbzAoruD+z1lX4f7lbsDupvp4NbZ
117e9ZbuD+uY8TdkOaC9AWjiaNJEPyqYvdKl2HFDw9qmVJkzqxcvQ4Z2K8et4m56mnVfmZEbdjQ5
fRWKEPCrC6qZiGkz12oP1maqy7DRJ6IphcqCibad+/Ovw6B1KsCxfQaLaHCPbfRjKcJd6oGXO5s/
CdYHqi0XjDpfLRHhnliIlxfUoxAg3xcmHqJ6X1sDO4vlUwJ47x6bghyfBSLqHqMby18uL84SJe7R
MqYusyTomhdmhuBuPmf+owOutyOg3EaLhrfYbXhF0yeSgMkUl5fYZwfZXMGFwTacECrzm5A/FXy3
LPcqjznEyBfFUwYmveLfM5AJiXzc+79EH2wgRhd8uYtrrFWjAZt9Z37eRZk3x78nL7ekdNnI38ye
2MklioFaPV30wR4CqiWEyFxU0RNNvoeScbdcStFDMXKsvqyGeFfl6EKoLGlXmsjEUyhuf9YDFZ7E
FqTztT1NyJHdveYBq54cqcZ3iIlrHPvptnltu9WHBQLdg18d3+xLRuIGYpozCthxfYjUH+j4woLo
1XC4PoyIhzp3EvcPX7Ygij5nkXI/8s0Hnen5LEqhg2nQ6xGBx/uqixzwaIQlaBsUNEfAWqkoN8AS
i0zU9er3NRWH7UF7qtIDiUoJJ5enscWoSBJRjtb085Z7s6vaT1JfMLeRS7uc90fgGjpiHO7IxrMH
vlsX9JneTPgNIBqsxgInV+0u4rSxWtp6rb1Re+7uvo751ns3BhheJkqeJURQz5DnplgXwxG6ydx7
tO5DeXDohdX+FQcn5H4dMJtB8mseoSUUBT/qLM0gNF1e28JRtC4gk6SaEVPJtSQwQYWvM5C/j5S3
iutIyUj2Kdqbe9RG6/JFZ3G/D/TOldjz9yOjgEfFe09V0+oQYQTg+BlCXridA4JpQQBm1FghlCzj
GDNz5gZun+9ZmJ2OUKx5Ajr+bBf274mMy29N2LX5z5xa2Q3bNcthPXo9lAWyEL6ctBEzN0TFiSns
u67l1OYSfSMTpi2H7oy3oICDNaTEP9va4p3GZkdREHHVUt93LICIRyWCxcyqx944Lq8jIdRpAlm2
N6EiP8fa9LjTfzm0UHGdkTFEuYY3buH+pXbHKm9QZOjbBXylPXDNHy9gViqHvclYME2z8UehL0PM
Y2hoWnqqGw+sSymqjJWVCObfQ8YkDIANr+neny4OyprYyRJGIcl18suN5UHNqYy+wGfJGaV4C9Lk
Kedx3D8+KPhVQgCRxJ+X+xiTM/O7Qg5OY749ijevhjyqbnti/U0vK4hJjNmqfJxlcPSu4ZHzwkQV
s0Lc+X6MHlIS6dAXjY41ax0+PnEF4V4HtHhh9EnSMFiHBvXsXHXKIBCzHlz0chcIEz1LGUuyIpDb
LQIO6w21u3z/HhaWSW3mcuy7OxUw9X8VseUBb+NuuBvzNbkZVdbiThL3/kICAmhbAPmpfKShH0YQ
ityKozuvS3dDxPG7jV5KMK6fEzcnorzttJg0A6uRBu3imT413flxUEDLH0+X1RvDB70lDCDk1zai
ve3b/JcLM/h9Ya3PfNRkPbVeuuWlx+VNHT4tKncgktJRE7EAiAtwMEXIx4Li6I/MYeHwB9ocYV8e
+r3TlKTrEvJQ5An6mDlYrGOtNgfh8i04/DNNWUMnmTvcukPlnymzPWWWvvvI3Ck2Ot67PO8qdjtj
/0vrOTUbRE6CzgftI4FBlsMYJAk/+VjCO2Wu4a7+FCYe3tXAF0GTOgqwDrbyae9UcY3zY4yh+fUH
CwM9h6KmiktmkV0wFuQ/Y7z1ItVnAy985IKOpjw9+jbV6QyzAVZJ2jx3uhRROY7wr5+W3iaqIa3M
6BIeQ/i/zcG72RDyZeoHLuAIVkasRB+M2QiPjbLFOSZArqG/t/gNtOpBcYZHE4uwLuq0rt4PPcIO
CocAS71PycfeeqZkC4bh3pOFa0C6HOarXp6CzyyhU6o3Hdpk4uv+fUjfvVOnEWqPHK3NcS5gIA2K
LOtYWi7pbHp2T14pZ8Gdn3uZj/AuznVS1y39Nz5cCN0EouSkE1UZ5ie22YZZ8N6f1c0U+rq13kqe
+Zn453F6/uTW7jAk8rl3t9FcMuDgoA45TI0sQLqzepXYHx8y3klY/IstLU4z32uwMgIf9pFfAvx7
rUtPGFWN1WWrXK/1twLQWKUArDP6pYEhK0K03ib9BztxYMeDfSx5QBzYRKS85wgCFwLNKQoAePSD
9K78YGp6pwGCNkKKP09MXDxi+OMeDAcFYpV7d/Y7uBr9eRDOX9VS37SKc22+1EtaEkSPs7DPB2VR
WjCVGLddr78M9hBfLAya5BwaCXHhfQgfbI3EDFsIvJHDQLvgaLrPp4fd2sCwDsMmE7Ib6sFKe4bg
f0jTgClsWRR2dUfG/2LYqV5yAxeuxwXrWQKsn52SxyqzZ3d9KC0RQrS2vuoCuGtaQ3pV3szBlt0P
jnSQCiQ4l1Lbzan6L7UTkBgjLdrtIo49i9XA484VT8j4qTsjbiv0ui2+v0D86pNXgPWX7emad9kx
tKLJOEL0MboAFeAc9qOYOVoG88e/qcpzcYCCbW89pa1alU8MdSrsuA0iV06pk8tWn7srJGkvyTKC
NdYXfLGxbsmHyVuw+V0yEu737tCMYOBlz6lTJcyDCEbuISBzsJnceWBsS0fJ0ulpW2fdGXYiI3p/
yfY+0zb8XouBZQOaz8muW7lBBJqTmvtBhzd1EY3xv28gBnd/+CoiiYFDjUJulUVMTpXutVI/sHVR
TWlBVxtnGt6GPvPUX67ZcQEI9uXuh+lWh5LPCrYVoMBQA//qncQtDPFiq8//9M0tg9T0cL9PGdCq
N1SBTNzJNvNn+oM/YPcC3Po7I4ulhK8I0QhmbxgT3d+2zHDFZRCfRQF0Y1u54D1tfOv7KcZbTsmr
NU4jRDULjjnNs7/GJKCWez7jL1IwLrsmXzs5X4PYjd5G1sFCIIRdo+8nRxT0aiFHBrlJTzyTkfoV
eb3J6keNDkdEnQGnsDGisxznOHxboPLSU6DlOmTqq48ytovw3Zmjh397gNfTUulOLIfs89OwcJHM
VbSWkxVaJP1jE/KO92q1vXpgW75cXpLAGVeP6nyL6EH+iThxd4qZQbTyJbibgswkKGjViPf0tIfM
l+018z0L6pVOZCk7639oORa20hfmntlZnaQA68QZ2Q3GiQC6LsqosQGWmDVKD0Gd8JTe+eVI/cNo
K2sd4XlC429058hXDR38YOF4duzp3onCFjaqq2/p2m7y7Ts4XOlZHcpw4Zht47bZJLKAwuGhsl7A
Ei2uMMYrVDTrztVG8XnE41gRWegTYf00o1FlK3pEZGZ5JPCUL3NbiJk3MkDuEKA1dG0D3VH+juXr
Vfvt2L/6Rek6v+hD9EYojVN1rf243In2BXQxBPR9Ajr/RyyFbB+EBiLnj4MZzdqfXb4gwqILFM0y
EGKjgfxXWPGJOgl/yxZ3jK2G8ywy/ch9z3n7Ua8B5W/nuKiTRQO/y6onHszmTH7/IW2z0DZmB852
CfvVW38jSOPtDgoDk7O/2DrwDtWZjVFNuyELoH6wxXKJm4U30F6IgVKrpsUZHBG4EP2RC2prmn0W
IBOKXH1jGhtUrB9vQ/hogcPT15oX3sEhiz0NTfiWCmEs0QLV9H88yvopF/TtFSPee1KnFcpJT00h
7tvS8/pxynBGfC06IXSKh+PxpENqY/FCgsKbwHgVKdd2K20tdkNlsS1qpliOl4NG+uBdB4ock5Kh
tsPF7POi6vmgpsq3OW1TCxynuNBqaNhrf9SIKDEDchhgTJsuk9x5OM/aHVHTk46KfVK8Z2GwB7ua
oMWoMGhBFd/2vG8QglsQFigDD6ADVQxuvY4AjQE/+XRiqcc1CNEHgyDIiZGYE1QwAT7SZDfn9IFV
JLF4woazt4ErmAjQBf9TQ5FbLeN5VE076ltFu1UyMdzhmnpLgLbNCacPVWNeJWZFudI3lQRnoQvV
OF/1t3IfYbQ2Wr62vsoWr8Ohn8CEmA5BF21/04qWlD1jsLWeHOiCQXZxrGHZYBuISjxYI09SckfB
2yNkWvSv8Np2CyoOT7jOuUMEtGHNJV4rkJZYhaNFUkcphcx43Al2FS0wN50TZnvXudzjOqnbQK9e
2o3LoyQu7n2BRijZQgTuHYRb9GZcOARWtuO+uGqpriTd0uGYUlL/U3AOGCGkvfAqRc/Pf+92L36+
vlYEU9vNH43LgldJ284SVStvYz9v4VU1UFbhXArYh/5t1MSTo6VF8/zcym+DMskqknRrTG4BN5KJ
5DYbf4amWfXDk+RVurKUlB09xQ7vOkiVxA3Y0FBFIucYXBIrYDResMw/DOkThFePZHXX7vaLfwFm
5zCs/UPDdIljPdOvqGu3F1lXPxsMGlgD9WdgDWB/+BqbE1EsuUmYgOzMkTgO8yZDOhd51D62/gi+
wl5WW/4tuD/rhF7GFoWTOnV9EDEySSVsKfkbekWaz2/fJUh70YPFofzN5Cx+0q2U06dBG6S+K75L
Z/LM/rypbQMSMa7h60Jo3m3B/49fkKr9Y+lYc9o4jUj4KfFBgjUCjk1miO2kxUX2lv6IYj458KsW
xbgf8lhMEcNceKwutPKGIGGIMDbB1oGRrb/gSF92fqB5xqRBAwY6wveq8X1012zWB00QsQ/TdbuF
ZEQ62ghtlVBNSQFTHio4YY+8n96ZXU//PArCLZqQ/h9zNH6qAyx+FPQR8SF/9E0gKXzxuaS6YXQx
s5roU0bDi/EGvmZ1KLGlkGMYRs61Ad27xPj9SCpGzocGkiQ7Vv+CTYUUhHEhZ+gwNW5xO2RVTHcx
g90gcKWayuimheHd15vjyEgnTpfi5ZPnSBvA/+7w+krQqPmlkbfsIyOeFLnFPbU1hwEdi83y6hzE
Ay3U0IXFmRtTn4GzUJo2NcHqSz0gfKN/iW2d++gSt3XfMcjkJ+OCISXfajiNgDbV/QTqGWYy6AHk
nfaIZWYh6b372HZ9IqQjJd+zcL/Ku1gPFLe2jt5LMnrrX3GCOGuow2UXFrnNzxFj478vtxsaJ9bE
XQwpDNtDjG+esjq6yZEczdIkl0odc4myvsk3ycncviUwnw8l10g5QG6Vsh93wvoOkaryEzaBYIJm
hVbBwfTnDTD9GF0BxLCnNZCJ7wY37wMcyHlEkk26C+7T3uKgUX0+3x0QSZqfsoR4+yOy5+MVo0FX
/Y0CY+ooBsrjeGbypbOI+PjJjBaXOcxAHjgEtEVCEQ4vbrzjIedHFd98WAjX+mUOYoMvkOZkdu82
3eCVU6HjtlqYHxCDE7RhVnBIBsMJP9isbfRSB/sjQbbcL4ayif05joBM0Q/E5EBCG480a7/yXjMG
ZGV3Fyo5yzCDmUM3RqZONG4UO3SHYh4QS4StLOKyzAgLxkiHRdya8EnBRWTQIOlmv/1as5/YNc2Q
vgNI+GNI5Pvoixa4NABEhMwW8rMQa1xRTBWkqpMOkGmKpHo0FABZsZ62UEp6KaRDy2WpTsv0dGaX
WNMHxLpvFQfUXTR3mCDzUdgp5h+GfIbwpkAYwvV16cAgyhC1baU64eexUmTWtGaiQU6bxA5eLSlM
0BM4YDiRFrU/sAj2ofC4s9UjWb1fOKQ3FnTqhcYS3VubO/ggaXYnEK+fPRAPbbq0QJO13NbvQKp5
qhcImr5d9H6ZogJsrZ72lfpRpDqcG0iLSDhSh2ETLwdnrjqYnKJ/XUN6J78f071XqXewoSGwD2PG
COB5j3elyuD8PSfeWCx8zrAb6N3uJaRziNGfgInx9cfR8EGqhYhC7oQOXILlwlbQfda9eY/nJGm2
33S4zJFnaCvisxk6E5b4Z9A9GGsMgpp6zVmTEM4CojbhoAaKWlS6ysW97u96HVL9rO7515bJinj1
RQ3DIimZHxp5bwenYbKng/cT1E4Ia7XFSMtlVlx5YbHx59rdcT6gjlObS0WW/iGBn4sPsXJyQ0lM
Yo3EOF9kNh9tXtKgRIo2PtWDW2ZNn3PUdi0EuJcbE7U6Yp6/B30d0M2fz13X0EjyNlb7EtK6P8fm
fI49rEojKgZ45cDdpqAso5Hf56zm5F4EEsTP0t46WMyVr//vwa1xjea3TEJdcP74nLvMDTfQyjfl
G6s0YGGnHMXbZg62XlZCl9Vux0dKIVjfQY5NWn3DYr6ADPNSqHZ9JSnB6LyPR7XbwcGifsqh2PWX
2XsKnzCwms8h9ul2Slzbq/LUNpcPfriYLAvCUMdYALFeuKmseJYI8P978JJe88T6o8qUdkarzQxA
1g7dRCSSd0cHVZzgr6mW/yeFVXJ9scfQIgbpmVwFc8Bx8PU/dKB1l0e23v831ZT5eVLX0U5dPlOP
NRbDVsGnamwenF+VKgu30rfBvwseH1CTuxcnS8NP8YO+E3+27AQAWOy+hlvn1CkvKw7SJ5bN9d7q
ka5TIIQv3DWkFLCM9DXJwmpjSqUBLLQyURyVkgiOFnci3s+YTezwlz4ZAAU9WK0BPy3LgWbXlCPL
CBUG7tKWzcD+G/nOILbGDFM3W3pWSyoYI7eJ1H+lVRND/b9YianfarvZB17pnzBnb1uxqqUMB7od
P/QJ7Hzo6hBM1WMWjYHMLH/ugYhEWiK/Ap3VJA3KoYShHBX3Y4SHVAEn8nJPFfyCnAHDA9e/CkFG
gGO3eKqRJwsfTEF1+TFZKZfU43y4vUorr1pPABV1FeEVlFtlKvbkAEdP67wVcqhsqEziJa6p7mdG
n6sKXJAxmJByyuEHaKG8MXl33cqntg/MBnEJhoNLxTX0XKFN+9Nuaj75w4bpdC0FqhgbUjT/dTMh
S+ExKlCS70jWOqfKFhVPjd6HSZE1ye7lxuZMzo5TgiObWlm3t8cvgUaUKYQN5+yzq+wqeIMFqXxM
cYclp2O2YkrtUhzeRHAp3hQAmkcCwLf325QY5vZfKiWfDijE1hGeBZ3nBIpFGY6GVTK7rpzvd/ob
wjpVDvOXtT1CZTxyrdw/HtZQHlaot5w5p6N05praMR459enG4mC/C6A19kr+Ke5+7n7Ri2RlJGU/
Z5Fr+M3GcpKT8nIKw2DuH9pJeiqaw1cpfEEcRHx/HApMZZVmNbN+yLeDt3dfUZvMjwXBfccEyqIs
MY19t39Q95Qhtdj55krKhRVrG7bEkpz84jW75j317mitpaiK+Wt6OYM4vMhUkGTgTZwHioZYhF+d
0pjSdiLZ2Y/fej0ZC7BbGKiM+z2w49KHAOAup/RaSU5UILi8sM4f+f6WfPdKieKSuG1tYvshoqNv
oObXBhrxR6+X3t0cR+OZWaDKRZn67cBz6apcG3XQLThq1n5WZ+tSPdzsgGaWYz/eb8txVq/Ixonn
8fzsouNdIpHWgjZD3b58TfALMKUXWgR+JwHWQfGTXQ00O+stxIczWQNpN1AY6ldUgMHrAItTWbi+
Yp7nT75tfpurasg2+lSUkGl/zA703gwFivF2mTbbYbfo80/WdLWM3aP0SKr0dj2QxaKSmhg5+9Li
O49kvl45aTEfYcOk16NECY7zG3VNliAkav79VekI+Er+Dd8ixzW4do9ZTXyKHJDhBvAK/OWQguu3
Jd+0YTJQPC2zvVpdz4oAtKMbnntU7Do6Ni1ZiaN0Sa00E5hB+3KIkXWEGz8Oimvw68nRI/l1n5TK
8YdRN4J/UqsSu7cfYdtTdFntn8NbSmZF9TBzaneDTytjcvNQ7ED16uGCDjkz1X7phnYPmf3X9VqZ
lVFLn12HJr3M4KpZ4/RyIuVx/JmPRKXh8HcHqXxa6iNWeQfguYOsSnuByX9dzDYIYbVS9lFucLdP
b9kunbh0wMMg4M7B9uHC9XeFLOjDiDTfRpURMn/FDJIPWPdEiBBXxUh5y1h0LFyKEvB1uObfWxRJ
7rTZZqPkWoqG3M0yBbCuM4S/Gq41Hv9kurMi4n2iOt81Ri4DAmdflYu/E+SHCGmUYltSu6YQ+V+g
3Z9ccFiMhkjL/Md2mrbfHPWIQ+2Qqv1ORMCXLCXttDKxCBKuc++Kd+I/3Jk3oXl9MqJCiudZPVyu
td9BMhAa/Ka0EdfiaRMIC9r7Z0x9bFPvqS8RL8kiSGlfJZNvnI+B5ubiauH1KzzYa1qNpQg02vt7
Ictath9qjpKLSOVUNb4ydSrgjMbRTH7mVwhjDbUqkGfXXW0ny0jgEzOinQH/s6HLyl2vPF0KCwtj
IlICftzoztPqPRkh8kjFw4infWGfCvD0JcFnT186JBq0R+02cTUFWoAZWArSP4jVPK68wY2FR3h2
h6Uhhe6o6HiNipEmnLzqr9iqF880AAJgVnF1Vdw6ryBCLceKRv+XlyUr+m9idI+O2l0cjuOppUA8
GWXDrIcSeRkSmQyKz5EuBFDUfEcNjlXKpOrC3WBRy05xxY2NFNI0x7GLfY3lW/GZNQ7DHLLaQOtz
jdlFcLkc/doHS+IC5n/3rQuK0n1Ukldl9Snn3FS99E3VK5cE+xv+uf1M4NTwf10BkE/8broJi9DF
j0JkTYL7NwohzybjJgOxjIoLMtn/lBcV3PRMGFI9LAqhSJsu+70KUGm5cmIfAfRSbEgtjw7EuLvI
nS4J9Dx0XXhoLZ2QeUEN8EPxSVt1VS5ekFk3mSAXwGAT2xOB542jn9NyvZGO9KqGhAa4l8e3D7zx
h5Z76UWIeV6orY2CLM9sBOS/bRQtX9MUawlnGcoAQuxLEfCzgfQyZQjR/ZGBDEQvOs5yrZZ3yKIb
XYlS+sZd60sx3dOG4dImJFxycM2bgJt3AV7gV5Wa/1+ChFLXlZrBhbGL11oTNgz7XlZ8M94laX9M
3HUWVP9TEbQuWTYMsXX0dpycDpoqmZNTXUXEoHSsYnCunFWSFN4mg6xr8x2ZLSyBM0xv97cgvAjj
xPzkB07bsU6Slx35Eb2Jf6EUysFzH2UZd95XRJGA1vzobLk52U4xq8rh2LddM59Hzwjid0dDuL0d
4Ckj0LU2KSINMl3qw7LgK9v0YbMJbWXWzmThNCIjwIkH2lQjr8UQ+6V4KOpUoXoZbUcJK+ECFigR
uqQk9jYr34Z3Phmae+xfcwNwS2oxs3iQV+FMecbZmXIwWKq7xXcBJP3saYbRWst6/gAy9AOgbzdx
E6oYDIX6DAR2hwQ67wFQeOOnBsb1csjRWXYD1IbyDDRvVyGaYraYUEwLfzc2tEBv5j77zFg5ct0L
r3cBD6hR+LBILryOzAfiHp2lTdqFynhJhK18pJ5e1a7JfupJr48/3s73FJZTxkFlHluzfFuc6Bui
v/rgQ1ZNyrAU2Dug7uAFVv4FE7fa0Dtp/Z+YFNsSIoc1DiHHPgIrENv3reYHQXk7CMYpmfaL5TB7
f6HsAUMbGzTdAyAidXxlEvauHaHfuM9YUuEUN88/K88rxb8sxZHIifXXaecWMmmGzqVQEIscr4+4
MLsLRjx1HcTcI9NLiPv4ThMpVLMd1ofpyxNcB5FG0MbfniHGV/EYonV/lDP0k4QrKcEWHLeV/DGW
Vxwr/SasR3CW5Bqbf5imVUr8h28GHLJSXVo8icCyN5JE6FmVhqS8Xn6rV+5YOOmCAH3k+y4NyjNQ
tLRwrRXOrM8xakVlouRDD+77jwMhQ3tpd4ywWITFJ4xPrKkMlniyfiBEygYx2aSRSQ0rIwV8Er1+
EG5EYE582IzqNlRr7agm+SiBQ68Yv0+tR63ncHVl4rLdnwfEPaZdstlMZtkYAF685V3EkzcX6+mb
1//pPqEn7h437H8QbXC00TRRbPcPmky3U5ezk9i6AK1ymwy9avXqu1jEoHJMxFB5iXcphV+6vuUt
MC6TUV1UGhfZFibtWhEx8yCc3SSc8up7F1i9Wg702YnZZgqWiBsa5gCjF6CmURpBIjeR93tI5I29
AIWQSwMptQJk7dcYfiFNmK0EnnQEZAk/6XPnnIIc8Daa3GCWgrQ04I5YTpj5Q+DcQdLxezki8wYI
iVJZK1Q1gB5NF1YQYGqWdfNVHYMJcyvXxSEk1iRkW7c7wdJWCRoQdalyOStf/Tag0oE/kbULv6pe
acqZaLFeOJm56k5xABWnqDuNmdGx42gg+/epx22mAq5bcZD984Vx735iknEPEyj5eKfvFQE0eZU9
snwKxDo70xW59BP7rQArfD9w3QXJnfu3UN45EdZPJrKG1ZsmzWEBwAgSKxlFYttZGS3vJHz+zVPZ
pJnusbZBMDXZdTbXue5Gh9rWwylGDdDPKn3GGtbHoQG48fGA2+qT8nwp0Aw/X14PtV4En/Q0gY8n
7qrLRmSt4/K5OW37Wp998ltwpSd4o/rJxxEJ9Kl679sRKqAVWzezobsb77HZmuwOYQfGteZco1Im
jh9J9ECoKVeNYOZb0J/+Wn12DnK6ODgwKBOU3k1naOWHMh61tKml/Kce0SW5xYpEOdDOY691ZOXB
1MpyoOdUoEQagSh5vCs8jCT4mM0/OO25EXpcQkapm/zRu4VOGg4bByla+CezG3F2+DmetEKaBLPp
gHhHh7CYsasZfTe6pGr1egcw7zTYbUvKSvNXAs5lZIfkpDB4pjztT9WARoqP5I89w2cXJY2Vurxb
pV5BWXLM9AJrd2reXopRpgjBQw3nYXvIcG+k6hDstOhoIO/zMOPtEEgoYPFptS8ieT1UcNujl32s
la2fHjsEJ+A6wk5DQNgnb9u37Q0cKUk1SIfTYkLJr/Ku+VpGKiedMlJEI1X/xFjecfI/A0n2iV/c
NXMr6KFZ3zsYN+wZUat0oUGTdEIQIrZLHzkVb8W3WDsch9mUCBbSRTHqvw4tlP93bjQksO2xzHLS
yt3PkwJTEDQiHaXC0qmwe/Cfb+2W668wxPYmb8xfPQtIuh089IfrCHVmkc7RcBo4s+r0LHRaJTv3
FkO6CRIO3ygSmZKRWGelTkP0hb8YcDq+gi2pNCiYR8XUrAHb/Myzh3vZby1RGYsVs6zrIDucR61D
Vafdg+rqS3h4GMAeZjNexVcZTeWmN3s6bcizo53E9CbctTz/GKQwgI6FhRwM3yjFoQ1CSrjIHtdb
GguFq0cjTFSp2Bu4uLJTW3NrpO+7Ugyey1YhDVEoJYx/rimIrE7VpdxJkWvFGoqiEqFcB3XDbP0+
SBkPYbnJJ1BLyoLmimyXTZxI1JCeMdfM47vPY2075Uj3tySGZwkKMlVSYeT8T16lF2b+WHH8Lzh4
kPr2cweAqcAh4/ikGAcsouP4CIEuvfnADRvtBf9B2vYg1sc/g/IUqPcfASLypIvXD+2uIFBzE8JT
8TI2COlhPYjGRx//4azTRLNgkVbkw9+9tW3qXcdRAw2uC5VKPcM03MeWgv654T2lcCVkMJ/tUmSG
UZKXtpF8phg7cGaOObIR8poGL2K6NeC7MAe8pXRMhdFGZZqvhclr0p3+O1xwLshLdzyHa1SDGS1c
h97M3D9kEZ3PmdYwZPrtGhFhdRjTVX0+JpfugA+IO8wWSjXmg/SuhpU+TesLn68lPM6QPqEX/xvh
UeoUku7j6QJTpAUOH/miK0q829+O7NrY+i3qqNMqqChckZ3sA4vMqa+CkBsC1g4XFFU9Vd2Illaq
eC1y690nlkkElYbYEy98eg2GIGFQk7DNBApD2DNnPQQJBsPbzsR2d40XcZiefC3leo9X6VRoBggj
Pa7wIbHF0g1bjVSNOr77KcJOeiJmKtfMcqd8pHu0EKh9R77ezCZVXs75x05nqCxvTMEuUipWN0WB
NN30I2FoGIX69PnPy0OhKqLhhSBritHXr2Jha0AjEBQ28tILMxgtsjW5Y/fls0pYW2bq9YSeIrEk
tluonE1e5/QfS66tmIVe+BtBE6S6vbk72M7uCmYCBEHKoQbjQnjXn6F+rgP5QBVqR/5DvbmrDoZp
C2SRdybj8pi/hv9qxAUrMm1ANwCnRV5ESvf9gm08t5c7eHkQGqn35E7Qtr05SO0WltogK+U1CUR9
8qdGmaeDb2EDLpIAfIJozvmO9OmVA/3LKD88k/TLmo0mIFSgcAbIw2wsahd6Poi1nkV68UQ/3Csd
uT6HXzzML85rvZ3KWX1WHu2RoQ9DaQY95ejGbLd6ttYbCusQBFX2tW1LMkB8c/HxX/CsH/e/iaDE
LvPHkYSPLxseNolncNbOBwkrckMDV5UxCFWBuFn+zGXpB4A+arQMf8r2X87bUGZVcrIkS4fwvs1p
EE6zPXKGKjU/a+X0M1HhCft57HMY/nzx/6122BvnEgiARki8ZeGSA+fU2Pg1pLhccZ3ywAvCKq2l
ZsH9GxUsQWawmmZU0u7EQkWfswgyeay9z2KsOyvHFkU6N0vk1Iakq12Qm1PeassVs4Vvjy31WFYn
XP7Izczhw0Cg5hRYVbmSJ+F69/Xz0l+ppBd+HY4TWEHfcPV4IJvVSDeTcYb2aW6nxQDCM/7nO5rj
eeuPvHWM8JQL7U/0i4K0vWcOWRIhvn3flYUvVf0dJxAF5RdLsuWH0x1JKoXV7pO8yxuZ0Zm+Xv7G
4CzL9aQqygWAnV5wrcs2AH2htjrZ3QlfmD/XYD1UmxM+4lPORaIxPnrnnglKERZDLmLr6j3XDh1L
fA0ezSiGdcVwO5c6Ftkgtm5859n/vMe1NF0i1Swx1zBCimXVcclXodexY66wgTBXjtYbRlMUj/1/
lG+HwpoYjK2gkaDL3DMdkKJoqpzCwAj9JxyPPhI6p5Z6CnrYN9ahrfJWRvbZi7PcUa6N5H8qA/hw
CJPWdTvw2icpaPrdzSy/sxVnu9ARSwXPFIfUR6wcXBycAjzo9V34MeZhSKtoS4k2XjG3vxTX7Ez3
PynWniW8cQuMnF3Dtkq3t1jlOfwqYpqN+HwgO3aykPOg2HsynbiLNq1nL9JOdvL00OWG+oZbkB8d
Avc+DQrGVkDN8lwA5Y1mUpBXPcEC31k+1h+pA6n34SbSnP1q9Ox9EYyv5sWqVtHhxETX/KE80z3j
JRROS76EpvHDaOZ0a+zAWzT86QFOTQPIiFQm54ftgCRmZrm+d1pDuqDpWQSBJ+ynQIZgMP2oKWc7
ByRLQHC88yvGRxjWlmifiD1mKTWzoCiVRH48FW6KsAVg9A3sGu17MrJEXJ25kN+BhyRYpmDX7vq9
IaVDGCIFZ6mIQJmmrx0mOgFyafX8uqnVrsyPrJ7F+pyc56Xf+pdRlBkJlJQifqRuqiL1fapl5l2z
9Gz+4Il/Fvc16CP4/NZOrcI8t4buitqxdJwyNf6kHEXY1l49wnKbZgo5xWGLgwDb9NboNXghtoli
5AKw8vF0Rxh1K0dAdSRzk9tVxX6yttCWwRlFHX0pU+YHuGsSPrzRamV2RfeR/ItUm9ULk1s/F9sV
gHoyARf8zTzV2W/WnPX1friOkVgfrPXWkiOcixRx+cm4INkC1HOC+Sp6QZ3Je8h63NktOaN1xLkx
DXKNzh4qi3m+W7OCT6kBBE0FZkdU2o2NNs82O6VnxLxWNhv+BPPAX5KNd+W21LNlzxihTf/B17A4
ZKutR0KArIuw6fWbWLWQs46VFDsNxWC7l74zxr6gNHtYWIjHA2Uk7gKNYpkcmdI3hMoMD61LDLpk
TRJPPpgxQ3dPHMrAWgqbIVA7npRUdTTJkTGkAd/u8JeQY4M1CauAeqUQzGywWLP6KC0xNyUJP9EM
75PwpSP7pfoouKw5+NoCiTG2k2wF+P608tYd0+Jn4kkI3mcWt72Z4K7LosIOnJ7EnS9SWKeAcaHu
O7N82MDLlb2k/JFgAd7Po8b3mUr633+APO3/uxxMvSzqUXzywpE6UNk60mbLdlFi5FP+u+mqJ8XE
uHMgE2dWRN2+bML2ZBKtcoWAdJNS2y3I+CN36u0NUGnrMxNl6c1mp4tUajVlKP/fHswj3iL/2mda
HdFrYwi/lUhPoxvYAouI2rzv0TdawVuyDc4jy1ah0bRkyIzcfzVHjB8oGGAAQ8CX3kS6lxx93Est
yksY+i+P6t7RyFyyCq7NgN/yd73EUhBTvJONEphwBecOvL6jy3Jlo5+Qz06QxbEvJE2Yn/BGzIJu
1kuZYcqM3iHa2g3ndjBFu5caNqf8Ol3WdHgcRg4N1uMDDM5x3ddkpuV81C0OsU7uKifnRUFW6int
7g9JBn4D0VUWREwfUbzWxDXFNvjxCqtM7wgBNHZ1Jmea+CwqToDhomj62t43Qx4UyoRbdMHXyJor
sJyKtQngqQWMjlGbcL67TZlvgwL4fYn3foz+wSkJYuNl58/8Pmvi+jGvDAmjkgEg5qio/HZCwsaf
VHPoAIRMAhEsKhqsIlbeYz93t8/5L+Uifw48lkYqqV2qGeck/OXAUmvjIIRSkxwWQU4gBZ4OiWdc
/5r6V1RRQ5kk7h+Cfqi4CQzA3lhQkAkoQmGAm0CQo+pT7A5azc65SOQmC3urm4XYiC57FyvGxRBP
Qztj7M22hv8+b4QtK8ZAq+y7oD33oeSBdhMg7B3bT4MvOWu5a9qAcuHQxVQXVDSi6Ue5XAgBniJi
VRhRjFbgS6HaNxY8sxnKkXlmYAY/ZBm128tQqBkWozcsYdHlQAscBjcah9CEcvv951NDhlngjLMH
VBqNVSOgOuTerOGJ/ix4n1UbkJoTHANmycr6msiV5TPJbfiFIziUMHtyr9fe1fvXpwsubO6PvWYh
Yk/rKOYbTobcjyfALOW5p26NC+VHaTkB+yMnAIVPxT7Rc/kwyofyq8QGy5gg0JHoihISJ8dVe/WV
XeAN0C+GiYV84WFXxAO2mKoNm5bIMafybxVDLQneZ+rJGrHG57G6lDw5fcImDqJbEJpb4CC9jGWh
KWf7TEXeEhsMac1/zbipnx1KhmiKNn1Qob4qtqs0lBApX7tim9Rf7OhVdb9bZ1JyDhqFCyJnUvXj
ZVrHB3wxK7/D6FglCKA9QTqcZdV+qbCyGGCskR+UlnbIEKFmfrX0wj6pbMSLfYNV7Qjt7LVKPD8V
89EcKrcL5YosvHrCbHArhDnJPdPWy6sSlBu60JssP8JV2HEmk6yOh9PLQVzAO3qJ0MXJ3y3dOt1C
kcWANpgK5+sHO8edjOnkKqkyZ/xxBrPoxzucFJYZ6RooLi7MnnvKn3hOKFRrPzo9R6G22n/wzysM
RuD/QIu3KCfDZ7c3oqtPaJvK+N6ob9yxpzz3rILDkBc9GTA9ZczDXkZvCM9cTMIfJLXGHt8APcYh
6RPGGTc5RmPhZ9J12+ypOHtB/dGn1wJyJzBQumgUyHr+zht+iEoIc4vgZep1EnQMlfmc76nwI2xw
31aBiP+ejrObhBDRWwnliR1KY0C6yV99Bn/z2oIABCkiIrybnIsO8OKf1XJZclDPRgTAA9+w3wJr
6afRKbaI4O+o13JI4tOvQfBKk0jJjjZIL/uhyE10mmLyBVwYM0nSdfrdAJZNvW0BXiGnFa35ezy7
v5Cju7gnmTvCHzcfvds9TG+yeM0tGui2Vo/OpHtehh4Av0e/7nwuQzpEAE1Ez3F5ZFjRdtWmeD12
CI4NiEvjcrIUxBMKepTWU41svnxdAl73b2GeKpkpl67vtzW8yrZgq8eeaH+b9JdguybXzbzj+p02
Rf+8Nim9v3JQKs75OmI3t/b4/hcAJDCqykG/XgqkiQR7Jz3Re/pska1nluxDqHbG7uABfvSc9FUy
XOXmJxOuTCESKQkzrJIFy8VobADlmGOfdy4ePzIYo3X/76bnNGz3EdEVoA0EJd3SxIyWwSae8G/A
SLpcaWzTrNmkU913dYUsDbKlvJWqAigY3SVpbNtBMeP41LoP9xQGtbTpocULK+UIr0AtCcl5P1po
vWha3frfoY90vglAB1jEsmWElOFlkS/6Ttol4cy/CEeXkKW61r23tGqJ7cvc1vXpuBBjtEglq6Mj
1lFqumKdhY1l0uV90q+dJz4tWuwtoYIOZ6A9JqHLQ4B8WjOhb0mfiMvEuIl7wZCQOHcTT/4/8/ne
l4Y1tgX1/BLhLrVQpiGpwUhehJwd8wYFgooXb8yJY19ytb25ePJ64ocXDQLDHMHESYNe/IcWjhzm
2VmDBj2h335FyLP5Ou4HTcOLryImN9BAP4aaUscIAZh/AuoSb+Jom+jJaMAjVL73wl+kfSVcipSQ
yzowoPLfrjSl1uqnJBv2G37BjrRuYsxfSbfoN6atzRfJwAxCuKctXVZjJo+ipY0jskeHKAkXQsBl
Y3jhf2/LRGfk9hrUic1pVWM6evSsENaerIGGEXyAH0stfVQVVMMZyzjoxHo9/l2lr/LbPa1Q7nun
2QGh5tUqvy/HCVFKpqZXMZH2qbB/QarBgnooib8qtrk468mAxNw40q+t8Lwfs34wXroIYGpTGj+D
/vl/w+LKZwhzEfLhr4j5rHhcdbrgY5KYDYe/NBxPQHzukyg7+OwBzuVLWl6wFMBvHN8w4B8melwf
L+Y3r04Q9CkNPMwCdSvpewXBEuQ5LLe2H//JXNXl4DVLXwDUj+vT4TJeG8ZXpMqXw1A3j3yNmcGE
rVwKdrrM8pbm4n/wV/Zzsup2aYqKm5WOgAAx9rhEJkfkpjYouGflHMWMOJHQU00ywgy1GLqlpr2I
3JawR5u3cTlIZX/G03LflhGJif/ebRf7ixu6L5UuWiKmh5o1qlH+3MYhup6TV3Vi3tPKfRNbO58o
T2K62ZRh+JHuDuWVatFeOf51y8kB43rTLuuoferDB8xSIiEGI6mlBZcRlK8NjI/ti0AjxcEdi7bp
rK5dj1LhVyv7HSTr1DUtiX10UkWFs9s9ED73ftNRptJgruzNwbwiQy4FcLDn8H/PBysY/ptk3Fu+
EQ59kGi9qm1iiKABpTco+Tv01OziEwrA/uS+joFLE5TNsZYyfj3jVZA3pld/44tazDMYkv20sSvu
sVW4LMk5OcIFyIf2hjAbxGlwR5Su3TH5h/AUljed/BclwWcaSfouYge+021f3HRx7nAdxmJ+tR0v
O+erJH+BBgSFHm66W2FHGBgwRO0SleLQLbDC4inbxdAzEZ0QPDGmJDJY16lRqZl2s0gPC9em4Q72
YypaBG1pSXcm0NWftiIe7Eq4pfr5uz6tmJcuyrgj0zOKqhbBU555oXyC8/M0tEBseWyJjw7Az6Z9
8G+JAmMpFSiBMS4Ee11Ow0/G0cXRSjfvr44ZrwsmFm8DVM5DQhpYouZd9vJdmiZxDUKXxkkSMu7+
AyUf0LdnqqNyyximc2HJbyOEbAsY09GjIkTViV709nJQ4eKEv0B97cNVS/XwUoy8sAzBAU1Zjdqc
4uKRdN5LRbWhevU1PY/0cYElyQ0O6Wfxu8MFgsWBEDKBjUlolV6tSnfun5oTIv2a13RvgtchwRwS
dM3EFARwijay3K+dy6313SJMTonSW8A8+9yPvJTXdOOsBxXnrR7VLb2DY+IalOgvM4Th4Fo6rOaC
b2NC4e3PL2rOL3A9+ZjdVI3R+nuqfA+dOFMNsz4gi4GIRtREXLqS5BhFQzlk+mcetHEOO6mXwkM+
7RUWOAhiOmeG+xaTe+tbZGRzZaCN1imXa4Ttbw0s0n1vK5sx5kvyjY+CchcbnMilzEk3JgY0WlcF
IGvZQmGA9kR/snVk6UqzQS6aANQfLPwfkwN5v7178fU83wdObYOVIbFJ6x8vKKNTm0ntuXHK1IYl
891YKfl3wbJ9hFDNBoWl4X9IIW5slbE5UgT1BnoJQg+RIlu0yu6WBT813wr+TVuCgMWzPX/OppI8
FvlrBuqHm75C5sorR2XNuwYCtTSwb9pM9zod+UquWsHTJHXivRlXzIs+OzGYhiTz/cAx9Ax1fI6B
c89p9cIMBzSfMBIsiXJhvjcBpJaLLNK9tV2L/lHicmfWfUbKoLGHJz+gnrjNsnK+EhompYep22+M
45TdjoZktaanUeYewZWbbGbwBMLzgVDW82TowHDydG8fBh6DN2Mu4YKu9PZlDvtLAxCYkJo7SzOq
MbMp2ULDNhFU22ywPMMygGS8p81BG8VF7QVDIuMKkgWeCru/cqH132s+qenZ6nW4j7YXsE/sUknZ
Z8MTpu2r2/+D/SaI9thC34gaz02MgewxWKwPR7xsBJapbDsjneJtYj5LnaRVwn3B6kERuzo7lH9m
Yf3hCdH/eMYke4nsGkR9JfvmeYlH+F1ql9FX0vvAYVDNC2aYUlIaeYkzmA5TjFOFwy9a+/abd+qj
EiaZILgviBeuilsT8CtHTJbAcqH0e3SDWKTiWmuuxrj9+uSswSxWZS87Vwno+PJpsX0OK1MBeOpj
R0qQusaRsteccZfYSsZvexOwbUrE2Esin3J1J159JBT3esCURxGNbKTjm7zQLWLZ7lMc/Vqwb9+A
GZYslnMpo0XKn5IkbtnLnThwFylxANx7ZaQ2vqdpsQrp1nOEw6MtsfDqquqJA26JM8eqXTESb6gb
/ZhIjDDdn2Dn8sNUQxelOHw3HwZ7q/kWgAIbkvXQAM4qDHKsxFQm9kWKhYOXyEk2LGgK+h7qL9d8
88dUGR98ILym3moRgzwk2QMf4yt/sdEVK67auiIrC74EXQtLHygc1fJWOBf4paadbHgMOKnXCzwt
8K4aH3kw5E6j2hu8qGSegApDM4PKvM2GCRYEFFu3lv0NIbDjZtStm7j30+iAg6K/7XdWg/Iuc+/y
+NLc3sNOX2ppNCMJPSDv28GaDMJ1H2QPEVN5XHuVIAzOTfWmAaD7YPOeYnA6OejzAHhDpFtgt0gc
3bA0rhHlPNsUbO+CZXj2pdFrLZJHKhTYK7Vefmr1I+k+8zHbYvSMvBBSQBZWPHVorYjazDpbo9Gp
zrffKQSaKWJJRG15c8ADjsC+h2PlbGCK5PrFTwdbleIdUtvApWajB2EZjm3+tKbDzikK+sZ98ql0
hcsSusIo9KzXHCXogkjSUstIgiiK4rklfDuVaJMvztp5V057PNz4HnBiDz0YLVFNIhQN5mnDjNqg
31i5g87vUgu6spHxpbEA57qk8FLzHy0i/JmfgvC6vY/l+op3Ne224ny8RfidVXLQ7CJDeJZNoOUl
2fGmhio6UtCRiRQxUg7Yty/k8QJSeM84G0XHHSUSmxFqNiIn/f4ZkQVW08FkysfoUDg0QMOT4vtJ
Y8ARFFZ6sc9NIllLnmbDnLkWC/OqVmZ9wGsUtEi/Lpqm9qhYg2k3f3bMCG0AXzTiv0mMri3LHLr8
hp2PeJsceYMTlJB/rRf5WwlOai+rDL4xozkrNquumVYvZNWXtxEl4oxQ5fPDl0iMsru1oyhFbvWN
xaOzHvzzZowqNn6DBqNmUYu71OxFoak/9XB8Lz5qtKP9Cm4BErPy8GcOEfCApSSl9+5Ck4MJ49cB
Rk7cOTKso2lsHIqeZfr8Nl2oRY3lnwPLYjb1TXd4YP4lK1uR+m9gU9fyC+QxmKTdoBUc7iEBdEBM
HgBd7Dq06XxPeA6hS6c0NL181YQbtly7RlN4MYcT1+bw2OLUCsNvwJRL7QRbxv7Bb+PY6EGq/xjc
HNWlX46BGZAzc7wgQP026dUPszmUJ1mL46K0VjoF9aCe5YykIEJguzdM7iZVgxa4BOFlDuuSkneo
DX1WEMxFp+Jh136xNCIrXDOfkiD/e0WvZZDf9YY1auO8uY4gSpW1aw/0+/K6H1IOaUBlihjeJL7B
OxX0lZhan1xxAOZS5b0x+zbYpx/3B2FSp0Lv+sTaDE0GBpxdmzj2fTmpQaek7C6jNVCr/8Ab4tD1
KgN3Lpdc1OGcuw5ToHVFQTH+fHzOhD4UG0zeDDRcj6L14T6ihon9WL3YIkY1SMNrfNHcsYXCRNnv
sDvf9d+NQ/x2GS58/V/LuC4N8VC8xZ3vI2lP7nKFz04Z9gjRybtEaOGjFT0YTEdp4eKW8d+EczzN
FdWPJp0nc+Jetez9t8aTwN4IVWBN/jhe8Jzf4fnUm9IowiTxM/CPwHql5X//d+fLzoqyFbrghCes
LHsH6t2IDh5pNNjmK0ab3dUYwV5PVsLRr6jFIEuH1dF9W46BrBDSTeueINl4pUft91xH93qu8Fo2
q7Pj62PK/wHlX7H6/viTqviaN6gHZsS2YUuO+sEy0fZZCfYEMpFKj5qRFDr4Sly67RwzRH5NFG07
w4fEDnbIQ96S/pt73DXMaT/1kCCJMMtojjsoihMYe1/hnQKB9OroS2tM5vAIY4+oXVsRjK53G3wj
hGM04DxrJTUJf6ABsq2Z6ocWQq//lEq0EIawEjCUaXHxATLmPTOytZ/SCOeSg7R4s2MIzsLSggDM
7IKhFAtYnlYgxDLjqFSa4UAzIMHsfIB00PqfW5MqelXvqZENcOgBEEN+lO1j4trDQnTpVxaNH0hi
aRvr3ZaVD3P/Q3DulpwNgrZnUe0Na+bnhZIhHx7yWXXlriC7635VY17Z2IWo8U2WjKIaqMG5B9fW
2FVZ1V6booawstzA6XXUZzlFjMPQoOy2ZCuUi1+fOnIYM7WgcwCortWNRQtpinUWMnKMq/d7ohPH
gxJtxzZL43UgwsCh4krbhj5FVrSy8iD3Pel0jBD/UOc1goyAG6/6NIByj7xU/4YzBwf09mtuhK8S
U3nXp4LI+r2fSEP1TvReFr4Jl5deLPqwWxHiEt6mc+PXj4HyHgRvhDvyaQ54vO1+FTo7bAajBQaG
Gaof2W3cVgTJoeKU4jlu1+UqalmVAUjYB6yEyo2pIQwNuSw7knWzoeRcrFvNUNnv/KQy60/KdeHp
VPUMsvQCSgZL1+XBS1q4YLKRZj7MBbACrFOQ3lVbMuEmUeBrpQia6FkNQoVRnibFvrtI6UV1IIlx
oWiI6ggthIbQaxie0gv+MS1KaqFpz+mGekZU00AWywyfZNawP/rRIOE1CjH7EbdH+0zRaEhqIEUC
p1B3Q4a0lx+l5KgydmEVNNiVSqGFXX/VxZXMpZDaSFyrTbynkfASmyQ9ct/5CNSRtyVqx/WBF+CD
l/4gkfRev/WcgI6hiwA8auvVnwP3AfcriaSa5GKIta91/INsLWMeW6nAlj7VBj4azPy/z9t2xBaj
9WE8AZN7sld/2IkvYJEqreYsZpE2XP5PmJgTMrrZ0FrGul4d/+K+VdXQqybcPvEceegZozbfOjlF
1zTlckDb4wA8razD7ykRFuIE5uAdf2DA5BxXjYGHTeYEBEvoq20C7eDVWlK1aRfDebRcnzn1sLqj
dGsKYeFJ4BHYVGLagq4bw9diHoL/1RYov/K7nm3GG8H8w660vzPbH/elW6S1EMAxGUE1whI06TR2
jFDSfSKea8ggjTzPg1Sch/8byax1L/DiHhJlEXFJ424EIr4arjTr/K6bu095/oZdB+BvfVgY9CMh
nqMOuO4Br8649qlN7LAwfs12wn114Xr7bqqXbfZcmohVX1dP4m2GuadkctfgSmn4y0aDjNXmdoP+
jrE8Wie9YdrXjfYOJrXvZu09UchMHnrtHKCwRNZsQPe+4shrJEPIzEZjCniciHujQSD7/0rDDhhm
biB6LZIuAF415z61C+IUIJ1TJ1wIR0I+o807FvKwXMxlaWmOArv4lBEOZw0+toInfWEOkv3IQHHK
w40mVa5KvqST1jW5GshzOyDgZuD1lmNV2bd8+F+HI6wQ5Xj7D3q+pFBypx6EDFggMhmNBGS3HZ1a
tu2/wEs0Oyxfq+w2VqGkUEbWkN2WfLvkxVN3vwbD1wQno4lkXrV9IAuBShlUjbo0bRQLNs2XacwV
G/WG5vfT0asF+ElS1yjHhYWWkd1mLDIWBzaH0FWjOMQwier+3+nlj1VBmZP2Qg6lMKl7B+wAsWwM
iTaYU5hrKQN71sbgG2rHX/uXMk4iRgm2uHaAd2A9r4GEy2B/gZl+4uTNOEC6HoRkhQsiZAvAFeiH
gzLgi5lDX7bhMTmhIS5gkLGOZqiXSgGTGTUXvfDAOCFV57NlreeKYDsYmuryCwZlh9tFeze9Ax9F
8svjJNBLampbnpmCLQSPxWAfLx6a79cObYKJjYJemNK9nk6szE1ppuC/xG3WYC+rKEuaCAAoR+tX
AwRg1joUB2yMlKjDjMCyi3zl0ZYR3ZTLUodLdIK241BrsYJOZdXltyXujs6NeAorF5ZUo8wN5/OS
cnD2B/k5WI+Dck4t4G80GRDyRJtMSILI2HTiJP+o9Yq0sUnHtbiQKC6nAwgxLK+pWp7W5092jxUm
xyU1xNNy2OREThQmbWe3xnUthA6xZjEndA/pVGzU6ixXfzvhMXIpTWpsAc7TMoXvWKoz46qq+4Gx
HDDaOXkdFa5W/4h5PW8nQtOxH40TOAMQZvNcXF/zsfi1BN35G6J/rLEfsLTYR5aa5BDNurD7msLx
1xOLH4l+3bxwBNXpZqvrQDVQr2YPcadsvRovbOoVRImjKMkPX9xdQ/+MweYEsSu/2iZED9xoyLAB
p9JRjbwSZ3rMC31tdc3zojGzUikoMd5zx79SM4vQGUdyIxHK92muXByHEfuZt0xAe3tNJRxYH2fS
fUdK5Xr6/l8pf3IGRlzklSKM2Gq6C2CAqeu3tJCtBkUA1NwSWykPpw+dXXDBj83rSspmdrgxRMss
4CMh/36dczu9CratJ3a8cCaXaPdDREAHF6ENyR1urqte0DZMyt1K5qMVmr3M6p/F3gsrU39H1RMo
5QkT7lMDrisTQNngytwIUXsnhzFjZ/bBVml2m1H1slSfHKhnegdaZ3+2RC30miTKcYUcQd1TKTAm
LKZQW9Lko98s3wGRFfCmMtZWhAHGBZCVLf6uTjweXNCZZKBCsUCl3Jh2rsGp+H74xbIG9ohu6rEd
8hRha+ZFisXH6A8R77uwheVYVHN8TaZBNhxJBMlHD2POmlsx+BnbX8oGOK0GKYAllY1Nof2cwOqd
G5CKJfWAUNgPeYV9FYd6/602B3mtAttY8FRrjAXBBq12Fc7XbidUfOUZit+K0NXPr/OvVw31Z3py
Pa6zICvnABnHaEGdwV6zQ86o5ydqIWzZAsvauotJSq6doXGXlnt8Sp//RG+OoGTd33fIqKckI7NE
f/roBLoODRry9imzGZu/hPRXN1ZfXUCKlpSXhc+3R5fe4Z0l41sP0xArD9gSUrQfVmeqaF/iLsNW
cf21dxg4grvqPq/KiZ8jYyV3bU0megAhm7w5brdEkZZerMbdcYp7d39kLyk2bLefg8jT0JC9U2qQ
UToOo2DBQtslTEG+zssKoDnr5D/m8W61PzghORaga4qkKez9VwSr4OMR/o5T/NNgyScEX7nmsizf
MyZ5tNR3BW2kEOmvg6pbfrQ492dBPcbvoms21gK4G92vrvwdxYtGLhFOp2FHPjY1yBjToZbjwMQs
sdkfhCFh2MNLZUCPuHyAOMDhVs+P7tRNoS8lenoGzEsVv12E9fQU8BWpA9ijaRBQ7b68SxRwkUn7
3fh3RJjSYK2WAeDJP1LC8Vnksiinw4rP/Gy4DPjhs70lTWGqtJT4j29s7m3dLmrgiDqrXWZRqHoT
iovA9LQFB/zyJcKFRaa8aYvHANAzq3EFSMSETF1M09KZFl6eImMb0ulnio1uSZ3wFMWwb1RllOFS
xW5Ih2/aUE0YZdaEnM2Hyx2l5luHpXmvb8VHyAJQtoJRSR5gNYq0w/GECsWjDj+TK40ufd1B+9n8
RNt2fYvl1RSQZKNpa4YakDKJ3zK3YAuXuKhXS8WZVIl2Hc43yTYr6YBmg+PJUqyXAv/c28bmzAMu
o9ukEBK04UeG2q+iJFXeyFq8uekhFgjxdHbWvpg+jCUpsxG8GbWu44rOkLEvbunlTBiB0JRR4S5A
ug9dGbPyEgLOJtaXphonN4OJW3eY8A6WvqGBth5Ph38zzd2tcrStopXHIox1owuI2ysA3xIZstE/
bShE2DEQfaov3MIiJZwyc6P4V2ssuA09eM38VzkFV0dplZWh2fugmI1NzrKMQE7PDDs3evsiTuez
Nn26M5zLQIalUDFDqyVHrWREx1B+lgaHIahgOO8MyhUWls1askzQeE1nMcfew6yJDQHstqi29WR0
SEQ96LCYfWSBYx9nKi7pNtACl/BEMFrKpigsPoGap3hNcglNxuOhJkYaD+odT1yenj5FWEChAMwS
kPKdYf/usPEsx8CBYzfxaU8xm34tokepl7H0M5IAMv8A7MK0cWqeW2F+2tiZ8dO82cGeDVkFQ8uQ
e1xqZSEOivu4rH7Z/S/Un5aX7w39FMJT8hcC5SB5WVeZZSs0wsbs4Fp7jBqG9P9y1oOt+wn6jf+z
d6j6zzTGmx0wZcGU1eLfAT4hBgeMRmzmr+CNm38d8q4tz4F3ECwoAGtQ8tNvGdCFruiohk1k5dg/
8JMM/UWAwC/Bdf0X48hegIsI7K2nTZlMuuU9a/rtu0lHnWTFEjL7+k2V2Lt9WgakAXKnj/PhqTe4
5g50zu5iMTHCk2h0RAqsXKNXo+n05DVKAfxU5V6hhxKWuSu318kM4eU6LFnPJO2efImzVZTJlDcg
6fEAbMt8+748atL+a5v1pwaZyc8fHX9P7Q2VUCZOvMTE06rIvSpv+x4pCXkakl82XZFhxIxDC110
2nX5E+Wgmi6XnrcqL5/vslPNoqZXrz9mmlgqyN6G29cYfYxOr72PkcbHs+1obUVvbezAsJIXz+QX
ZhxjyQt1eCBbacfYjMSXp9bNRhR7qjqFil2/zS1GI14wv4HywdM2A5UlH07AUGFB4j+q5LvMX0UV
Ay9yuhfOSSmvM1Xgmdrx8eaHxAFWMIgE3j3xodJGFWwlOrkkHsZlvsGSqCsmsTRAuIAN9APm5o1m
K63pVGEVgYO0WVffrIUysdcfbojsy9oI3EMxZGmNPpNFGBv3ecfuYG6A7CpCdO7N5sWG5ZBbueU3
fJ5aq2N5HA0/iyAld92A8gd2RtGSnJFGX91ZRTsk6cpw478xLF0yqOVOrV8g2mXC29iC3qFRNX78
CW9fE9f1BeOysBE7/i8VXEiHhzzQnTMLCyekDTcoOkXZlF8wz/59qGbTbvGQbGuA1BDaVJ2nNa9i
6waZ1U7q4nIiIcn9jkw784Nmm9nsz2Q61DVatkuvPv52zfRYkBh3Z4XvfCNSypcFlmbVOz9AG+9C
Isov4KCOZ5feK+BUOzu9U7LpMz6bvfWyg6mS4SlTpXhrr/KdD6X13ktqRMfekcDJJlJQCTAxAYDv
DVl8FzGs3r6wdqJRKAexaVi5T+TglQ5uLmGmDZn8piLDnCStBtAP8yiN7GfYKKHv+JIMaMGdSVkf
NJG8tSBlQ9Ic3Hkawz5IsLUWOKQrBCAWnuWqUZ0tULCDNkWxC9qqK7j6bvVFBIEdHSmEf26kCncE
brVyLbtkAoOnAA0eGLsKjyBiAEQCTEMKacGPpZm0uf9nX8E3hf4nB4aI77Aq1eo+r7ovO5WowZFY
6pimiHrgBjCet1XbJxXFRisosxWntzeLuGgv3qmJqzzI7Dcqt/gO0Q58L8y7cz7DIn0Av2Zea1DB
iAJcULLJ2tz0be+uKIYDxzUlTNdhgP/xUp3pyHebzIrBKphFIEjUwnQCVZjyeyGfbc/90Pjjy/sU
I8dpFYBkLGgvMPZkybVsN4j2XfA5BVPv4690fFsXbK8S9AwHk0ga/F1TGg7oaprus9P9mgvjh9rj
E71d7CIhPG9af8qs9f8fmGt9Vaw9KN7IXbjRHe65Lw2wicqWqly49THmLck8WvK4EiafsZHkfcNw
EoqlcI7OliYLMPnnSVcBUNwfPy2q9qVy2ehlIfRuVJPZBa4a4q9dPb/OpOiGLnHPc+Zmy2KJd0SF
JPM2GXghva7stQQFgnI3AsVtv+3RT4zl3A9eqWD5zM7d2WnyOEhmCvShdXz/CzH8b0opQzW4Z9bJ
qQfAo0pjTfeVm/wVdtX5/lRqfUAFiHKvLJGEPCcNC3Kphy+R80c+1MTeI9hHG+/HV8pQ8OuYp76U
jkVJJnpaSETY32nepxwSyM3pBcLD1gqd7WvX/q/9pQObUlCbSePImDiAY7kWq9dQtIFKcTmXelU8
AheLCCmmHSt3a3lHPSkktT6NxevoG+uqNxPi+jJl7kwsis6arpAAERDPuxP5e/lXf4yaFL4kiael
INekJ7TuHcjYJbw5kpy7STAoX0ZaIl9WsviWjIaZYgeVSRE/3Rxv6EFUKBuo8Nxu3BSm0a4O8dPb
KeZrs5q+FlNvCHpoBlrEsm0UKHn5ldnnEqhL9YPAW5bwrCniwwinitjB3OwkcPhUR608pfmbsMKx
XDh5TNdur45yqvKBjRyVt4nCwcofSQuT11yYxBa3h6rDK4yUPYhJYQPPPwR72uHgVVscndaPa6n7
BRNjCGBlvA7bDQjtXj0Nvt8fvEBcet1litaxvHsKL3kuBtGPknlCNhQ3ZI72zGPQ545Y8FGXx/7J
YAbOsT6VG/SWmASZmml/dOttqUScvOGmdajpmCM5B34tXEGk9Sd4Kmo6mP2GNbBOEpYkiePG5j8B
dKTrm59LTHGcbZkNFujgwzGUwjm+PWUWeFMeM/Guz/jpdJWX75Lup7KZvPlyO7Q2kjAhc+goi3NP
p+iGs3M2Wsp+/ahDFi+hvw8So1Gof/Weyy5S7ytd1jnH+/wBhNF6ur0pRr5gI9NVb6U1SKQZsc7b
P/ThhLfGxM7XuoISdKToMuqBMLD992xluiSwNOi1jZBo+jq60f3NeJ/2WXyXI5AeF3w5NEydANW5
UIA6LxfRWvsL00/eWCdQ5dylBc2QLRgbweN19Gz/1ieBoONPeC2VDxvzh+GIk3sQMz6PG9vrZC3+
/mdWYSlz6o/oUerMMfsRNY+YCK5CFZIzar4U1sWRT8cVy9c3q80fUyeD4KiC6xHh+Dqp6vQRGg8K
6EKbUEPHr00yMCPpk3sYRtHOc1qsELSdabN8xDKeBsSr8SGmZWGCAQ4zhUDBhKo4aZUDTErPEBVO
/2RAKk7lTo7JvyJ6mUlVMKGvVnMXQMUrxXKezyeOwRnlJlvhp7WGZK3L/YMjk5URpMcBkRxrJAu0
tBXiD8Dbw/Kp5vlMx64W3FOaD3Pl7xEz8cjpskO/DXMpzRTz/Lw+bqIq3Dk8mYo5AFLcErcK8lBC
P7g4gScMDVvtjD92j01yUk1GUGVp9sIj0N2f62K64s9k01ZCdLaLHtXEZmCSrHsehMNDmARma++t
w9pj7vnMA+bLw+YkIehzCIHVwj19MsWr027mwibK6EuDbbO7avZKXg8rUruwrHak9TR2pkGQz2zN
Akh5MNJeAhQrPkkzbJa7CIJq9xg7z4pxBZY+ewjzNw8VyKGIaNranwHTkEHFTpgObgDsLj1xgfI9
ZT4RW1tUqXsQ5x32PPdU2O8/OW8sg1b+YqBSqVXxSmyQFnUSG0MJ8/xIG/eYISg8b11FWwMof5x9
MzETNowIwQuxQEt4HdY/O9Jxet4AOFaD4QVOVQH36vTp2AKcFILAKMaDgwilj3aCD70GJrBKp5MT
+ArklI3NBNK6GZJTX/OMXeFwMQgE7zxlANksXH+oG+c1sIqGFOhg5DgTYYr9IT8KTg5ABmzNmr0c
B++5I2CGHhYALqrc0d/c4f2GlAsuTBiH9kFiOzneguyloQY/ZWGxcfzC/BwSLnMO2FM/qiXRxioV
ld3cL1kKOi/eV4czlp8auX22K/KClR/M6IIfz3x4h9i4+NXIepOq/1Bh45JTcFmvIL/zEA5ESJmZ
adocEVaEzM5FZ9mSA+9EajR6wHtaniMt67ZyF1q4e4Kt5tG7rlS2PiXVjGe4dGsJtJVY596VrypO
hiZ8xNeKCyFQ/btobP1Eq+Ownmvr2g8ySdAbFdm2lUyv/tQUXfR5wQwfFfjp+fiKp7ZW2caT29mW
5QgaDoxyWEwawEVD6WmL3AUCUdpgx5WobtlPWGPTWxldGRDzj4I7+15EYobyqSaWfAtf2AuAduOD
+kRfsVOdt+LlIBpcpqxZfWYqpNLYDWdDvVi+DYhdIzN+qxVA50odmMSBd0KCmLS2Sg58Qku6HcHR
EyrkaQSZ6kitc4DSL/iBK4ZXD18IyqAU5SoCY8XcmbuTuipGnhWVuxibkmvKrMwheBp00XO7Wzy6
DFyyCBH6284zBIoD3n8+00LkucHLnLB3FBHraDwj58f5WJajdAI4OlBuD3418ZrVFtbz9s74yCgp
YYVJNsoWSPrCX8wTPiZCIofgVTxiG7Wn+wkIEiLXaslPn6oUVgP/aD+sIAlveAYw3Uuf/GEK9z6S
ItMQytmc/uZLgMaVJgRkG0WkIMifon+YhtnUsG11fvEeemk32DiuhNjF51vr+V5oIxdj1KIqqRSY
YtPBH5hHJiAOpMI/yeU5AKiGL5cusgc2kY0DDoxXH5C3KLmEHB0D651q80Res/sXxO6j+Cef63Pa
OUVdm8qvOxF12utznISRqTb7bBvrRGjqDpb4jqEbaBf79TQx78Bl7MNFd9Z+uTzUbt2VgI5hLxHA
cx/l96IAYA43kZBvd/Oun2OmIM095y/U6yJAB6Taq7k8QapB5BpKkCyA/mBBKo38o4NztzHESSGM
ihWpb5AweMRXZE1+2hXor2O25gvdebWRphnaIypzoZIllhcGKKxc9te4vKcD14g49CUnCmjWIOPv
D25J7Bp8GOkqMOSbMGlVi2kQqfwD5PVH1QVZEDuRYJ8PEg5fYYXkl0IvZ64vso2ILgjTQ+19etCU
u9vlZASGuxHGPBzos4reqCZY9+j2ZWmi/9PSkt+RNs+XlhMKWLzxo77//2oMmtR5HxFKL6u28w26
iRmZrkYNVrLqJ+s+3hdfnu5FpfZmMPMNaznutTZPxqzgxXKnhFBaqIaLYmD1TsXitXLLipOeXPHL
L/rQJHbrGm6SMb0D/FFMSrYDQi1kMSJTxM5Ao4yjYaftEvaWbr1E285UL9WusXGhwPSUTFdkTogA
6AGl8fdpQAubFnfO2vQ8fKQ6HBs8ZvYBoKywI0NT1UPt3QamoEA3AVYmZ1GDhV97Hk9nG+p9P0ws
aoWr4MeZwB1bg8dUnrtyIUPESamegJLwlia7XcUP5gasw3yRXDTDRkGAekK4E4x0CdAPN/lQEQ59
+qX/jUZoKsrSkQQLSAu2rsuJx36C0PTNRR1bvnZRp5bh1rdZPCF1zhfnXYs0ulepdvViKCGmqjtt
nugQ7NYx+oem90LkgpH3e4d5N0Nrfq3brBrJVIE2BJNySGcxoRVLMdFHCnBVc/8KUfW4tiMZSea8
b2wLszUtDqA8b6Pfo2yKxq7FfvfreN5a33LNCbs9ofvq3Rrxj/Gj48BzriD0XHkiXugUI8O/5dV6
V3TXk2p5P0aOiVsxypC8Fg9IqzYaukpVfodTjNcZg3IyUQev6u7ftRkCA2MBfqB35Rx4vNl/u5Lf
l0Wq4sVuLCCoNhyOwYnR4TjkCznt0S7m6ZXq0Xq4aQEiKFsgT4BKPIc2soqnPu6oEGTkK8qBEDFY
CYq0aXTRjB0242NHm1maBSdYTZ3lFg/CpM3+c5FyyFNfBqvYmCnHLIgMwuht8f79e2SoyFaMIhbV
JXcmRRPR0sBEQGNR47OjqyG7j/7hAMYwAQHXjFnBB3xYOwFcghw4Pu/Dp/o7tGc+DO4IsMKaeHjq
mcz8LjmfGT/PtY4yxcTNGr6fgPpbBNefDnxxVPVVoEexWfMb/l9d2znzA7T9xyIS82tdyXFhp+wX
jajbo9Cz5tIvPOTO0ZSrbSgYNZyAddbHR+r2d2UkNCgm3z1E0f+ug3JcYjGc0NeS3QZt6ykwjl6T
+qoYNJ9U757LwOnVk3oUP0m7g+UzRCwvsjF/DMliY8cSs29+t4lcNeT3dZPXdNkyD0zSXEqEjZ6x
6dh2xIwzjJ/nTRNYxv1kHmMljHOSgzeRtNx4x9HfyJfXjt9v0Yq+gePspWCfTXx9wJD8sYKnbupR
GzkbawNOVEbt+6y9w6Yp2eqdKivdw+mXCRL+otzXamCsjJTYXm5Vcbuy+28FhqBf8Cao9QYS7t+f
UG37HVoBF6kk14R42N+uoMiwA7s0DpTY773gVTt+/CFt8eUhGVYToNeXWEWQBU+Yvnyrmid2fbR+
Lmv31MvMXpUbgJSAqRoK3Z+fTlJRVn3EaXG9jZKm0Fcac4ZbHTQdQJUoXXuqiGJm+IOhJpVXjLpZ
zGtUvse7gnFHnlRQFfRzUfro40QQFcFBJEKc1Yc8lRJ0VbpmQmYfZSlPnnU9ajP2KBltde6S/FDu
6BvVnjJTKVkJkv1Gny2Oz4uCdkpiTkPZBKSTR44MIv1X1lyH+5lxVX13rbaQVKRP/6k9Ni2rN7uN
Y30Xvi2ISXJq74D3ef4CHbA948Jq1GgRRTqg56cubXRGOMiXfhD5wYZNO98QeNdMPVoTyRX3Fgok
2vn2IuxXr+B00aCZ8BhLJugWCTTYAD8y6HcQJsUHo4DEiJvPqRCTRJOWIVGSHRJR0Qakja0MOfaP
tm//ei/lv9nhJ5ngAFia1eLllZrHT7/ug1HMKFMDLODfK2Lh4gHmMrBKK025uNgWPEvHe7eqF/+A
wgnhW+jvwY8plQG0MhTUHzewaMo2yIZhNVg9/ojcne+j4AddkUPiMSBe7eYlO9e1saDiq5jDbb1E
zNV1Su2YArt7YeIo40U/APB+38Eap6pMyWSihWeszInuSAeBzY20bbOIj8CFhFjXP+vlwAql0Fw7
KaaCSWqcCCqTy0cn/fkZaNSptLBE3ZyqltZzg6Uh4TlC5KNdumWuKYEazmE86boxDHKsAXuN3K5f
fMI2DGvPG2FLSoYH2ivHhgZJgnvn+rz29mnQjzmqiYvka6SLPDCBddjEZRPwewxhn6eiJE7c77/l
q2TZCn4pbv/3JO6nRq/rAuT7qSe0kXkxNNZPdv/ZbMZMbV3nwlWY3rMiS0F2omko4VICALd/vALB
DQNzanxqfrX/vmNnHkGUaxQzzpSudlX8H/mH+dNy8kEBXoz6UatFUzU+yWu44/Ok3fiebJKpMGNo
HiVZSYmgYk+jEW4qdyD1TJx5/pohEIXQfVUN2S/b7Rb6XZK5Fk4BF2YCaI0/5bahDZNC2KS0VXZw
VCBjcaMSv/PRWNJUkbcCdGwtqKvOBYbwYPiTB5kd1z5Qa5lJN6BsR3IDJTjCQfuSGMGlKRXcggW2
O/wwxTdN+zovBve7UTpX0ITw7x/FcAsv4CjDA29mohGmxDlOBotHx4lWItKZbQ1kBK2yqlilXDIE
qV1md782bm+Bmc/J9u2gVKGY0nAPY0IGzowQrCsqgW7jY3TLkrxbrJ8jXlgyqkHa0fId4oHard5l
ksTIylrIRAl8oCQFCUS438eofsCFBFtYzNmJ2DwiYX6CUjCZghUgMY2jFJQklsbAk6IFR38LnB4L
fMgSDRuqgmvd+4Hy6aHYpHH2p/lmaISvxbi1ZxHFiomgnHFUr5RHE9ZK1xgA3MdYN5H3CPnHP9hs
SSHq+rwuq+KzKniQamEtS0ZoZ8mkO6QcSFWXjfyI6zXz6d1eFREAgj1KaGnldY2MssM7mI3uWjlI
sMzu8/uhpxSt3JTgrwOyys3I4czPjr7Uhq4sYviPBC/po72lbfxeGuc6EOKXrr6NiRPkCD/XMOpq
n0cCKpy4up2jsxvz3bqlQD873ai3ape1ee5kvJiOflpqy1JbyCWvaNd+gayg7+6ZbC/dCmZPYpz0
Sg55UtpV7ww3m/j/DTi7SpR72zqbokBeMflLxL69B//Nd9nLStiGaZF5D7T5XDoMI/twqE7G54i3
T011/5iwnCem4AY5ZcyqHwbNcx/LYGTNTZ2AQ1OIKLTkxsASDb86I+x8/1dsc7YMwXS+vxPExmP4
iaoEWr5zvqb/lII2Gl0DbJwMFWoh8GLOT8AuhmykSm2Kkg4ujjMMphdXqCc5Z6aQtNW4LG9AKVkZ
+ynr0tqqdorBrpkoDBTalJFf8p4jf9d+tWoTxNhnqlLTg6fP/8QFxl8lLDHU5aWa8U0gFD6IUWMT
PSszr1yewJS75bgAJaQdvW7C76oBtVJkDZlxtl36u12XNfhIYxU3H1V/Rj1vHrMRQrjlPCCxmi2W
dXBK/riVmCv41RWZ3+PrVYLqhcIEvsXBgQKHiakCf2Jl/oXsanmWfMLqvJXWD3p7/wCl7sGnBzFi
HNLlkVRcqR0geRw2LV5OZbfB/movHzSArweT1cEh7y31uPd4ME+FewZ1/zaLI8C9zecocBvkhf31
oAEgkWdAOwt6Z45rUHemnF+0ekktwxaktC9+efo/2+Y2Xv/eMDA92lLbjJolBRUh54c3ec+eJat1
HWcFRBvd25sxrHOhNaX9bEuZ/rukv5HLS8WjTxcDinYEFr1d28PnYW24NFm1a1a4IkWtm/XyEDPG
SnubEGH+cjev0ZIs8AWIu8BPwIFCPy2geG5z+hD+EBjfB2rDSGgTUmoBtZmq8w6pFD5v+D91Lgmx
nM+HSzGig5Ea8nXsASuGf9hG0QYGpn1LFt7Kk4ehwil6dM7RgkK43edkYBb4qZ6hWSvRkO8qtQZv
sAtDybKQauMHnYnSdYYOs77/FYu5jWtVIxavLQC8MisddTpr0gaj53fPI5o/r/aVGcFk3DOHZkmO
N8dqmR/AD+XoXpkf0K7NHeue2W0xlKwli1Qipa0w9sqlKF+iUZk9Ri/+S4U5o6uM692FaKYJvLLf
lQmtEfYhH6JKgflYkzSbIoXCx/agCbgauucGk9H7ewRd0jjgOEk0rJQsYNum0WlqSI5LMIU2X1G6
UW56i4PKdTLVZK90FEC3cL5KPIxgqYV6lyRHrgQxthPRS+cjhxjxeLKQW21YwtpPFCFKck3MDZ+r
TnTBKAY7XD2DYUows481xQK1fmN4o/+1/gcpOZQlsa3GtMbIVMEdTqs8jdQd5YGSSqAVLYJuI2WN
m5kiyHsjZxbtj26cXNXmuk96QvDeR9rEG00BZCrBWvxNtHNljN24h77g2UAhK47vK34nlhh8B7s2
VIL0gFuMjM4ETdnpJYtpPPFL4bS6fWEvQrK6sPB+0Ovq2RTEt6Sj6PtAnoDHWQmxXclCbQ8Szszy
CFBG6GdvE8z/btmWavcHYo70abTFuf+4kTNVwpegyBEafrHADcBQrLzCK2XwhL9O/py1NFXhLiJD
6Wo5oo1pXeMUw+mHuBPONTGYqQNvHwXpL6wwa9mPevJg5IHxeWxMh9cmrWDoMK9DUa8FZaG9LSrB
1VwYMnc/mtgu2zBCcqMR5CyLJe4IAnER6JVL4CnC8dsOrRMN/V5SvnhYNDqUS7w6VzqPayNh580L
+R4qSkfwiMabvM0c6SXFqxuO3TET3hPilILMv7IRD2AzwLFCRzZkAxu6gWFSk1yvxoEjVQ/AaEn4
OaZ7etrUwE7ECNbUyHaw/FowF2pjx2jWANdhO4SNJOpPdnCuGxGQCLuKsnQPMTz2TaXZt1WrmBg3
TyXEymVOWD+nDYHYXqOyxORzn7UvTz9sttJu+C9/vkOSnvATT7sbi1mlLucqnFpmcLl2i3oS9kFG
wS+dQGDNzoyC4wQ3LsvjcqY5W2c5wIH6tpjP/kcfVOWfzpiEQn+pJTkIRUFGhht+1TlIZaThpkUL
E3RuUVvKGe9n1Wayeb1mK0eh1a6J/lKvokGv7LEyxQjRWH2B1ZJHidlWRH6e8jkNUkorTmzizYLl
XZhSADgErbTUUzbebWjYXnQc3lCvnsRqTG/RnSLJZyUEU2i+MD7qTZm8VWraHJ+GnA5hierouYkl
KQPgIIr+/Ea/kxXjluh8pSgV1p6LwoIyKCPfdYnvs9+rGxTuT/wNe9uIOem7LHgPsiw10UA0x2Gt
tCbfR3XDbXg1+A1Rl6jmTFuu4pOSZ63JrZPaqKhBoeLWcySgknsIvTWCooYGrT1DUztAKrmaSlST
tWZP8HCByYuMFyQSTvXZxYJqTd5EE1Y81hOQVjuEePk3YcTfccjl2q6Py1/z3XbLHtpvt9UuviJW
tYOW5AbiSvwTayaj1uvhgzASHcoPFmbOvQL92bnOJed+iLu6MrNXWsa3slTMLZ2VYSVU9nRtTlz5
PkWk0/+jouc2lPj2Kg0Yq2zZ62KVji0MHFu2fwLRMYzCLV52pg8lj9FrnOoiYFDkllszqtIHagFc
vtyt8E90CYnRV7OWNIAABfDRw7UXLwM5xD8e29ZtRc9Nwd+4MLkJBT9mOKIbpSxmLgbrLvb+996a
obZDPtN364Sk9TazVHGslezsE3bWxQ3hs+N6Bj77ymx41rxJXoIGWqHEnzqUDIp14pQd2iAtvmFg
IrmGD1ySY4M/RuBRFEvfdQC4ewMKLk/8ohaXK6RnZeopdMoIWN6iwOe6Q8wwsozPnbjQXd2L9SNQ
8BCrdtKCRMa/AZv80nKpcepB4rCX2ddmQ+A8T5pytfIteL1Nwjgh6R6bYG7QMIHI4wk+vbQ//r9O
EH/OqfeQ/4MmDx6BEh6k9oinEmoE/mBH6jOhuNuyQk9PE/XnuOyagfRYKlWul7Sk6OLW76wPHyDb
hH9zcCKa044BweaMxY8tasNn3kAgm2REDf++UVorZVy7jE/mHZRTAIy2ViLH6BP8kpMmk/kvtxAi
nk5+qIo+rM9lRpTYBJo8GaeNLg1BKoxFseD7jhtSUEB7OIABP0RJRJJNhuvhm+46csfV6sDBI7Km
Dt4pYQJHoEuoYbZ++Pa0KMbXXu0IK27pnF/iYDr+hAYBMCj17A/Nzat0k+LsaNwRK5/fiQxm48RY
LUl0K0XAl366xYRdYQRRcli8pQLv6n4oYm6Z/PF1rBmUmmMyR5hS6hkxgv7/AKtWjAzWp5lPBDJY
7BNFbvJdUybz7HutABgLJ7fc5TD23xYX5jU1pmsRXFzOx4o4Ta/GcWmolql4MZ2uq34q/AJx8393
nbSugXbvo/JxtFc6envLleGY7VeuWo9m324kmXWjDIAvfqOUeB0UTjKDiG/H5WKIjytZLy/Rc45y
k8P0IKkIQEq6FXQYl/K4aPQxKJGT6/9AUjBi+7EnED+sG5GkHU6zaExEIQLhhOYo5ueEbq/lZBHz
qUpeJJT7JXHCKCj8NGtD8soDJa6NMW/b8qrxL+vdHJGpE7sZUZjo831GUH5SRveJF58hquflv3oq
fAe+yIVtkTA9fYAi1brIp9VLCIf32LK5hsDbHzwvM7Bj0ahuctexEkeYHJe7AP/z/21sETn3NOon
3TRBlchOEauQQh5Ox6KnG0Loag19EkMfpKU1ojNl1pIekcNgo29pl83LeMls4DGviZhJueb0EysW
zM44dhraUGwfbAraE6IutRJTkFrvyYcbyaYZmaXOQA6YJsvoHuXxnYKMlsd2nF0lxTitcC/1FIEE
PkxK8R43bAi0cdEczzVfLVr7QUAh39LcJontHIOQ0DNZYObKZa9foztLPvTCsrT6ds14riW/ISgB
lgLblEgB7bYBpRRa0OINNOGs+dcNFXZJDxfguaHVl/M+NhAY1L1mV9zgBWjIUj1702ZXWBAymS82
XptWFILDt+yK5x4YEVHKNW6cXUEsGA6lzRU0zEG+YfPrdua9LfHPBP55i8R3FlZKlnUwu+4FtL1M
/Jszcon365gKp4F+6RWRZgvziRs4RtOit2PO+WMi31bJTLSmb/LOVY2WBKbaVw10RBUPNlfVz8cT
0Q/ynr2cw/DXAOtgbaEEuCctapsgn1x2rzi37I5oq6+zeox8wuTzmpKIZUYPY/JTAwunfTok4Clu
Ou9gt4mt9P9pHc/BiKT/E1fDeI+UHEi0gvNWMv626pax2+O3Dq6SdOBdrMUrcAo038n/cWaLA2vX
QVmAUEGaVR9WUG/pGKUkeQGfbnSIcTt5KufzAEhNFpFHGBMPjcj2kZ+evla0WAmMgCGuvoHIlnyx
5tj9VmHbCPFLU6jOThosyt6PQT8IrGvOWqnFs7vLZM4ZWFGVAwUSeI9HNM3S2lFNIckrxBEtGZAc
+3Nz6gBWOrXLNgPUE4z3SS/q2wazaiAxeG6XK7VYbFoRMmDcluPDuVR/rM5lxR8dJcOk2fnklDXr
Xyl4WoPWdtZVJzDRgbej7LlQ8chjACeTzwaSU2/H+8E31VZDVFK9XjtCOT3e4rzdEGzUx9gM0GtB
C8LA4lUsh+Ev/7Q/9ZJV/bGUrOp1EiWUUROe+AtrAax3AUBAuBoOJvHKpLX0xBENUv868EO95PCn
OPL8zmh3Q/B1zzL3CKprTf+nRmBGb7rlXVDGN2hl8GyKcV2ehUmY6V7YIZQei75b8Kl3Kfxp3boC
UlTL4/3PJEcsxpSga7+GWtMlpCBE69vTVMcBJ/Ha9xqAaEcN4b4PB0WtiSwhL7Q0FeO6rDTZ6PWN
Sm5jKFqFHGiwreVOWM5DE0C9/zJxmpJYEtcQMUUYeZAmW5jChlsa3CPUemBTq9+evlsIjtTvx+Vd
9df8TVxMfTKaG0sblIpazbRJmpLFZ+EHUwYdiYBuVebakiZk/PDev042tXtmCnkqfDt3+L4u9fE3
hIluK74P2XVOrEOm6GwxX7v4pf50ExWdXvgFML0ySXJQJ3z6DJWnaTZSRuY7A/KFAWkvLRHIZdsy
QTbvqPtvXDMpu4PwOUpeM3IwDykvCvkacOwOZuJktAv59e4LSasNoQ+lZKvMcldBVWn6/3YrctME
N06IO4kKJXnGmzwxc4bpkoBXBR3nchUAcxio+CWdOy/cwobI5wgi/QOkvpkHBeLqYXWlu82Nj0zk
Ou48J5o/e+rmHkGzXaXeLe0VFWZGc5WW9Ms3GqKOdLVn/2JGwVVA7bbcu0Vo7g6kP+6wTZGtuV0T
ZYD09DX/gCZn59+/VZCvrxLi3YOl//ifUDPVAOLLCRaVFIp+pqnhbQc+fXGBKZK9tgZ3ItkV6f0g
g7XrEqRw4zviwuQGlDqPS8e0viXP/kJKywTZ+ME7Z1GZNv0YRxhye4W36qiDn1cTskxH9wQgcl+d
DtaRmq5b2Y58w0SYPH7r4W3uO8fXCRHemF5ZuR5VMTru2SB0mOceQry6zkPlskSMfHIYAmTBvrYP
GCN0BVCPYnqxm/0Q8p3hh51ywpQQkzWQuVfieK2ZcTTL3U9jbAWFyWFbpEJ4SG2gGOo/RVASSM2N
RRzsQwIHNZUFFn7rzvIEnhCp0g0ujfV7LJPzipWtco+XoxUEE2/uDJTZv/D+FfXeYK84CF8cC5rV
5VAxhDzIXMT5dZpnkDs31Bn1GnqJSSaWLa1oQf1EG628jHi6IsSLO4KFFXkrSiMeKNBgueaxphTU
SCFu62qWgETBcq/k3vSelv2Uwk/IdzYFEgQ+tiASflSNUXZsCu4YWk5kCA1gp0OK2PgqgqzTX69q
oz+j79YeYyqXifDRkKL+3seQahLQ+YCqXqSM5/K+WuePEQVduJ+JwZyPEE82Xd+jzkdMih0PAxSv
qlY1RVY8sypxntzqTp+X2ZFmGVGqz1PsaHJspZiFCH2g3cd6eMqjfkG32NjA/8KvlnvaAioZHE6r
sH1kZI5S5bjkKurxxz/DU2ZcgwgIdRLSbSGwsFOxe4ijMiIUSOPp8z9cKfE7ZmpB+1LgJrRr4mxY
rHC/7L/eNCkyOw4luYSZ3silDVdWTPBHYJMAYjWoUax+PEjcrp3nMF13clt0+fXf82rijYXLMp8J
YZWaflMYWw6U04I7XVejncSuJBExfSCuBMX4VmOg1qgazYUquVDvn+pJuFO4CJgnswuYFOXWvHDI
hf6fdQZXlDQALyw8oIIUjzsXHoiUCswDNO24a8+awi8Z11Z/NEETEe7TVJ+72T3ImIFvJWvum6aA
eS5Yr1aNBMjg5PEo6lk1tqDahv2jxau4kyd+FWhXb6oEoxAbhBYPce8le59OQyIsYkDNAGUAk8+Q
aiE7FpbFc6hVpIn2cptdCGG5JYYsHLhVce19MjbNaeNRc0gDkSVtQFncBpr72tbJALFu5NSO6yDA
eEA60fwMyKy2noL6mkCGFFiorVSd67BM8BE3coxearCWyyTBsPZ3rp5liy9zlbIJ1W+QEJcwoIuF
yP3uxqS1+WNPPUJBIzU0Do0y9ku8O91l/KHwmdiMLS/LO4+Yw7w2PIslVAr/1iZRv/kuQXU+fFto
MUw6oKj1thRQT1SpI7AinDQxa3kumvUud/TlB8K42XUZA1Ifrq1nnFuw0O475TI2vle9/3TmG9BC
UulSW0rWIFTMyGiB0nhRvyHIqCfhJCqkK131JLaFXYgrBNY3RDUsS/zeflwHCW7Gp39JbqZiujxr
+9mU5Q/GZ2doqcgXu/M8wr3DjQVo8Q/ESOFoE0FYq5XhcIFupuyzH7bxS/GIibTKaUJgs7vAc5tQ
tQZqchdfQYhmUkvdk5g/kyY+Ur6Zk48bo4seYQd2rueexKF3K3T/VFl/ClQsuIUb4/rfmjxhnxlW
innTni/YvwIi2onAaln7/U4EhioGX/Mb4R6C7Ob8M3kxC00z/RirmNYQ90qXRXhBKana9CLzBDWE
aDmBl4vK9I1Sn7YkqzCBjDnTHkvAD/yACU1C6/+5tUwaOVUSNiVBHNpGg30LCEXCLwoYniQfM0hy
grhaOgIEc2q18WnNszVDjmkczyEDoYP9pBp3JpScbAHEfwHrB+jDJsrx69vdczFTmQSo4s2pHwNe
4XBJk2ctknE6xIzypSxxBpU/mcySpHGAdlQXWYpYIuKsmCLLv6e45BvTwFz0Gn+r1aqImEr5yLma
Mpcb7gMUwwxPQofOch3XHqZvGUtRL0dm9uNJvLnEWBtImKVyoc/DtnwrEAqs++SMHDopaWIv4kOQ
3bJGBu34FIktzNJsQ5kMhqt/O9A7e20NBNGaysalgDv2meO29JA2mTXjiJ36ZFic2OkIYLtMapYb
kQvbwP1ecTCD5+VMjzgwhQwqZq39ZzKhLQSu0ipHIK9v279Q85S0m2hZQPojgaIy0kG0pH4hg8zG
S620BqsLvCGosROT+TnsK/1rluVHHLC6SqjBpQgRmolQwwB9fcjSFBSj4YtTsbLoT35vvIgWquZ2
AKRfGmf4yFx9QdLiUMXO10RsPyry+o25saAuX0EX3a2MN6xJD3ZWEzyDiZXZ1B/CvUIJ6/E1ru5O
kO1Y349S5x6BpDqZ9Fifb5JII4JhAbCieRbgxccH9AO+WS93fiat8ybvvdHOCyXphdNQg4KeEJU4
I3jktLLtysxM0WULd/jaKQXDCYt3dsX6PKQkwnvkj+IKhE3am+/CuQ0KFvsbLv6bHpQ5APETUfRz
MUTiSpsz2Xvkn6udqiWfurrKOJaFtUZU39Ay8mp4Lcofu3TLWpWQBoQAiAUQB0Bxd+uobMe4W6F+
YQlc2u5rJwPiv9E1xlYhZZKze1gS86PQpi6qxZGSoRsHjOZIVGaZDRLbPfTh5cuB8/DaA9i7bVOJ
N+DvSBC/lv8agBaeKHMAhII4MK3RKXEQ2WivQg9GnbBB6/IbVky7vI2lY6F8lr0sKNSev+I3DrDu
hS6UdJBeIt876BD9rjmKsHEONYbeu3ou94qwtMlylmIh2OA7ekRR7F43dKkkYNY3pg4TTSINnNGd
7tFs5Ivo1nR5S+lvVXPxA1kuXVJ2ZZFu/hil0BeWLQ5wL22t/5MkmYooCc+qDCqkmKwyRFj6fiee
gb2EUovCW15WdNBeiq+YIERj9Z8ESeWn84qQzd4TXqybCmk//FfUNk72ZWMSt0uA3xRUA6GaqlFy
8g7rUDh/5yDNGCnmAFQ4xoooLEfo5tjdtmfw58zBP7PL92ptgAlknmjCe/qjq2K+Ibu9x7UFMdhL
Nvu90760QiZ62HMJkkKgmlH6bcAueHClUSqJfruiuhWm5ItfGN0UAVDQNjpDgcydNHkEPKA3PXZL
lCD7PF9Th+lcHj/eqkS6QkJhdPna9YN1QaEfrVY26BZUn3UMioGqzinSNISI3Vmx24e+Gj0/q4pz
duG0uXHLqlDr2YdujylGkTQOQakJjKhdypuoGIzv3pQDyCmp0LI1/k/oa8st9zNL+DM6zrBKdY36
3ei/ype8H24X5UjaGutcck2V8Ju2MfsOI9lrCmU08R8QxKyY2tlMXe6BJ+SboXcn8zuRUQklZ4/s
3v62T0tF/8i85KIVokyUCBMVA87h3AicdFKIRuSSS8szJpT3iJUNhGMOfK4W9sQDVOKRk6jHQvE/
is5l844mX+3MjIX2sXPlKP51NG0tJFymthKuvF6ad/P9fXUQWZkdanH+YsAaKaH02/1IZ8yGTd3J
KbVQefr5BNMmv/wTzvTvRvG5TevkWqRSRD090yfGo8bsd5Fjq0ENCImMG8rjBXR3R2Ft01iGRE/t
Jops6U7iSLbqOVBE2eFFR/xd3pRV0tHKRZZKWcQK2il8G0AbdnSR7QI7gBsP2SDShpEHa0YvPM3O
y7X0TR2LXvlx5AhbLelap5AwYY453fMTw9Tfj650PqUaCuOTcsF/MrVAERd/gwJPrTIomaE9F7Zz
qEzoZAjAxCJKLWJe34jkNgHR7lDoh7/bxLMdw4jqImyQuwqnAZNd7+Wnek8dIrlBX8azzRGoC3mg
KJZqIZ2TGID5b7cjVyYfmJ994KFA+tuP/mTMlNETFinE/v5ymj5l9YCYx7kKK3A8hQtS/YZff//8
qwUvPr9L2OWvqZLGjAHoT6sp28WdNDJZU/BzejG2tbIaizURydnc14lzaGRD5IyJr9nbjudt1mhE
mKi3FNwhsEYsj62lGTSQqU3y7prre8BScHE5yM94v98w0hKiRoF8Qxx19v+BQuOQPt+OwM/A7jeT
ep3qWTkfv+h4iDeJengsykJY6vtiPOYzrHOxf30rz9ScBAXabl/XGuCa/tJKEnAyrYlh9eI7p64x
3l6Db5cVHGQ+/luR3nrs+bHfV3MyYSYzBl5DNYtIr/DLyQ5PMDyOmt4N+3V9OAoT+Ya6iMFU/k+b
ekvKEHscg+DnBx5GR+9uJdJ62f39rlunHyjfp7wkI1M4oGb+/qr1EK/OwxtVENAbdLxeC4ZhlsoU
tytT0ApIxXPCuQ81YfkJBGz/YBlAAVE4T7SJI1GRVqnEhX1rustynEcD617uy8WL49rmFQljKIbZ
YOzlPuGj4Jm+x2oHLG6e78emLosLT6s3boypwIR4w/jHusv8UKsPU7ciVcxg265Lg+DZApdkXl2v
t4WRQIJmyZdTFF5WfDgMS51UxmfdNYPopsOdw0Pp4bWGxEYx+DNJtzT3AcXzsE4LhC5YNFT9y/aw
Ew79nUGW42rsBzSzrZffCWoLIyXCkSqs5ZvMAeBkz3Yw3HtIYcCL8f2xO5robYHFjg3HOax0C3kJ
cwRv4cDZVG6KIt/Jc6vSzRUD0ah3QbmXxKmqwGjCE1OSDgsyI0HVEBKXAfSCJiGD4scnvObwiD5g
RmsCh6kQfe9OwiySbIoc3xVyLpFz57F5rnJxwahuiVzOdS2/Oqz8CNsfOPMF0lmo02yfJTmH6csy
PLSpr4LSBvPaxXdgqadl4BARQCNAn8BzOoEsXcmJePYwCXm6gNp8NdX4tn1uZbTutxOZnHoxGV9j
UXtAmlPvT6gj+QehuhWaWF4ate9ljGaEZEXVuNWVoss4s6w4iiuzLH0Lv5ZJtoYN4OA9/wKA6ejb
lURc6tScYdWxjPODrFplQzcdY6WZnhqEbGJfEwnCET1yT/NKEYU9oLaGFjGzuHCjHm7utQ2nvELv
A0zn2X5374aBET4sLknAScaajmEREwow0ILi5dAdgOgFUqC4oP0jhtm2vUtMeAXP3Obiv471w9yI
wwrtTu+aX6XlddY4Mis4n0sDIfhG1T1Tg+ElVd5nAVlu/hvM8JoJIAb3gCwZYQ+jp+6zZHLT/wFD
vTvnkKz/XNmCS/F0m438TzgQgB9prJWsMZbHOn3S9tTwppzL4CzLP7WCqysTLa5MNNQBcHZK0g3h
lhNJwyBVyw6jf17aQsqweOTjAV8JtLXXiuR5FzJqnnWCVI4Z8gLXcrEgKIfPBu3XSopL3FVsmUDT
1HqjwNmbx8N2Yh4I3Scy04W4NTCW8yFr/+DLkVGfs58KgAXcMhpIQKg5FYfH4OVFEf11TdnFPR3v
bYiFC1wcmJ6aG8U4DGhlHxu/FbSxsCv9ijKUQIpv6xzTkx3ZdSfX8JeBJLj15597NRYaDaZAmFnF
g6T/Q85cP3uU/pPcMh3d/p0dEmCxFc6knxU6YbX+7Qgnrov8ybvHytqObrZBCcN/fmghbyJONpJe
GZwGi4TWuMvpOzyAm5pKIJ+eMdgNGhUzx6+610czyyWx+/8na4a08oBY9gSmrqNt2K59Qq1XrkB5
h8m3D8WIzRwoBcJMRywHepspIFsJKlxuGHVTsRMKvnWeeRG2SSi8OzcgWX0KJBNGok4oH7MpLnhl
up/cN9CtxfcYqV5jU2ydL9UsKlwtTzqQf/ACrWXsQOnIr1FpeuoY83Pzk5htJvtfUvjPDc0oeuLN
GIChbUNI0OB9XWkO700AOHS1XEpsUd8AxqaORVgWK2PPYuwnKnaHdil7e8joK7UKxxL45E6a53N0
5c+CGNWEyAarve3EMSZUFx+A9uFtOnnNfD0xSV29eTPYV4wOhbkPeYTRzi6m3E4hFG6bdnN648BQ
XwER9uMuP2DleX0jvhSKOIuYbb2KwWB44rSWWN5D7evZYppwexc45Q8BuMaxDMXtPG1iVtFFMG7r
fh6NXW9T37d2Tq5LVR7m9/Qfsni43GRFGJbnTUfEfPmlGfdXXS87mKhA/6KNJyoatFg44JnyTKTI
UPhrx61h54VqPiHPv0hteuMTbHzF2X9JxxZ4fgaUef8f4kGcu40iP8NnLqWGp0nOAgAVcnXMUJ2I
Zx/ZrN81nXzEF4WM0g1oYWKP4VS8phDgI3wMBuE7N6+kLtDlmHsmXErWTwsEyaDFbVeHKXo/qXMe
m2/z85dql4ZyKM2roo79zcChXyHaH1UEMYnCFxYEz97/i+IyyxdkJp1Dlu45XEYZg3y4Q299ALUb
f4vYKZrGQXI+YsG2Q4dFdbZ1evi5YzVjjvMM2Xn0NAaOLiAWlUcJLBJkV788I8UHf/0MeAS3KzbD
IS2VwUufYyaSCLBTfV3Hoj7+EkWxM+r9QPa7VmwgKQOIV7YnE2pM2YDb1JDwa33jXg92bCARdWpw
4n4edOnG7xgN82kV8iVkzUfN0HKV+z2h/lnCvhgbUA15dRoK8uynD5driSN5TH77UcJr32dlFc2q
uQhi97cCPbZqli1WFyVJ1G0SgRxsi2ScivXaFJwKAzgVpLY2KyNcime8DUrQGq5ltp83q3jrlc2v
9lbVC1UV1CnXP/gn0A0k61cN/yAPpLrL9tNoviJSpFO5DfgpRIpjpVqvSaKrzuK5FxtJ43HIc6xp
jPlPxB5njOSWu8Ki698xUOlGvugC1illB8UybuSw7DB0rSpPFyq+ab5YFaMeTlzxzHH/qIznc8DF
0OX9djTtC1slWdHWbhOnHMa6jYVmVfUqjaZqt6Hvfn2jXsa6dcRKNeZTjHOO+Rkv8vHknnkuuH5m
KwCRVRMj1B+nGqwXFM4fWtmohqMueF+ELNQZPplwOrhMYoYlQgWug1ZlY8p2PtdXL/9f7BVTH+Id
Z7Fn0DF7IQikTcYnnZyq5PdQ4zedC4cXy7XUm5eX2fTfKVayBggPL3lsNNVXabl8Bq9VesG1DYyZ
WizIXRaNACQQQ+o1b5cyEotDKiab1skaGpcaGqN3BLBnla0FfZEpMD6Wj4LD+JWNUIMpT/3U79zZ
IWh/2ML8c4FINZmv8IEo9Y4/QdHQWyi4Cuxc24igFNDUu9yvW5qkH/Kw9TgD2WafHPlWCTAoU+tS
SPX1Nf8XYS8naLVcx3PyD1h+FXuRXk2l7Yj5L5X7Fmoq4ltbtQdp99w0aYU9TAMsWbPk1C15rAEZ
5YpsvTgbYysrykcYDsc2G3+Y6D18OUWfPJn9K8uFpHQ5gkDNeLxytkc62yMEf+p1tbQurmzV+7RX
dvL0UMBfUVOIbdkQ2UAAfGemSsjH5UxIb3mhtdpR44yI2n0OnkDxzj+2o8ctvJU6+4xgZj5ShR/i
CJ4XN/qhtqd9EBfsiqccs9dlrWLqpL0vdTsQ9gliAstL1S48BZVJI/Dlxt8YT2Uz/Z4ihH0738+D
pM29e7ghloE6ChZijEk8yuvI1M22FqanGQmJsY1WimGL2uT3MWFAA1FLZg6jgeO/IPG4otzllJs7
VmvRHiz3F8lxz3ywSOoKr6XdYeaEQzoFumxr6Tj81UxQjJhamD5dnJ0ULcIVmmPFA2nnVyBKg5LG
9viy3AH0K3Q8GEvMzmOm2lS1ZV2ZQ+waw9mOSq1JlM0fRAaLR6LgYMwTaEKqecLDPZISJzWpq2Z1
wGlKZ6/nmt0vG3am1+pGRJgKepdqK1aZ5qr7XRsV6JHNlE716CmhkzTRiDDgqx5UBGN41fewV5//
YUej0zo/7SIXK9Yp6QNzf4vHdSzyKBgawU78CCnJ+sBEvoOH/8Ymfep3ATBgaD0XcH+6fb3uViHk
gSG9y4wRI7BhBaLNn+z2H21hTxpJvce6+gxoyXF0hxQIBomKln/GoJJKwqCaikI8iq0rFUKb2quv
zj8QKmFXHmW4cRlM4gUYuIHYF+ih0WUHVr1cWOGtqjjMCWD08z0VSxgOGG+55kK6hk048+KJo0gc
QvZOGM8bwqthZn/gSXZzGoLG3gDl3nvjzgUIWmlxiOY0aagJoYG+BYrjEKtM9cHnLghpLdzJEDLy
dkhkqRIRttgy2K0ERbA7VRjSGAjGJJb4xGft5R4mQfaUI+TRa9jVdGhfOtoJrNwtbXSro4MfSz1f
MGiVrstn2s/fKMlgTJQ6YcwbkR/Cu0OSRV4B+u/Bcue2XdmBJetmVhvuGuIemvxMMsmqCaYjaf1l
7uWG4am8+uEJvshCxgKlnTTWT6cC0jXgqmPJA3VUYg7xq6w9/g3MVooKS68cdbw987rFXEs/v9P6
UFfEmtmEqAViIAayk8cpds9oKmpDXVB7bv0pxv2Ppmu9rq9Hza8KtxdeD1V1u3d2gMxrToLzf4Q5
fDSiJwmr5kHWppX/NEyq5qPti8NAhBTPnhcszo/OTlYLOl/wpGdy4qmilYOb3ylCH1vrzddyT0BH
a5TUQkgtLysmexs7ynXIrcI+as9G01RN6CU3L0fLp/48FKA1tolcqdksFXANWtYw6Bi9QzDl8B/t
SOZmcOaFUbvnvbGGi0lyb8qEllwzz8Gulc6ynMVp/gdXOkoW++fM+PdnVpiBVb3Hn0EWtwS1VkMc
ZYo24IcZhL2z55g34EZdIoZoutELXTENEx0877CcIHskPZmKA+S8w7y6yrGrHM+RbEwcxgGmI6EK
Weekj2GaQC8RaluDhyfoFer9SkFHXaia++Rq+sv9rjZ6DBoGWclH5b0N5b2ykFdwyV5JADUPlQ0h
1/+XUo7joAx8KZk4su/4PIFX607uvLZBMrk3YASnEXTtveyjOzLc0yJHUy6tDi5/RjOkk/OSHE2n
tdXsALXnoyYvJ3Q/CIm0SdTgQKNt1MDpwUBkbBIlQS2OyS99uSwwovGmA9NOpqpa7J0X5jfOUePJ
WndC1LV7ry+F9FpJNcW8NRKBA/NamrsilHSvzmsGWa28nVUyhUupyLaNQY0gDSH2rIp97gjoMt+z
Ji5kWdZUkkUsUOyp7V++LY/TDxAe9ZESvkFnFR4CsZLA7J0MFPK4l0SIVcw2J9tlBPIihYct9AVt
bz9uyykcA+Zn+EA2XvAgGmtrWKdHDS7hFLFlFAiGFGZBQa2Rgat62MxbqswFILBFf5nJZ7yt+51v
LtFnp+adEBaTlrYiSsz5NUGM9PNnCrDl+q+Z+JvQPMdA8bAW2jru6SxLGXH/ZKX+00s8QI+D/bO5
BIExFbIQPjkJtSCHO8FsAxpOEUTNDMJaouGSiRFPPESe9PkA7ONPhOtkzp187GKnA78QYwyE1oul
y5WgeiJ4BJFj/1nkBeOK0EVZfuZAqqZQ+Xn+c3R0tZMPCW4fsM9T/Tt+pppv7yCvvCdrOMPO6ZKo
FZnjkgwFjwYQ2RRIAKahOy1xTryDRWAhKgVALdHQOdc80UV+eXH4HRT3sUGgxziUK792GxYfHwrr
IctEpKXBxmpqQNKkI9sqeyBKGbmr/mYalYd9PGyfhMVcfu023DdTsMrhp+XGsz3s9fR0QeyvEnGV
l7NTtBKdN6rz1IktcJZUFaJvPVfD7viRZ6XWl3gxFTBs8w0uc9orxfjC1mQWQn3Y1EIx5FgrXZpe
gDxxJ6ExXN/7S41ZhYxE6nQC27a/OI60xsx495BzeAZf/LukxfmebWvXj90o1aCn5TnUUuqrU9AQ
skS82n69Fku+geiqPkpr9Cza349VlWyzbebO171lOD4qPk2A7BktD/8NE/EY0Jvd0xYUB8fq5pwV
eOdVCurQBL/cxmyDJ3oE0Ls6EERvVnDLt9BZZUPPsXOiNdoCZ8bj4vdoW0zA5EAyoOiz6HEjAbnF
eQ/0gSk9Z8lUR9dhlJq3gP7p75nRQm5K/LH6ws6oFvuHxBulwEUtdoibmueglxO8qQygmC4cRj5r
8wRj56/fLDHQ+Wxmq4/aWt8jDopAr5Df6bF6B4zyzeVJGfc0S1hShpPg+NkSboyMM36IkV9ZYoMv
q1fatIqXIWry+YuxocG9OkZjT4YwruaOXv0O0RByDCkdaNhGWGVyahujZZWAXMRlNVnw9yhHboMz
0W3CGSDkTQ+3TzuSkI6XmlcJGVqHKWCNF7Qj6wD3MJ1uyMcFvGXCdYkUiNiljCBhX/4M6rSusOIj
tgxDpGLM6pUw2LTyMXYB6GXqUn+J8LgmnHxwAXsgstk8Wvf291j9hfsv+GPaFKp9dnOhtBb5VfMS
TIEIYZPMfzUMi5fvD3ZeM3XXBPtehLQaYJKK9Zo7tPP2L+oxMmzoLzORHvKiw/cdF/6++/gN4DAv
H0R/Dja3TzkD78PdSP58b9b/fxgkBD/yzNiwi1+QkH0UWmM4DAzml7xoLkzau9PT3djgYMcq/V6H
QtYGcsTk7+5O0isSI9IG9riIfu4nixJ7HJzjJ7Uh3X5h9NjpnEQFwVu7Wtx2OtAkCOkihVjmzQGR
FlPpmRwILuWih6eWR2KUItMB3I2x7BDo+WPb9msoqXN3ilJWYlULE8ZgyY5OGrx4gMZ8HC39/JYm
mDcZCDzf3pT9qTF6fgmIIYCaq04yuRCbsibPIPJHC3yoi+GHTSGaY0kdE9sQjyUHBooxo3wbO10g
/bc1DHXCjS2gjnDc1DdftPp9OPSdPTGedJfuFZnz4ebZOfgtBjR1VsbLBwMqzfJtnhqwPG69Z9hE
aaURTchtwhZjDU8Ehx5XYixUUkeIbHOr8qGyEFoUVAoyq+kmHGcWE4Sora/cmbE43GWi9tFllsVT
Yf3UyGa9Wquh/LNYbtBLFfPxVkfZLQR2PFcmzeln8o0eK9FlmP3YhP9iApbgNLkYYC93aBngrMov
MmoEv3s9NHRrWjVAuuYAuUy6cMqRumbq7DcqAz56WvhdRD9OG6w107+Az6Fplkaoa3/a3qGvKYi+
qRLoBHSo9kM7cMETKLrNstAfFxLZLgZFRY/njYdmT4c0S6XqC2hALa4VEZRLt/L4fje1FgQRjjQd
tTiOlWN+C7pE6ypxAhskc2KdzPQMTYrCzFJ9qdjkqIZ1VnHsFs3+ZZmwJWVZHOlyNpqtTAZkpwI1
9tjf4J27GP8FQnSG2qaW/tpAgNx53QkMvhqftcBaYUfAmnlQlOmKdcdZDZ8Z0pnBDvF3CW7uH5rS
y7+7OqUKf9HdG9Pg1OWBu4M1t4biVWzQy8ZP7TWtO8p8bnj+5soAz9xspFj3+uYaLlOBH4wEhK4A
5eM3P5c6jb7M40zWOFu5ezQSIdRJvPTt957XvOGjJkm/Gc+TEIeZM0fHPq66nr546PN+DJVIeD/9
gM11DGecIOaS0wL5A1rmit+k7yB53q9vsqawWGJKUuBzrYCeS1ufIYb/JMSWH1zp5LfyOfHmkzKG
j8eG54UqM69xu7KAq7eDXNUgv8yvsLOot0QXQLWNlETrULTEl/EJg/paqXS6QAE3INqGiil0de+W
GRYyoblbrgeQJhEEzGkOPrm5h8JaWpVF50Z31A4dNe83Chr5/axeH/wwjA55xR/U2C0s0oF9y2RQ
6WyUrfmflSCC2FLA+hUF1j6ZUfcDmZ3+TTSREr2cD6Zzp1Nuh567SNml79rn9sG7zdqV7ZQnjti4
vnP1q6KVHyFJfJdRaWyA1Yt1IVsy5pNSJgaysI/oD2rGZzGeglLi5oNX5qQ67RBkNYhNeexvptP1
wKHrBisZBWpsvCXWoU47pis9VrLGxl4e8bgP7sSFPlsnpCKbERRZB6eklB2TkRSWpQ51azd/9ABq
/PUVrHKMNnkAA8qXAj8+U9rT2TLOTJSO7uxVinktcRolWHQF30ze97YJEzGY9EnKoywt+MfiKQCx
XiQIxWtqQQLuiXflZuaYRLyVxMFFWPmoy+oGM/An6iSPzTVhitrgyksZt7szBf4HM7gzGxzuAUUK
EJJs7iTckGo0Ux2j5BgqHhnLY8XPdXgIxnL6naFbJVSvrJul0rKaUeANrYFRqydpb5VERlqDt3J0
90uATf+j3561UyclNgFCZ6h5gBp+AF+tSvWH96hSiXNkw1I7AvXevumKNhgbaDHDHyxUiIcNiG13
8vgabt+CQMTPBKREw+2CEb3/sWnzBSYOfgFqWwBtX0g+Mf8NtHmRw3M/GtjWUpz6JfK/2d81EHY6
EAdI1tIKnSHhVjEq61LUdLnwsA/j+ONSSrSqSxnKlq18u4wAaN3GHBhBsMehojgEoae7McnKXi7r
xsWG4/vQRDXULyKMWfOl3cGinDPHgjQRrgqNZJq01MnHSikTyuZKHSdIE8oJxWHOV/1t4bCM6/4N
Gp0ZwuI8zZFZWHGaWWo0gGLH/Oki1H4PYiWGdWNGfB7gwinmxqsfGJ+3hSsx3EdRoEo0cXEysDzH
NSh6+09rSthiFAgqAe71csqUvpRy2zZ2bagymumn/mXSAxdls30pFtILA80o8jtFfPiYXbBoUD5M
z8GjSK4QS4LBJx1HrHbWfdCK7ihcRSs3oYgKpJTzljs+z7faIVWplsHUvZOqrxSh5QxiBRQzskZV
EqAFcr8aWGBbt9szWmVTWQuQo4Eyd65I9JX1fzD72RfVVEOWFWJyEqXKWzpEC3eOjtvwwPkjYMqv
QGD1T44ghN31hJZPinQXaAgSTAid0r+IaiPPuPr80aYKJdORNV8Fuh9QvPRt2f715hsXhRj9Q6pm
3qPcFI5fN5boqNOQ54WeBH0Vhq4g4YYaTyQRZoBYZp3w02g5qDqLteTVt9XkzrjcCdTD5yiMVmSI
aZD+J56p9/lh5qP035tPbNIqyLdKAiX1JNcMkpiq2/BnOe7PjrkcaibekxSDr3eyTHbiEOxvwjs+
xKCAy9p2xm5UPPrtjL35eoJ1aMJGWNQ8fN8U8Wzc4U3OzEoLdEhKqsuxdmXd4fFtk+6S40+nEYyV
CyAP1ZzBNj5XlA24xGDVlquOC1h9lwvJ8VmnYneCJvo/CTi44cGtvle4AFM/6JXiKMZ83ywYak71
PsMee+3Tb3uxiyG/r508Fzz/4nusgmyvkrblhZpXd0kqEVK5JmCCYd6BTzOrXC8U+1L5wsj8AFKi
AIHR34fFlzp5Q15jEPbW+cofGkaLHqyXRV5CoN6h2yXjurwDDryp6YgNcOUlvLdNFsr68iZLFFhz
cbcEhPole9DoYVCi4vzwTOWdpaQuDAo+51Pn0mi9XLZFeIfNalu1GF1aB3mzQcomwIpN/rZehCZd
OlwNVX//eWmel/5le/70RBT0kkjFsnRFh7FWsFuRzgP4XHe1PE09+7KwduAFCzrYLBA/G49Vc1Bq
OKGaoMdYVykMPMo0cKm8Wl8IGptU1kdpjWyUbwfoaeWkVI/YQMxNKkn1QqxIjXgOfOCDzS0sJFoy
+XyzFKAJSB95QFgEHy9KL0GRCnYE8PgyxmkymqEIwQjDv5W6K6jzJ8vszIP2Qwg+KkeypPUQVU5P
ssKfXqzc7aUiJLyw3W2ndD1+EZvVM9UMldn7LN6QaLb02PU6P+ijBjDTd92jFg/RNIl5lXP1t6fk
fv5eKjwfRH+WIz35ksekuyDyCgFnvL8UR9qrBJqV1OkYYjr/vaLfB3YlYy8rplTDNMiD6byS+o19
fxB4WDBPGe+4y65dYbZcDBO65pntaWO0jNaSoArKV1ENBrQm9RSlROSiB/vLAUGmggOBzsEH11Wr
jh41JK5jw93d05PZBgATPcnXFpB8MXJ4TWrsHu58gjllCQbzFpskkMt46s23FEQvljJCp93jSNfc
usS/Ylgy7/kMAs202Y+VBlbbxPO5EgfqcJesHftDYSge+kIP5dT9Ys7m0z3HhjKfGxvIKZKDYL7u
KjJ337BzG4rnJ7vubBEGzGdnTq0ruuT0xUHxIBoyh3b0m7yYHgYcVUSDev8s/er50BvbWfODuZgp
gfJLSC4MzrKtzqRYxlhQdLreLHSlw+hXykQp4BmX1XBPRJw/3U8T+vvnzlWHx25YtcnHxPLqYcey
1x6JaZQ+GKM04rLHH7opi8Tmm1AQsEfX5bgrbMSg+eEL/KZkh8u4tmuK0osZS7pcR5V8e0YTamOA
qTXXaGiaEaqSkoHJIoG2oPN28GqRzpWSJlx2frD3OWeXgYGWE/UNMgjeK8E5HgZ29nOvxRmg2DyM
VnZ4wBiLTLzrYt/9sD6cSG7pLGlvJfDoWaEHUg4O0LUPiQuKJfM2uPg2zucgBGQZu0TQ1xEp26uM
QEe9H3pFYGUlQVukkDGIHZXr5OWxpfUrr/lacnXGSdQeiKLuEMTAozOqjujI+KImf0AQtVpXZghI
WkvxY8DsnaWrMUwnk8EL2ck0NU3zOTx1g6Zp1lDrHCwc7toMYjoxwPJGCXGbRaQWcMq1Gjw9TNFG
PQUFsF1xm5uYMyUmSZzw4SaC50tfVMI9EVxpIIFy2BvFbhjlv7ilDILPJHQG0OhKH/2DU6P8dvzi
c5P/OpWG/NOGklrsQfE+iKgUPd3Fn8Yl4aRXyvQ0ipwNK1DveP9bbuFdWx9as6vm4SsxD99M9F5K
TCo7wA5Zla610tyMFirpKg4DVvjGF8a+7Gd+e4wuuUtYDoEYQfV40dREczxC7t0UXZxJzbWp5oHC
MegMDfvsjUHRfcOHfkAUlBJnQ9RbE9FTWU9fUX7xSd1AfBEtUDFqW2BxDZ6jpooWnLaRjuwysEJC
TkiDMcIhOeRUeUtg6uGhzyUuT2Xmvsw9qJxhZLzJiyPGFFfKLRInvHvMFvVL29prWRhtNhSMTft6
IUTvegHpTC4PGuz2HHl9HYaYQrZ+KOK1BbvxVTbd2e4QIiTjwkZSTgqzI07WDSeaoLiPcmM45PEa
GcJA7SPoy8HLrC3iV4fSKtd5WlvnsKl4gWNu86eol8OoKvVe3lpjrIuHehHafmiW7il1HdRbC2Dk
eghQhzZaXD5+qGd4FuVKLBCTR/+MecJ1/pshGFy5wX7IynSq0TBgDf1GqqIlmbN2HbSJwU4l4qRL
X6nAuasFkD4+nhXCX/9rB9iVg1kR9ZqSllsR1bzfcDLdKGOM+PthMl0YVMDlem2ssCr+ighvmBAT
+OngC3EXeRGQM8+5oH6el2vzem2A45UbtYfuK/3KUCFjoeJK2Up0Xfri53uYCct0rFSPw50pGPzf
BvPSQfFXCtG13QXuVe7KrdhGhTmxXSN2myWo0bzZS/iYjb4AoOIPvaLNZW2C2n58Pgy114+tOlpJ
XCGyR6mMRcxuMIphg2yIxCxjv5gDliXe6IXbBdJH/gn6NT2oumpSmliKmuvJ1ExFptbchu2P6ZDd
P412T6J68fuB8MM1r/FHfrExSeOIIFhJRM/EOOwJXl+q6cg8MtoxOYqvPd1Xx4N+5GUeduLXUw4q
7H1jt/nm2j/s9FRYCGq3PotMGGLi32qP+bb6TIqkyrPIL7etPUcpZHNcZeEWy/a921FVwFrQugII
wun5ZCES6WhT2gfkJL4FDn38Jmg8W7B648Ha7B9F09BMuBtqr817Mjrj/vLm9INGryGtMjKH4Pjy
0NUATzqW+INAeRWcE0pRQFv9daOlhfWRM7SQcha3vG2skDlc3tj+V2vQJJRLxc+BykpSTsE9xn0I
sSrRLpqn2T+haoCELiH6T5zqxZJAAQdWW78qXafa2Blwv7OidRWOyeEUaD7iGcu/e6+ezylsBUKX
h1vCDtf4/jp9LfTrxek8tFShWRqFg6gjqc945162AGXNAlqmmqSmaVUvzA00qCd1P2Krci5UM/sV
9PmqcAXO4KDaUAzy+gXcFv2AS4nsCgdAl18yh4LbP0wkz6m1ATpqxvIttVFUrUjy3kmX7s5/6Y4Z
FXM8ELpK5x7JrvxflS2BzjMouCVkmFnWxlTEVf0GQydbUB6DMUYekDHGLPmNNgZefL2ZYAGaBvju
FrqtO+eQVOsog4Q/g0fWPmEd4gVyc4V8Im9zKv8DthWs7+iWm910X2zkHfkAg7gSGGisn33XstOL
ZWtHBWRlNeyW04jj6kB0sqU9xnuhA4CgPzo9bKb4sT8o4ZRufBqNwbm0x6CQFCJWVrN6R0828RTH
/X9ZB6UjdPoNW30UG8Q4uYdL7S5IcBKCQr73S/6cdSHt+mMSYgt9da6wNJhmWfeGMKkxHQoPWRvL
8UKGxqoZeJIfh8FlWw3A+g32HnaNYwTSe4Xy3NJBa2vADgypxheUT7Zrs1WKgZqsXDzqjUxmROxQ
OPlUkL5/Bc/N4Y4eRFsTlpsThM+5aBJ/pEUADeRGV2Lmr9N5LBrQ07rugogCb7GpAF/KmJfoe8b+
ITxYjF8x117vU3Wbzhb7ytzdDpEB6DNeib4KPaS6fitB67e5aJpR74km9GvVZoVNXUinuf9ciuQu
CqlBk53rW4Dd6g2hJ/K9EIVpnQQhuXKxHVZZywbrz66coTTZy4xzxUX3YpJr7daUmv4QROvvYtbU
zLisj0sUIIVMzZDYFBx5jmZHw1cEZHhBxWJQQSTBLck+0ZwVGdizcCTq5zRbL7oAdL3Iml9V41XU
C8sECarD7sG8nzxJ9bmMDpmXiCpJ8QcvNQ6HAa2k+EA8Lg0d38UWv+P0hFE0VvflVR73K5zJdp4p
BT4fkkO3eDsIzVU2Pp/4oTYNmQcZmpzD97wBa2ZnbhW+7gm4qgkrkVNtXSZm7POu1NrVpm3Y7daA
uSF+rh6wUcqpxHLwNFY/EtmrXzYdT8Yybnn/jE3OEE8jhFsp4vKBattgfGmpOTBJBEgTostKsxm0
kqZXYZg3pAhE5uSfLupJbjU8B7To5Qzg1rpYpVO0FgJsmoXxSLHV63gA3iP9ee8/p0QQ83q0i6qE
MDYHJLtYTLn/WUweb31xQCNG4lg8wGEqjq/Nc5aozEJEDLU/Xsj7yw5FfR2Ei8YnOpFq9W2/9wgk
DamtYslZmN3D+L4GJdIZB3nWfMP1r15+Mm2MAaQD7TW9jX9KFvMb7oKkKNEh23tZLZ1SvsFSuROR
tJMqWv2hujqOLfgJNJTvoZIG8iBZlpvlAk2YicUQREe0DUesm4rEu6mz/bKfciGz9+yT5bNx0wCp
GM9V8M2ah3BsIEBKulQ78ItiAucii/yTrJau/wBjy9xANBJ33ruZiVWknhXFXoig/6Au7rOO6VKq
Q91khbMAMUPeP2NfuRrg4xey+77qZVswL8X8QZqJEHG0H1w/5MT7lE4ylUtDlXnsjg+bCjeEpyV3
xDvsbdIEpZ+QC4re6NC5v3KqmGPbQBJxt2P4nJmgzg0tPGjxjH8efKTyRzPU8qN2+zNfRQ1O4XjQ
3O3hh9g+BXlSA1HJWNewgHZZjpuUucFvrw6Hf9cmRN+rmxmtqtyr+VnUTFi6eGH4x2XHut+tgvqo
veMrElehfiT5eFQv+zeqmcF7ExB9D3dTzcxKrcSDPJn94LvDBOoMXv/U44Jijk98uRKFtGwY8izH
gIxghYprq42HKapYOGLmaztd02yGrT2X7JO6uJ9927AK+S8cu2WBEPTjbYSkOdHBA76bHmN9wqJp
lfsvnLKg4Jgzv0+JwqbzaTAbunpdNl0r3CTUrvDneDSaaWu5d9cC2oAl+/xd0fWQ1+yfyBJjvdfw
HlNh2ei7qAwETbzg5GdeCM+bF9410+mr+krCcOpxLruth+LcuHgItdEalw477UAB6TTQrj2CLWsa
LDUW6OB3gOVewRgWG1K4G21e1XQRALsUet/DELCo9UXrwFis+TMRgl3ewLGrULW3NbZSJC8QZR+d
VXhJrTiGdf4s5zi+LonaPNfVlTpGzhn3qRQdjX+CVjGN3wV9ZV0RkJEQfE+AP4OES++zgoTh1c9U
hAHm9GLF1Y9xLxXmP6VhngoLwuOtx2QJmF4LfMMcPvs9tH6PgjRrf/6V1YmRCHrS0PBAnesgqecz
u9hjfnKd8reEHQfunaqR4ilVPBSmWJLwwoX0cjqPgC/hieBN9w4V2AmmI86cZQNEgHRpjStC0FK7
eX2BCu2RrLoTCYixBpLae3RWT6LQbScwztzrW/YwlRQpff9erDtRh/xAVfa0G90jv9mttBGlihzc
Qy9oB7DgXzeUbw9IQ+YTnet5gJC6Xmrvi+1cxmIrMMwkuzGnmWfCeyZmpl8PVhBnrFP7amD+0//B
sJ3zuAn42+vzLqnbEUA2PI3g4QaLinFzqreujy/a7im8gKGm1xgSxB/5B+S3aMBIKRzTUtaIoqv+
u2ZmydXsAu+Q+t600h5/y58XZtce3bTFNqcuD2QkxbzvKy3IdNC263NtJ3J1hQRa15nkBAh6UWy+
bCX/CeSnTSFUAnGsjXktfDJOVzT2cwBsI8wBkQRd6p2MQ5nSlrwvGPutTOLIauJWwsFPN8cq042U
RxGgIN0pYCIYOC+OyY6an6yvRAGw4hDWcjng4eoTes5U5IqNjlNXq9fkL4pCDauj8lk7W4Nj/tAb
4p3ALUFUCaR3ALzl7V4ogwckhcj47BgDhknsuHosBWT58/Vfe47+Rc2t/wee5SqahRfQtAlt9v6b
NV+e/BO3nzH3UymH6MVCMBZuW8obVHtYXI9Cx6937CcJ6ENqSlIEsFOFdrwQyOTK7NuGQIHV/rOw
5Bah2s9NHJMA0EijezbbqwyFfWaRtmP9+pgIa4MD/Nn1KkSd6BdvZ7Gier1cbJeNbjMdEVGyaMMQ
mAslLoHhpq6fv9aEjWQrISY3aoKwmbABCIMLf1mfNnrx8AQT9XZEFTIGP2SWANfUsrk97K6FSXIN
DTh0KSXjTJzgHMCs4ayz/i03zHSIKboleHFIVamRGsouVwIe3EM1cQKOZP+GdZcdmoXF4tcCGvZz
NTKkHaEl0yxAGqt5KiNQIjo/8XOTDvpZFLinyzfAd2wRGLfVjQsvSx8akVjwHtUNJPmCcLgfCu5s
7ogJ4+56TOjHT9LJtcRNSQouHylSIkPfdTVmnLSy6dlgbeT3LpGjhxUCuVDALslhvNb35+rQc3mN
n6HRqnMdRD89m67dRyMkt2BodQ5T9nF0Nl7Zr0N/58ymd/mLKiLuc1rnRpPnXo5W3Rlf1/aJZVb4
1BAd5v5PD8OFSI+HcmSXMvpdtLI6BkjxHFtvcXr7k/g5XoHWYUqvsrISTksAhMrVeIs81GDRWHma
/a36yPdRAf/SO5XyLiCcya33ZBYLzKyIZm9V3mfKx2jDvmqpB8bT4mrgRWYqIGPvH1npIvWaNkFG
TBFNE5ddavhNxOzP6YeFx7HWfX5FA4zFumjKaim8Q5pzGV3vP0h8WBD7vqV7Fvj1zx6S9G/aPgGG
q/Esl3gJSq92Xr3duWLpnmp1AiRCMCPZbSkN0Tzf+ZNYDitN1AQjAoKZyTdJWDRR6OYoycvpSqgj
IvJYLNPv04Jm7RE/AQCMulhKd2ns9S7KxCPDyvbD5BVDArCHI7ZEKIil2rnRJ4hTRPTtqd86jvsj
ywXZi5ngDOYyLWkchLyx9W05Y4cCbxfypN/KR85qmteIKct6OK8ZgsEVKdLVeZxE26QQEZLra+c3
0Ka4u2iGQeY2srVZXN01A/jXWnWLIQE9S4AgiUhmjD+OXe9GTD47/t0eaw9MN7h2BG2J4MpZ/lZ5
T9M0ZAGBSNSadwCSptBBaRQXlFZzT1xvMZfqDfhtjTosDsm6nQUYMnXwLI3gntvifgrsbnPaajwR
jyuwL0agVvEP/FwaplUVfGjLMCjadCkClT/LClrwHNBXguJv11dcQqGKapYYGa1pzgliCtTGF1P7
fq0FaFogWS4G06xFdaQri1Id9UogC8NkIdfi5ImLMLhV210Kwxbj8uZN6xmhg5Ha0kHrvHYuHyyz
9K4qE0QCCtHonAm5i2e40HDD1vvs3xthpXux7YpCoiqQ4TUa8pouu5CM6F8FzLTYut8VGKdQUDr8
Ah491TZJUrlxRPhN+iNrcNgh5G4LQHrp/9/PMh0AopS1whwV9uub7mi/WjUJdo22CoxJx29qGDJ9
1iqVcaM7vfGosMGfKZY9jP0PXN1yW4JF6nQBXGjlW7wO+NBSAwnpXx0JGwiP+UWMn1axbyL2aKSt
/FNFfUDF/3izDiyGm7WZ8Tt2HA4qmHTvm2wG/yB55bdFyw9VW4tpLssIVt9NoxE5vujWWk2+7e39
ltmHMMFdXL0r9wEl/g29Fs58ZaD8qw9Q39ofW0EpdjyBqqDWj0urWlxVOcxn88OKLvg83UxTvDrv
fg7rRI5KEeCwyc7MMHMwuLQSFfuzuBC3D7luvks23deBv3S2PiyrcyojmA5cvpzvp4f+2My40fuv
lKn3/zYYA/NCrhjH8pBYAcuqGvpSaEggT88BdRUjDtvedQddGWC4ms5fS3gKuyUarY86WcgWpPha
+yjmR4PDnQHL0MoF2mzb7Uqnw9pNpmiummN952QtEF3Fyz8twd8w6MBIdPArKFeJxG78dFk1q2G8
YBfkz/fU4vt30gOgi0b0qkBRYny4Rwdi2Dctq6ASNHdmLJapsP1P1HdjBS81DUdlKKjFzQSUojbN
H947VVPOix7m/riyzXflRHO8Dya+j680mzr88iWSZKVBxK6zOxcdFl2qWRcX3zCUkPpEpeacdeDO
bTRp/Nu35zzfEDhGLNZzlqhC4/WRDZy/qGy75bqaTKPCO1thkygrFMH4zXdCqCIHglVDXPPBFZcm
fAYvi8aP63NCFa1KwzR7++Em06dGXL1DRiygcD39objXjGfrQpBJa+HEo8UnAHa7SkpSTsy71Obg
ycLdiq3ICSji1ih9UIRlg+3PMEzbxezFL4hUZC2DbgdhMk5W/+x9Wfwf6vILSH85qe41FSdh2ZN4
+qXUzNw12kECtViFp5KJqA5M+eW3EWs2Ppb0vzLYQUjYr1BUmQIH/hdKt9BUEYQEf0254aypJ8ZL
OIVZdYrmgIlb+vw45tS2JW2CceReQ8T13mBkDdsPHvuq7czlWnGHJaRvtpJSbh+G2FC6lDcAiUGJ
IIlh0c/kPW03sCS+tKAZl2aCHiC07wnpvPr6QAk5g3Bs6Wwl29AP+FjvmC38VQ3qfqKdAVMIoqPN
dJUHmYJWySzP9Huss8WqXrAyWRusvRz4kCKv72QaHKQGqMDUJsy6DETh0fzY2j5Q0dorkPM3NPXx
+7Zy4y39l/lrOILYtPMzCUF3E5hAJeb2NQOVgCg3kc2V6/pAWJdsZcplWh9NBm6Cqq8CXIrSs8jg
qENuXXkZAeDA2g3Vw16GiMqPDL1BJJdkSHDLPFweBJTU93Y5FqVEwXBhE4c9txEEJiD8o3mUyvet
oGHhSHHrQG4voGN6PBcauKSMD/cvLpeCEVSQqAjN6ZBskZO+bMWCJnEi7kiLIOi6tojUrQ1fuTAq
5n2FgDboPw5pBoyfC60twshRf0YeKFUOhSI/uHGb/o2GlSn9HliqgM1iiN/uFXAyYfi427H6fIj0
Oqa+QSV9lkmhPGucCrCkgGfwujEki51WjZPW39HyKlBnYatrdP/WPbCj/Td7LoaNs+UjGN88Wqrb
GeAd0a2OsRyhdSYtndGh7qfpZKWScPp152DcLIQulutVjWqXtwKIYicAxfQx6Uhd8FS8oaUnJ7cy
4AVbOKyljLWwpi+nPNKbuuuvepTU1Qnfb9uiTXxMBJ2PnVtL+jAQrT6dz4N/wXDUjzjYlrUJqOlA
cTlIwqeJPu5+yAQIK46oCWqKCCi17H2vvqkEY5imPaKJ8VaA0nBX9num0ptD9UiucBZjg532iL7T
efPL3rwyZ7OzST2lBOoeJbNdSJCLubg6W5pJA2r0jWkB7TLOfoWZC3yOmqGEHK9WNzJgHXE/esXp
ov7ILUIsSTcqTnboV/yaesNz7FUq4NbghhcbqQ43pYF7nG+etYWgBBd4xv8KhboWADTQ/OJCnAgs
BmmL8nLltfqCW7ArKn9FxMkl3EWJGHUHGK3wCSf1Fv5bWkIl6FikD/Iwn3E/0EPRwK+1tqkyJSHT
G4MRU4n3YvMSQBdNPh4GfPeENLeC5CVjh9LOlyaNdmWEWkxZpb8gA8tMfJn0gnId6ooeEXCnmyiM
zQGs5b1hpb1wu4q3vpDFhSS4RtMD2LHOh+QbWanYvRklmLRgxIa0qXefR4GLWgMiFVVhI/uid840
xxhuT5O+PbZ8y4ISf+jYJvpsLoP2iKM4Ad0PzWiHyeIkYmG6kFXL4fui2nFnhjtgQa5SZO1mAsh9
ZP0EK6ftWKyrwwcqHZ3PRpNQuB2J/lSPUpgbJjnHrni320ePpa2REgndPaMGsWp9dD4wEdnsXUDy
pdV28T9mma1AVg/m3Mr4mQGh/SPk9cd2ZFfC4VhLIfZCqXpqzUDSXBjT13TA0Qvknk3hl5BX1yOZ
H0AQyuMMQmmBXFv5PGxHrs9S75Sd1wTDFf+3DhgXHhVMhA2v9pHKYlNRViwAVv7L0dtRoFsaLaGt
YrXGlEjqIIfg5mqrTzqOh30e91KT5wEffGVQTzMHKPqcOicov2EHRKHpYMN4G/25sYuV+vWep/7Y
ugzLBFuJtqJXgT1t58PLmHlwBjDJHPFCRtPmIZBx2G2b7ClviL1J0x1+qNxlzl8ganoCEy2v6e+9
ZQgmpL24EIqCBdHpnnmhObFgCAhNFscxqjOOSP0pgWxDe89CT43KgQkvTJJvRXYI4Uct2Mbj/+EN
wciZM88Y0FUfIqfn6X+UGY/9qiT/Fqk+gYcrxilnel0LaHtBpnzM4vdfs83yR11wJk0jxkNoYnhb
ILd9qWJFA8ZEsdu93jxMcdF75FRbTBuOgQbM28AEPLi/dHRZV5jn4tkKnTopfxd0BRdO4Q29fzDE
Il+RfIHR+lbFfoYFy+wv6erJ6E0oBI/QvctcfzFljzlV2nABKS/HH5Nd3TceQ+xHPgf8GtmbC8VQ
gDlneYBw375OlNSGLO9bKjMB0oOe7PziaZqnNPy90YdqFCwQ5Rp2D3CKtL5vDejTt0jUz9AgUjeV
u/JjuG6ZXqyzc2W+K/KRgWM+yotXx04L020NNmeM2hlwNz8t+SJCvXxVb4rgKZCxTc6Q1+COC6uJ
WpQIZx2OlF5pmFzv4/C7tv7dboDtfuCW4lIVK2XRzdgElOJCbPybtlFwYKiG2bB8F9UL3HYsyIqI
7rZRhFtLv9DVsC/gka17IJ1f8sju/kIIJyRFzNAbZkE5/RS2oOQ0678/oIiRqGgh/Swej7aZZM6V
U5GKTwMG2twBSp97P/E3WaQ59VJayChPa3ZyfXe/i8a+jZJndoJmB+tAw3kP9OJOL5DeeTNnz/vS
uKibwSYEXSmZGZNyE+bjEgpwbzigOTV6BIW7Qb9UJQKaFxEp8zki3naKg6ODIkXOf/1nERdHiGVK
ef0AnFW1RnOUm/wQel2UlYRUQpwTKgYELmyjHhzklgjIPmKIK/rv16bn1LFLA1NVIXGHzEwWm/yD
qMZW026iFxZseMJP6a4m97nY6EBey+IGArGr+8GyTIvaTGqWsf+sX7dwhgEQ66jxr23Yw8ysMSYO
Z+nyTrPzdO59N1Cq2J7K4qhKoOdKkmlTGoEfXRh7TN/TY9FgN7wsu37QTPMHpUCjMlRoVDVHlYxG
Z/fjEeaPWTPDwMK0HnClEpky8zJ2NG7HH44cV9A1T391uU0Wf0ziNUcC9S23UG9apIn8N2V6VBnu
ScataYTA7FHs5acxjYXTQHk3gJcy7+40ptqQMqzM9uo3IwVTHX7JCIYcAl59ID+RYGOe1PncCxh4
ikat4WjsLQVaP7zY9gy8hXDGw30C2j+/WrltPHJlx8/SDEj4LTVE4kraq6VPxJPipQxlEeeTUw9f
+q0WP65DXE42RIxjiazu7smVsy+8AU2vzvqW2T9RJH1L3G6vIesNIFQx3ir24WTqgjYVcYCW++nw
nY+1Q5XKW7PaSVjDXpxvnbm3KcslrVENTZFRQod45aH0L2f7JkpAgvKKqCza1aabilFZChqMZuQ2
eB8d4xZ7Djx3wLdsiZkGncjiVA0asLCCjxETvIVbwvVfhbrSIaqRYfrr3vr83QhDwdNB2aflWat2
D+4wI5E33oVPMNDNvjPzevtU0UigAc012Sy1r7kUTTecST/luRcu2QGwOIAruCKVhiJRUH7PhX5n
lyWgiwHMPF38SCBzVdOeX3PYSFgmPKRsk0WnZhZrmoA3DvZGuuK/zVMeWEu3jkVT+oH05uTcCKPt
h/5VWJyfVfuxEJuV4ak/kOX5OLHdPTcnU+/ly2SwxZl+2rDhxwrFf0lYHcPmpDiNDnWw9Uji1dvP
3JorCS4PuauIEFadp846bYDXy5n2CbYqhlFQAN/EPnVdJ9yG3Fjy3GQyN1sXOm5Qg0nF3SnC155F
9PVdMfWWYDJ/IpiLhzNTrcoOCUfpdveH06Fu4wzOpBli6KZ2rs+sWlvciI2T5ycVQ8/BDuelvau5
axDPNpLNYaFGTKP+NzCMutTrKa381OA7kM8UW+rcDg9EMw0YuMXTSV5K+lFOPuvkHlWJQrcZhdw+
E69CB9U3sEaGIQi/wBP0dBXSfvMyHK9OFLCvAyYicgEmlxHBUN4QuRDrlaGXUO0gde9cNMrIuLF+
2oKB1tUQ6sCjAsJWDxTysxFmvBEtIqpSnbMSnPjHzoKjLEwVKFxEvvLhZMfbMt0IoYzU/JKVWGL+
BMODI6lab60C1/APGlUPaYfU5ftXqkAtHfmG2zekmDjQn3p+X9CyyKCsWWb0JtXBQqiwqJd8Lehp
FAkMSilshszrkJX1DnF35jkRTWgIJqblPPz4GbrVWV6iGKsNuSW6TfjzSz5djPvCHb4Qg2OBWDn4
li//i64CDTyVHzZHdVSD5lYNmZ9ZR7awhVlcFBjEFst8f58NCorQyztxjNxzaEPcm/F64wV+lKHY
IZOdiGQ+cY5G/K6UN6s+Ixf8yXqGIJiJ4yQUyxC6tjn4yR6MCodNwvSIZIyFISpN11aL3qBib/pl
0kG2nBxVff67PbgJcqf1ZRmpeSwwQ/KU8HEycY+hQqfriM7A1YdYTshMmMEyIwH5bAwTALeh3Wca
JkYAvGWaq7rpuPQBQNh5+iYzWH9p9SCmtDz8btECRsK63TF8dRY8kox0nNKjAyWUFg1GmCbjgBP1
/4XVOlsi7h7qwEwq9hSKeLUaA+m4u44GwKPaVJ446kmDbldAVFi5zxC8cssg90UcBQk7CvOlmyDJ
nmhen8c0cDFgxI3nb7zdWBLmG3bl1Fioy2D9CMGFGvBMStEDMSnpsSRG3bDXkyHp0NzHB/P3Z/uh
NOIhvMleuFp0ROyq56fS22X4wJUq2II2pFrDhFTHHvr7xUS8sIh3LweDTkMJwCZg8KUgPi4Nf4Gq
dSpnQmTNMmnBW74BNV+9aCCr6GV8gv+sY5LmKciTEBLRpjX9El+UFEbRVgtcQBZOub5ip6ddwR35
suA1W2MTwCya49HzR0cliR1WNdP4JsIfj2cVR4VLDAiy4WyR3LejiRZlnQ01LFRQPiOC7pTZBvBX
W1ad+4MaJ83yg4X82/jppqlkbFvyMI4SydGmLSV3Fz+litJnWcdKVNqBsn7NqII3sjuxm8naRe6W
KEv6JHuIonbytBkkcD/JfqBx9DqVD4fgfbd0zqrjp2I2OAAw+RfxayyKNA9/zRFWTMnzpYXJaGuF
VVcMSak9o4XD8I7iLZwfBKYKR0mXNhJMD4Srg6PSHTXiRGMycojBM1y+oHWcTo5SN6jf5/NrrwAV
ptuBLYYmo4IE3bjRNGRbJZNqH8jhHvVut5NI4/8rU3GPOd0bgo80vPz0fNzpThIwwiYrVDlxpld4
kPnUukhEhPRgZAkLtrvMx1XE0+YZXMVtJoW6Zg2I4lYXLYZEpLQBNAEyp78AKkdyUgqP64sevhvp
PDwcuzqInXAl8/LLxSOpN+t2YMz2IH4xIC6rqziZtPWFJYZYSE7xEM2+FvjM00D0aJa/QMn003+F
o6TH5LXDrT8jGY9FK12WnwKIqWm5ouMPtDCBtfjsFvr406YeeHE4gpUaqZ1wkynZ9lCFdZ8Jy1nT
3vn4JtcRSfSWcAllGGdFCWRFsKViyQ5I0/ZJyhjD5Q/XhSFmhlXxuLjfdOs5QghXhIoEXj2OAoS9
aBQzV+UF5rqj9VNDcBiXsbJ+DGcHUvUa4ELu3VCHS+1hqgJn+//CMcffhGB1uB7FAoZMiIg2HAD2
xeG9xszhkLK07ucc9k2COsq8Eo7nQifASU7ICMO9TRIas14/ZASvz0AwqRe8BhyMV3OGSJ9fU691
lO6O/3PD8smP7bGZgb/VvnnfciS+SfWpfaxRATBemeEZpls6IGYZx/9t3xlQb5jVc3s1ndGbuV51
QIqiTOPS0+BAn7PV5yhYuIU5qs4IAD1oYhthm7ZSp5qvLgCi1yBt4CaEYrpCHKlX6hG++uBrw20n
8TxLHchtt26J91bUq6LNLCq3HPUy4F1IFkz8KmfJr7tc+PB647MEsekR53xm5TGZQcBxW/7btkIX
eMFdMl7VOp1ruPqY8D7a6Pi9dQ/2LayLjQxxnwzzYGjfBJSuzuMtyv2NVnzj8qgBN+SmaYZRbfkd
gYPrX2v4EeIZo6hB1AdBZGynXhXp3oCD2pb5gtEcp8JpVzrK6ZUEJ4tVnOrhS4xHOmPCz07Uc3u+
gwDrIDiegw0agvHM7sqoONqFeAvKp6h8MJcn5KR5NRffHQMZUlRa0fhnwYIqteEsBtQ7aZTvO0so
O8X3AgYOWDLdE6EpKr9fgFsOzKd3zXQThrIlwaNc1dnKWXHQZQZp9mmhSO8CN392jh4vEmze14QZ
0ys63veLGOokvZ18gbUVm9uAlldn2Age8z8EgnRqEeveaUK7mR1SOlEuMmiCP5ZQjvFPKX7W5u9I
iEfRq80EeslHUWTmnBHvUX6cZiJ4FGmB+X4mW3IgnaI7BYaFlwvLgHsWKoCLpQAU0Li33gmu/fRv
+3VaQ2I5Ic52dXNnn/ejpq5vxcmfQ+3EYzH0WwjI11s6bhcumAVk2YOQ6Bgcw3hjhJPU/vs2Wwkn
yg0cHygpwSD4nfhzhTh9lzqY+CHOOtGRC0bY3sQqhXt3CNIwWUKJEb0VQbz+bOObnLet5Lhfb2Fh
F7q7ArmtTLZFlByddL5Q714cLUsYVr0kxI8Z3oDbHqntGTpUu+nbUiLDtF68ZsgiIttRTs54uizm
ctH3OYGKIduRvsRspexC/8hPpuyooPxMF8tgSlkT/Sr2FUaVV3TYO2r5kq5g28oZ/lani8Uj5rJv
Bo6A/9fvTQl12AWV9PoOJAf3wH5+W0T38vNq5erhnqhJwxGEPEkK3zlbTzDAq5wmn0BwESN9l3TT
d1sEKEQMq5SkjaO27kM3ziG8I67IBCumnBFUf3iIYcwY/HXO1piCKBCdyJsnf10nc3/6dI1O0x71
jLbUzvDL9JSIqpwPjm4RY5cg4akJKWGgZ9KAJ84ZiRTjFYkVkGkY+LTbtxKz/X8pebwbZwqW2dj6
r/K9rZnMKi8cf4S4LKcRTaYOc7ZEwLYHW/GaWZlJMhc4kzdK4wDzg95gYiUDAiLDSAu9pktNEtQ6
Yh+CvfPap1BI5oKi8sEs4/AbO6zGLNkV6TAXEr0ZChsPfTEKTy/qZJc9owvajxBdupQV5fmfn1VS
dMt09ayvLKo9JmdKNmWTWbHig678eyrCfOt4Qkpmm+9yYh4zcr9kYQyYup5Xeu0VyBGqBpAcdsHS
tKJVGfgZQcBujJ/OxMkWw1+ysmS7MsacdpaKjjYu4r1rmaS6uk1F4qsQi4TXet+8eERFNWc7ybe9
IF8byC/YuTSi5Wk2StJB0Njwrb4LVtJbblKNnxuxgUHkdYvwYKhY308tCYctcJBEQ0P1ndXllZrF
xG4TcXqOO82u1Sej5evKHC9fl/7kbzOVyzBnvtZdQ/ZVAAfi4ezfiPL7b8KRsQaMEBCW+soOO841
UxSpz9RPaTJCvUCW2jLi/SST3O0TFknmdn190WWU4I88ZHrk+OM39OD7wyJoRNTbu8i2ymkdCYOF
hC63oPsoAQ7QAU9kMxr1LNvnyv7a1BBnhuHQOmw65wZs9vMeRytHSga9GuPwgfkGbJLpHLIcGZpG
UJu93BH9uRKxzKhP55cv752S8XhHu8VUXtmuxXMjNPQRALKmOuZDhyrZjFotep6bszzdWpELePHU
oqPyJPZDb9dLvXxLUnhqFK5xAYjA2HaxXTiqZTrUNTw4UP5ZZwrpTuL8tGfBlzFsqIubSTWVmZrW
Kz7HRxRa9QufjUaaF0btg5ZeJIn/YFRtlQm7Az+yPDBaynHBWVCU54C4+4PJR0zqGWYJbHE2nagL
2xl9rYZ6uWq9MxDq+UV1XTvPRBiE7QhkOWCodAE3AyjU0oVsWhm3ArYQxxcbftNsUZuhSHmRDw1g
GgLU6+S/HVdAHlUmkd6jUkf7OHdp7TzGjlkgIjZFv1///cRMKhCh4c9yh9t/4Rqlc7cIvjQ6xHxe
oHpysTAd4l2wHbA/T7mRhjLDi7PD6C22mM818Nxn5sG7adkwjk3yHfnjviWBYt5ZXfbRM2DMOFhk
Ga/jkneWMbgh3mxrsM3fKn70C8G8h4pNeCFKzw/ahEKDfp2olkKrGNEnBuVRC/sNLQElfX/hZPev
zAHVz+UkuXWW2tQiVmnIaKlrnVKRe+C77A4+zAZXnPxlkeHgXXLGAU9pEx8XYvCYeJUX7kTRUYaf
CKvtdac5kftqpN20jFVfzPeUg31wGVN1hlNF1QjsX3pP9rDp4SoidVQBH2WVEYk8FSFQl37akBE6
5e2Mrz0nNvU7b6wq82tN7Y+TAufd8RuTmFM7ff6berrR1ZLk9dPP7FfG+41muRw5YmPXgG3g6rll
1CbO+mfiiJNL2UIJQWnbBJQ4f9endgq1VMmUD/e0IeehC/ddw84Vd6hrg18cOlxKF9aFZzwCbjYb
iRyEBfBALiSv6oExdI5QWMuFuXTKfp3NsdbBqWjMX6pUionRbnl5KPVCfzc/hmJQg0Vgt7kJVWf1
XREhfbo5S3ypKQDhlAFj6P+ZArkmTsXjMj6gwze/IByMLyXqRrVMZCO8g7ws4rAxADTqqXOjOHav
d4nXNICGRY2B4OL2wzifpIiIO9vyoK4EPyimGHHa8Bkb3jlcJJUxp30VhdUwW5ixrckjNWYfjfb7
028V76rlRoeqR6jcjA83IPPqLKbyYNF+ukHHOETH9lr6Vbb/lBcVISQV98RUr6VEyKa9c8380Zlf
/Q05eRRWIFAEjUmMpNXZAK7uKcfCZBc/neoVIQgoK2EekxppnotJnwWrlOC9EPuKd7qOwk86gSjN
mWwJyNCya7p0oTdSisJwfWxdFKa6ujobPJzpEgW2jsxaQTtbFZDtreuq5pLgwnfwlbhV5vw2WVWY
KAqkcZbv5N+12xeMe5vq7UndhIAGvlbgCAtcer7tUoVq3XwXIQByE0VMKh6bcqElNOZEe4BdIe3o
qaWHiXICKcvcSQQd3GvSNoQUX1Pr7MEwZx+SE4mINiJ6H16EnNoe93o9rFc6Alg59IR6vLG63iFC
F5Xjppmp0HQ9mIp9BhQ3JQMa9h9jNwJXPV/X0nNKOYGDSuogGZE6+dhxJ1GCTN5WYG2w5ebDswhH
5cDG7m9V2iGJ6ikv79QMaHCF5qpN7aiL0iKitUDtnKaDeYm1JBPrUf+n0A8DhY4+LudwgVT5qrN5
viVQI725ZYThqkOACCdrjCw+QlhcbqtCdg5VQJKkWHdZuXvkXeT/qOYucnX9r/s3ttlMBXJdCzOE
kQxd6KoQZzHX4m/L9ybxrgjJueRam0sG+6f6c5Gr48vIionrVNGtNN91jYTYgHjpA+7AJsMedpx/
H36Pd6Rk1UneKq3UOr3oOuVYC1BqtmStpPJnO8vF7JKI13JDoZQk8OpoJEFkphFLlI2mr15flk87
iByIOQ2d4gUGcz07aRmwR+I0uiTl46aIGQStjJ4CDmTAL1eVVMDDNWjPRWo34a4SkQkMsyCqWwLN
ppBBM4lbpHvnQ6XcMxMD2bWkWFYvCEdJcjSIAPRv1k9Bc5S87PJpzGkrF0QNIf5KpDd5Rk1vj98X
CPMfDUt7gNAWI1OhFUJGyTEv8hkdHxicqbMvs0ZapANsIeKGSJODqsKwIbGEnoYusMz00REoBEMI
xAIKgbi6iB0uBF4qdefCSa8NyS6RxrXq6Do0PjVujDXw4H3U8Ydh9Gcg9921sYoLhvpVkh/wXLfc
jKhDNKQlkCHabAez1Elstz1+mxRFtbtBHnex2lVwsiYxI1nvqvp9GkAxCTOcNTXKAa5FyWicIdbe
L2/7aEyh/4Lulnl2k7X4ZcOSmqUltWK7PEm/8T1ALbMaiDhkEc9uiiaamgZaQeFkE7owZZcHn8Sx
F7MYCcoM06SUyjqBLbtdCFF625BE6dOLDanv7nL1Q9IpLm1IJRFADnxIlq7xvqsOK77FPWobQFEL
2I0GubwOYE7rxdnaDE/atpkGTpHJQj09zu4fNIQuhOspCETk/5rbivH8Ok/ROGhj4uUoYAq+kxdX
4xgXjMbEimI2Jkdfzj8OjHD/mITJ7AXYg7YHEocJmv01Gvj+2DeIZSnAcR8zAjfMGhrCUaULP/a5
2dMFAHMTdMp9gNcPjADSwnKgZnhmbz7/EN0MUEuohSbQzMDidWF+HDAJFWbtLJ54Ew9IG0FFsmun
Zhwo8sN0mnFMPXzMw6O71xtl16fRQ0ovZqHIJ0BJJ/6R+qFzYw4SsbcPCg4sHQDdk69ochAd8f+l
XjGrKmFGKxKTM6US7TltgmHMsrW7bSkD2u4y7EF6W/Cw+lbEm6H23rHvu/MogQYxSYmolz4INkbE
ouspW5td505B/re/e5FjoJyPpIbqIzaUdGLFNa2a+92+LlK3PicZdl1qg5nSuhsO4Pdp+mgzm8AJ
n8rltaLxwA/+0vzeMvHkZ4Zm3G/z6RZEbsajxQVbeDsR0qWHs3g2tIpf6D/d1YO8IiFm2HNzsmts
cT6Tspjby5o0GyzQVnNfN3Zn+EBBVCmVfdaDWQAcXQkzaisBfb6UUQOYO1y4BwtASt7s4swx3GdQ
n6ptzkYCiywCZis5xwwb7Toqv36nFhH/JJoiP3dYTsqfxempKuK3i4Vs0WNbm4m+urAPUPV7El//
rlk1LtW+Yy9XaDAixiEXrZ935AO+pyRij9L3IR32Ua6H+GvQkhse/ENEZilBfaermQotkgbglEnb
XpeNKSk5SnokyBBUjPJfOqd7lf/YLNVvdSVwtiLsWpIsh9XahkNkAmPxA1uLd7BVfg6fE5vFWT/e
rtwtZMsFBoiB2bKhg3/soREl/dELtafQxExeWAdgjsECEEMDHhzuZr7yX/tjigsRNBuO+W5KMwsR
eZBpgwxKX+86cqSE30nJqsQaxHRdwZaquDwSPmlzEPUXVLZFeKmvZEp4twF4QeEWfIInPGkC4Som
BTD+Wy48iUJEaqvt7ZZ4nNtvl9ko/gmT7Xf/kIVZNwZVdSTVzJRFJwRdJXZMuImj4yDnzEcNUNRX
aWaoXWFuKCxCJ+R3B7CyIxvhm4P5x5s0EiLdAw5mewvN31vlMG8EkmsYBJUI//Pk8F3QxB9UxRH4
02eEXx4qckEslOaliHTDoyi+Rnt5W5LOJ6UwjeaSz0rXd/mgdHW7WPwhwHxwWxctOtox53oxtxW6
MD5fioIly4epWobHor5bZ04Cd8m+tqsSxI1flTBo7ZZ9m0D2aomyJwl4X/PB7fvZWGEYP5gomOCB
Xz9cwy/dJg0la10w/v/Z4PzGG8WoTM6dM9SrHYn444LZBEygwQHsH29lapIStEIlfhrKP5Gl1O14
/cedg9yeeLhfc+70ERYdRdr+8SY0Ha8m6GNBRQVoQrBTEdu75yw+iosPWbX8Xr8NO2/68c16sxDs
kuV0npflAj40K6ZPwJHreAgy7gR+APbRyB1wxBWKfH7EINm0F6KOYK6eqYBM1UeonrELL+NzyksV
waEhmoQR1b1DET9PW1SWh76F39dD6GiW39uc1eFjEpdTtuqg5RZyVhjVbEBBTn6hEVv0lpyBhmks
N7RZLzTecSCNLoM3ht0rgC6JY7q72USHN6UbtrqCVJkyom//cAil7fhMUjwYe95ZbhjWFOeu7ZKQ
czvRF8ySWmW/LlK2Gf0iQgIePhc/flCHE4r+li2CdU5Jn7BR8j48h65UJFPX3OyYFA1kPDbPzclu
aXRDfBX0JxzEGSHqpytpN9b++oI/kjy1jFDzmgpvGVht2uSDFEmUZXzCYT2DGWSvZzLCUDoxUCyx
CVEO80atQHPtDj2+GKkGTZS62TiMF3vagrSaLgmJfct5RO+7xql5FxMqvoQg3Q0rBWZ6rWWe6pUU
QhvZcY1Qntq/UbBB4Kq1iPzJoUDG6i8GTrWyEG4xivHzuCOyF/+JHLFZAUdJbXI47ZrV3CUbDXaG
uRbQboN11O6avIVdprKKpakNAwH7yXIz5eoQ6Vm5G4valiDEwM7ouhdcLMFp/9b3Qa6rGCGJM0zn
WFoQZG1xoVCfaW9H0dmqUnoXUh6NuE4zrfXAvWjO/uCe3WdFejoihEZN9eqbVlnSb8x933oQb+7F
VcOuJKHsymiCxmzO6zUQfDkQ9+QEuPBiwg35H2htQFMps7wj4wjui+ok5w4S/IiPjmatJJ4zTZfs
UpLq+4tbE+Cw9iFrP8BnrvQZl3SoNxTSBmYF0vDqOXKTvWG/Al2q9ioOJBKnvGhdVkO7afpiSXHk
jHPWF3yzQTfZDPDza++xGyWnJTfX82keh0ThY+VEAse/GtshkJuoEo7SaKgRyKK9pGsXVZTtJzry
Ddw5DB7ypREtkYizMxACMaWn0CWJV7oBRfX4Hk/NsggfimD3H5Dd+L65ny4GxrUOJvQuez7ggZC9
+pZS3FUNH5uasgWEqLlze5BT0al+c8LKbbFyHJcuZwfWLdW4/JvvFKHfrX+xkP23Nzbr4QdxN4l8
GBSl6U5RasY0lZx/5seUi1n0IdLjajfG1/bgg6DGlS5CguCpCqfTUZTUBy3koKJB+PRf67ikP1Iw
jpRhEED5UF1j+TskxS1iIm0X3cGuLwT6N6O9wpyHJrBocdobaDXQd3yHQZswaXF24zS5V2+yzuUV
5Jst2/5M29rxKnCPRlQPlFvtID4HDtLMWSkCmUX1sGRZH5XhkW9C72MFU2vK28yguekvw9TDPyKY
yW3YVo0Qo3k3vHb/sPiwTpZpnz5zaDbaUxWAs4ZPXu+6Jst9sf3EogzYWEowf8rMmFOZoYP3v7oN
JdTEQ3Y90Z6ZdzEygysb358SUgpf/kcPtguplba23siZNUFd1dZgdFO4IWDo0XBls9iRobDeXcgW
ojH0FukZJeEffvJSzsy/Sf5cREZAjye7N7D5+Q3r8S7k8LGs0VoiucgWQCk7JzEfqU/s/Pn7HLBr
+trGYectAQ3pCvUhvrbvH/7xkbN5wTvLmDH4wuuAvowr5P0e9opB3uRy2IH0bF2wYQVGwiafb63h
fO5X8LgZDHl8OHJ+81XUx15d+iELViltrRGCNevJ3JwBzI/9WrP4BOux3WJrJ+UWRcGRSSQ9duEu
r99ufdvIDedWWLnfDsE0CFZ75BllMVYBe1B8GxLjCrsDme5kYDwoMy/7VjWTOyZSuJSE8Q5iWxov
scYoLfp1TJs4vePQm4Y+zywz7tBbHvkFVvbz6vcZ2nj5w1zpjAvu/sddodvWXMNUCAhav5gUhIRo
Rmw22cnCqtZM+P+ClI9O83qIdfqp8AxBECg3TgZMztbWcClpVr9C4satKuhbrSoD53YWQ8S7TVdY
RqKr/x/dJ1wev7x+7DvTJ+mhVECiRcmlHYB2c6YkV9wtLxD6p/LLQHVmNRtHyZK/KlMyh0kbn8Wp
QX/u1m8wv5ocUi/Em9UwoqtVahwi2MwcmxooIc1r0n9kUTYhXFkW/Yhh0YZPphcntpKTGGnrTiHe
bXCxUa7yCi/f1uottd/SsT1t7IixdYXqKdsp8A9ZyGv87Q6QpxuyLgqoywP0ZKERR87Zu+NqbDns
K3OC7A9HtVcuew1uLjhrR6pvsMu59gmMEOX4hYgANxmkcTj2uvJH9KhQrtEV1StQpu1XipRyiGYc
18oi3d4EPyOgxMpnn0yPStsA2oUkHcm8oHm1ADeIQPRt0vbDcRUDQuUoRk9Ujhte1E7EHY+drAuk
gmbAoZg+bT6BJh3bgRzSe9DGeoLTQySNpHFdMMy7/CDJ/jveD1vTKsFfdTy7LTt4mXVOPZoWGhGZ
hfHt1UqPr51VE/tvcQfQG+mQWGC/WIje70u4nZePKj8YknSw30iR8XY4h0eKS2VL8AFIJoiGUVXG
XB8xHL6KH0kvDM8pdTcWx32XFmtBSEUPGKbhkiUZHnGvgkB6AknOMIdM5TQ4X1e8tjfVc7Sys2tk
r60TSX6O03VDuTF0a+i1xXb3dxOYSLPpc+IbygRq3k1wchp5C0nYEiiIhj4Bs4kmPnAUzlUWFUGO
YKzzaBb7PZbHomWfhewRrgoOvFyjebvua5CEB2DtMK3Rffzvzwre7VO91ZLafTTG6557G9qeNBbh
Jl3pjdW9RNAT7a9lnP8iyW28fzHD8PIg3cLcGNhe/QaO2vXuHquxsJHvO729uSGp9hzCxd9sUaHw
DwS1QMDlAjQbaxhPV1mgPv/WTET9L8iR3UHHEWGaCv+weCW6mjmH1Vojk8ewT+3qvfVpmV2gBJBr
uwa5E2XL6Ea31I3QU0xZ+tcT/pFNLZkhPdTReTf2rztLOh4xKd5Y/bBGipjoWOpMtnXkASPCq+yk
Fy9zH3v5MiCsTg8G0k1NVyGqDuanD2di+AECh1FT+OizXhoQwHtX2LS+ucC2WqqYkbgeNlRA54Sl
W70htBIKyYjJSHXvh6k9HnfbJhIyRq736+xy3VDDF8Zo+oMixO4seSgE/9ZdzN3SAislzvl3TdZt
RnJXn5SclMJTghwBX0chmvEljkD0kjXSjbFynKhkzo00wTJIM1O1m9b9QSQDNjbjhUBZG7gXO1+s
knSrnB8W2fSB6wHTcrmn1DumfGlsgZd3UROtGGgWd+iGvCLM5wtg6nfxmV12P1dcNXGVoVYZARWT
8+rf+qeIw7XapD7uxxA6cA42BbCDQpkldSAzGhL0j3pXCmbuNy7ibPDP9/qbTkajcU7QTIWzSoUD
BblGJAXQwfhoUNvsSL04jCHA0Fwn0+7MJqfhxEMNhiaIIoTsfn8oFaGPA5M0Y/ov8m67QT8x1+OT
F/xVNL25knYw/xXya6cRCT5mNYeBvLUPLCFfymURqSFloYk9vy0mlwfBnm8h+JP6BQqv/lhXsVHf
WB5RHQ5KcQHjYta0W7pWZH0IP1dwNc83Y2jbhntAmUmgZ7kbONK1IY54gfIVFCJOxxYRxuegKI9v
Cve877FiFR/GSbn7Z6tP+iRHdUhiv6qv0IMrx0VoahgVvArO2fJ0LJhqa04zCjIb9/YtWjmeHpZo
bLr8lQrtImbeLYQi98ca0SS2irVVmztdjQ9CW39rUkJ5wKgdG0BGPfAe4LAppKO3i9FCjZDRfpvZ
aU0q/Zg4YvfSjHbly1O/KONVzIkxut9i38rhuvueF2+5KcCQWhpDWj6m28vx3Nh0SM+ruNxshp2d
kXpu4ZkG4G24sEo3rehCKFo1GEf2SH9TLOfjT1bW1M8PmOuDCs4O3u94E0AbF1kXjuAsGwCt11Lk
SD8v9O/b24NR3yeN7/xU6cqA2F6VfX9egaQa7+ahfH40FwtK2K1uDZDxVjmOmE4PHB6ScCnNUyG2
ziWOOjOP+PsEknyxq9G4UF5YWd3/BY4oyokDfiCfbN8/W5Kj6Z3AVnkZM8qWragMWWa21OgEIp+F
siZb4rX5RWf25q7nFTzwQyVGlqELMBduSJcLf1uQzWr03/UOmg3gHjpmhrQ+gsUZ+4En1+pqFEng
qBl97BttsMjkQEazgPCH9Ax/igV+g0HwjB3culNz6TxhnvKp+/6dURmjuJjUf/Toy5s4jkmbveFO
BiPBulu3BClRKVszCwkLnLRuYpN8UI3RtbLfbNJrQjUWwdRHGhLPIbQfHNML80X80W4Z7d1UHohM
XrHTfh8JfNS4WUL+xCMkoMODJ12vuve51MunfeU75E++ptfU6mros59EbUBlMdSBmZGg30i9xVN6
uz010e5p/tWXYo2wl74Qm1SNZfKOxS/VhAducg7aWsv5bdUY7Dr8s18myEy/y66pq0H3s8iz2Bjq
OxR6FYC2MowAR/K8R4maQEBiu8qVmK/PPAAZiQ+VtzpGPzA7Blc7yPw91MelccCLcJ2VDXcetHM7
4Ymvix+eRWcL2Pt6gTg43FpVmrIY0ZyQMbIreikD4YuAnXS0123HLOA1cg7ECwFZyDcJgf9JHYpK
56jg6FKt0Kr7a7jIxbXafuAZZRXfQJ3Rfb1SF8oHhy6EQOsA9cqaYiRN+5BQaCs+YtLXepgC76Am
ogm2ifNOhS61TkBtWBzDohTWRCRQ6h1vM4U63yypbNu+UGJOeJ7cfz6ooKL7DWEUZCTknsW2nknw
y6ADeqxrO7F/KNqOmMy52gtOg4av18CX4jb9uKBGTLpmCRfXfJgpKJQKxLL0g8r8XVr94uzKYt2N
TTrRfSykomOkr8Y7d1GeaTMKCTwLIgtGs5InfsgtdKA828X0Mt8TdiK9mZR13jfhlwip+FuOBGhu
FrmFtLta9CwCbyi6+7j475iCQFcRv3JUGE43ZtYj+di7+lulnUw5cQThX1rdXFT9vwDRcW6QMJ/h
fEnv7jAwZnNx9Ypc6u1bbuOZYb5DmtlTBCGN8pywi3uS7x0BGgJsTZNHK2jFvV8Ox1o8dd1JNEAB
W06haAgAu2Cev6/kYmL6ZsIJorGJr9vbs32IrZDihs58YRoKdyw31GLLRN9NPa69ncr/cPbtu4va
ClbWD2LEdt6TXj+vdFAEZhnLKSFcaamSLM+6zEkcV0aJYwPEA/JWyXIhJSMhwk14JGaxMjm9XDga
WIcP9g7wplJhpH05JjuenzOUGDN6uJ8DsCl+9Ab/fwUmDfu7Gxf/5mje1ITHWgghbY1P4exgKo/Y
TuLFc4AIjQSFjmERqet2ZcVtFKiZcB/ShWOI64Z5thpgsN8I+sufs76PEaIm3NmVH5Y7x4rO3UTH
OOvXcBJ9jSU3mA74ITeni+lp71Jy17gnOmDTX63Vb6yRhceSqDTkHZvdyACdXvQ0C6blp5oo8PFt
2eUUNJ+IS/aMMCRyqVXgTb8R+tY0+qkVFXx3HTI8GwErxlqDxljOsR9n1SduiS4+/zdTHgREL72X
l93NPGDEg7tSrL+jV4yYzPevaMe1iKnM7WwI+5pRVZXoQAgGZ4s3id642zCAwQ5zSSIQ7L63BrtY
ESP7V+E7i/EgfRkMhk4rU3hidvCwAVZ+Elw9YtxDjQQ0OwUtsxxB+GbFijR4D6lSHDxWqWfXq4aT
Z2/4Y3qNPUsnyqmZav6sXO2S5WTb27Zvl3abaT2ia1+Tm7KrAiEMOyA5GQzgqaH8hjSkg2UWZwNE
FRY0E5ZEtTav0tu91c87R9HjN9jvxdcZcqUQ07bQldu434/64aybL87TWzkwaSGuPxUamYaucpfJ
CkTd6vJ0B4DYt3z8Nnil6wgUtGgW+Gvs/ylrYYJJs2ygjnUBt5GMFGBNXk448eCtFdJK7/ntig8F
jj6YjcbJi/9pjIMR8WCMQ4Vf4XUeRW9/nCZ2t/63bP5WSe9iell9xBoufTN3meRAERF/PUPl6YpT
iIl0NprhHzJ6V9WUeTXpRm/onIoj29AaIC0OBBW6SKZ46FxOrBNTa9y+f8B/nY4G4NisRyireAmX
GE3FcNbs5IXDgD5rd/nJzkhSFe35zrLQ2+ayLf8XYc9LGA/hkdp3zqnChXDzywRKhGLdeWFks5av
xKU+/7pvPO/gLvx74Qy/J1GAZihodsubW/9DFVvk7FxPR9BlA0bQB29m5V84/iF3p4TR6whuLh80
+w9LQMLiIb0hoznm2lAZStLHOgE2NqNBEYtOG/bJCEIwVMw2azUcJ0xm6emrWLdzbZSPIdyPK7rj
QlQ+IIwIe5V5FNxTvIoyJISgpfCfkFdJMAoWTuexdQEfh4R5jqKarx8BACV7QJxeSWbVgMbD6ik8
kV9T8cyHjNW4Gqvv4XojAffS6qjT4vTHihmjQoOtaIIMLX5A39smSUU0Esxwqkl1WxKqBybxvupv
NVPL0DknSvdhceuNnjG7+V57nOHrpl0V8g1fdWQEDF7xjnInVHrrKNH+5CYDzoisKJs1LXSJMC7F
YDCJvBGCCu/5l+LVGIRr/qSQmx7JS8Mq1KileI6cuHqc9/kwrCUApsYS3mNcIDdvsb1WpV1XwQTS
zdMxAvB0wM0C0oSaaEyNPtZrpH+on4+6W0HfszgcYW+EbMTjc1FErEY/d7xfH/XaHJXuHwVG4kih
n08TwlFTQBSaUXeOcnitAPDofPDKLxZlqqvaN1+FPAtdaDkdHwIdRQIUNfuj+WdbB5x7iQIHZauO
sYSPDppwTR5wxwQYCiMkPBkGKsg2lrE5wY+zscvYa6VUYxfUaFHICAaqHrbaq7XaM6A8xfBsAKyQ
gofQnZrOww5+A866WL01P4ytJr/uw+j0d+MByZAzg6cMIOcMX6wY3HbRuwSzdripMjL5sR7YuwCT
Y5hn14iSqR7yVm6oYpvyVo+ka0misyDfg9NqoLdqO3axV5fdEVJ/0gsCF7qUi/xcXdrP+T+yDMI4
OVcJ0Ewi8lw2hoshkZxCBv4UICl3kEgXuo/XLfqVXpikvAs+PvVdZyTjdNntJbvJ6OA8VN4tsc5f
VnQ9+Es2PxMxO/+H75XSAk6RozM/276zAtmJcaBpREfbZTURnhLDeO8kMKsSipIRNRq6Ovljutry
vfCSDGkVMdXRonsAcfm2NaMaC9B9eBErfYIHi7i+Ycs9mhCzdweHZyUPri3VW3rDT1hVum//9ba3
ThgDEI9V254o9xqbHlssi/7XQvCzdVUsurC+i4SHhXXMsHMkoLRYwJbza4TAnmIdRx41m8Y2ry/k
scoS9OdEYvLiZV+ZqYhxGYM/EurFOB2fB1yJBO01UW3RQKEsCMgpeyhnuoTrVwvkwFQgowf64VHG
dxlmbJaQavi+lAgwaL221inWZ+DnLrEZop2ZmHvj3isUcRFGrB7lyTlAa809xPaCeW1hUYH30JoG
fWYKU5hzVoQAu+EBi3hsJ8RiB8ZSx4hRpbgrpqCepHJcPd1Q9vmPOjW3jcffk3RAO4LLEDk+O62/
q5YpiV10gcQicUd+O7ojgmRKhrslAANyVqVdzPqkShRduVXJfb+GzoUNuOZkotl9SLPfY/9CnO5x
+1e4rDiYBWvNnyovxAbhRru/f3yuQbldjnrts2mgRYqvgi+q8JUhaVKeJjvQaRYtdH2T8OddfnNY
0sIEUlhacvYCIor7ZN23ZbAEaSYoiG5dHo6NZfYcztaOgxWnpcYetydw3NC9wFxgqtUSNWaM8UwU
YD2+NhWlLPpee7BLtD6K/I+D4a5fMLW01vL7AvOysBaS1XT+lqEd0c8Iiy4FP3SnlP71QCsA+nwI
i/wL0rnii2eIy9a+FRJWhfEbovpHNmJFarEzbV7HI9Og0g3dY/nmyRU0dPw/6h9ArZ+U3Iom4lPs
JZt4fvXHV10vEZUiphDftEOMx5kmosMIHklDFpK5bdxykjgn9wxeZuafgwqdEzQYI9mnpbBOre7W
EN7is3bohe5Ufn1oViHevI2m2xowwVXp9lW6luJH19O/sIE5spQiPiWI1/UB3y9/MI4G7vkSXLsO
EEpF5Pe8Ha86UPQRtP0U6EKqeAFJIGWIMsNeuPoDsrZAU9l61OA/riQiJf3oeEOJEYAnqMfb/dJJ
wZtALLz8gFFgTG6adnBZ40naij6WDlxVvV3HyY1kOwsV/z+RM/vx0hDCF8OuVLfeptrJxmH4e4/Z
l833LIUnZgid9U4oVkVAwgHahp9j0NJnoP+1jtIIYCqw7ILPL/oROTVxpSgu2XnpeyFjMP7ch+MR
FiEzPAYiiv16ImAxIUn/1YsC2wQEpvHG4rPt6brI9xkMlp/NYR5GOyf/3jgKKzq9rRdakXT/PmVW
hnh3z2dmlsd9tbvGx3gpidqOxBHvqKsDAAYO55ziMR7su6ir7t1o36o0arNa5QzutEtFxBeJX0/K
byrK3F5fhC3vrE/VRZPIFj4W6JgHtP2PUHy366xtRCFL4sAEENJj2OMrXrSCQqkUK/KFjkJ3tr9y
enlSCLv9PlP0Uwe7cbr/SPHK5KrBzjxc4SuFnjuDi09Kcb8jd0zZZ12BU7q0NVUGdEGd8HCiHqjw
qmAJKJhJrd2DZ3hzLyca2d2OBaTSQDj+ePTGux6aI+Rm40tF09GWD9iJQ2We4pZ3VD43NlmYKSFo
6tVgOlOE1AE2zQbRJ6GzgGjp+H7ZpdXomzwspznuOo4VisdQ0Dko6CfD+g1Gg7WLRrscSEcoKuXv
SrEm1JGNXwqid934rUhpj6MUNCEj2vddo/ABnzfdYQPrls+QVUlcWFr+eAbEyuqRJ8aPy+lY6xYn
rWo9sCeRIlpFAM6EeJouPI95OJ6qHxwaq9nso4nqugo7MmOKa4mvmavqFdXdiRe+n4yKL3I0AwMA
qb3F27qD9/Xl0v7ZdbPS/+7amb/qqdFD/8KMH+ccOHTXuXRvxBUMSqiz2vhj8IRPPZBi6BV/3Eg7
INkuniVMjqsmB0NkQv9xAnI4JXj0ePevVxVTCwRD24V8S31lna+amxkWPiaH6+JmN2V3Rz+cMO1a
rf4W7Ib9MvFE0lDNz1mVqZT2sMRJpGdPXxQSwDsEGlpyz/8FEhSb8BNN+14jQbXWLkd/UqwPZmCa
iUI4n+6cB6BNoXQHOlCuq4wV3r/ceaL9gqblK597U7qVUxmDQdFVKQ/9ayl30Z7GPKXQx5qgOZXy
sfDL2d260Fb7tUO7Ihf5b2zWpYmaYyxkdZXiIV1w4JjxFYiQSWWkiyEEnkeLKV98f2+Nb7IkWi6m
vvoldk+wP4D2tGDz3WjEq2AD8jXKZt6eKx/ppUXQlgXuwZzaO/4mFYmtbz/lka1amomHnnA44aAx
X0lj+DM8M28s14dCdTFITtoWd78b+n0oSsaLPRCYyr4+DVXS8pfRpcZq/BSPnA7oyC4k0DIESO8n
1MaD8Hwc6eUGmZGJIOT8/UQfQe3LW9hqcxoetbYqlqOaud0WyHUu27G1Kfs/CHECRk2GrsWDsV5h
nw2jR3rZn8UWhEvdMjnyo/y1DTYvg06qk4NzMCsRubKj2i360t24PED3D/+L8+tEGv9ivqYhuTLH
z9afMosSBhIlboIMompv4SFi/F7IlC3Iga7VBh6cIHjeJeb/bqN87nGZHOp3VMmCLB+EnFgodwZS
tzTjwmWHW+xCJWazkGYQFd3U7e+nn+LkPKanghuhupnPq9npsxuUIfluVocHIIYHaGdihGgJJBVz
SDbmAbSKIx5sydACcOkcNVJ+lBQQdsE+fJtVl+uyEOI0NMgMLWnw+JmPNsSogmU1I2gp5+deQLIO
4ts8+3OrHO4lQMSQPTq9A1mYlXqrrPUrlo8JZdcCee53kNU2jM2+XuezrnPEnIRfEgT/Oe6FbiV5
c3Kq7q1OfejhUHbzLwTQndGAm1WSg68VdCJ5M7wHPEvCjOIiwWV6uYxdZqVQVkrg7AScZaELUkdG
SPcm2TnJtIKZxpwgBoxFeQJYcTu9+nnIbezEbJR1rnGA+wPTtKJa+zd7J10VOJznUQ0p4c2Wfoel
B11Ev6cIJkma5py6s8MFb2lsnMXXNwdo95rdD0aoFx8l1sz9PtSNzpJqVxxn4Z6dc5ebKymPEuXi
3SmgdjTSinIzrv2OJkcRXhlluf9wkVM55BuikgHCEexuh6wWuT+u420BB83BLJU/EmuZZ6MgBg9X
Uxh0+hGaLyYXEwSbsbHfDepzQbDJvAf/qs5FLWddXAZQQ8u0d4le1UnVWj0lAxaPpo4didPszC5a
eNVnIXSMXl1PQ0+zkFE+5J8qXibRtbPMQgCHKPGTawmZTyEHV4TTw/ZhpRTKQotwKktB0Mj8GqhX
Y8RUUaTVB5utfrECw3IpFT9mvFz9QhVPZW6qmiAw5KsViHk9UBeFqWv2xqTK5eFD1sVmRaNL2WZo
lgcm21U7Z/1HLve8fRaXHE+0vF7+WR30ZMTOP7DwN3ChB4ITgDEXngOd2y5C2J+U6dReQlxaLI+Y
iwOpgCQhnASxbtC0bAncs+zO8xKr4adW3b6qN768ZujbG4lKjRf0FpGxPHEQ8lQFVZ9+UbAlnE3s
fvFlf27KnCIsHIwS5pLWdN0IVq1uWJfteNqMCFLPoOnl7JlJi74wfday3Fk457d+tyOdeF6bNNg+
2l5TqVLTo6pYW8sq1zUVbqjapX+bTzrBPy0RdMDlLwP9v5phdkFcgGiYtaLV9X9Vu7+rMs0oy1hW
qGxaBkTRMtvPeOwL7dPECc9QWpx0oi4rVLR0C2wYqM2wmjq3LXtIhvgXuNl2aQ2iyjH4BWd9yhs7
7Kbax+eIl2OvkJ6OXtCNuEXJSkQJx+AAzCEC7S7CU/oTob6ocIQ1F2sZuYkQ3Yc1cBMxJ3+rS2bQ
kXB248hOVLINHqzqXOyk2e9/VkB8OY/G8KP1l9Pv+acsKfh2RStUV45UJHbc39k201f8VA6F5GVU
YuQMKjVxrJNFMLzvGUQs/Z6or7nl8xsF9zqq8W9yjoWtcgklelEWc81I11fKRg9BIcnNZa49u4f8
8J9JPZ7WulFm14dJgl28R1SM/EeB3NMOpFa0eIdlaXqB3fv8N0lcRuWitlWy0vrR3hvhDzvovzVg
/4SpkeXqjIhqtPo5mReKCqR6UpztemS5aicGuv7Q94hJNnOHIX59ZYH/GiagQUFmghdEMqcZGCFs
XvEqWXRrbVsa0pWKbJajxmlxXyB7dIWUahrE9nFCV/98F7rVfjUZM21kcD/SY2TqIIpnl9VbHiec
e6SrY9cPi6exSQ55Chrtj+QjxwCvpmxNF65E9AG0bZOD9PduqBftAadzrFP7iVzQu+ieBAdAGjMR
9p4TJzxmt32NYLe6lDK8YWjJiIHhsbWTQCZ5gIPewY97uUMUmO3DBWmd+Gettpdcw7Ab5p82FzcF
dm2NxUkPQdZpSDanyqAj0Q7DEeb9XFhC7n6K76uR5xBeQkCaPOxr0ao9CSDM0rBIhuB3Qz6PpKeV
Qu3xzve18OOvq1+Mn0Uy6DfSAoFo9rQ+PmirI2II2J4Pi4fO0rrbnhqEhErtjWlX7r7zHm7VDF7R
4IqAwSQYStbbnPm1lclT2vcRvBtdrTOQloOUTGjHDHIPOwDQqY3uVHBudRx8xW9OY/0H/xEAxPL4
BHFIqy2bK2HKlqprLbsPs1L7uBUcZzdwlQpxZKBbv13EddEeo9dcN+NBtOtDJXg0HTqjNCSW0w7j
PhG0Jq4cfAAovl/cktL/k3NQ+U+uP4BANIZZXBohL3Gc0Zo/mIbsTSidkACOkkQbc1RCa01PAARb
cYU6eXMBYcOMyVAnHt98WQNiZEkbqB23r8Ilqrza3wKL3YOcoHZ/dMQUUGsb0Dm0Ps/vl4J5bmXZ
/6H0/E/CNztFI2l7Rap5tLAX1weh1EMYDw2O3Q0oV8T2Hetjj6aLzyVSs6FGkGQ4QXecFT1f9Jar
T44NDWNgr+TpPRIrbdKSmdbmHynTCgxX0QNvXcb5bPHIhPTcvRvCvSZPYzQ2IvaDnyVlMQRBiyia
wRPf5xAHV7GdZibxHUiCA3zJvnGcmRXe9T57PfOK6fvUoPnKQ6VivunNnDLsnNnzmyaSuG7aMe7J
oWMDrcTLBTWcVjDtlOCW1K6hSxQDA0KNjbyR44EtYMzJFUY33o/d+skh+QCH6UBaxSK/5xGJ6hbN
++zCICqwCegIr0q7GxMx77k/5hzXzDrTBUrjIWiFjFUUyIVE3WI7Ea4gv0Y2VpAJ5VeR7e47B+Ya
Axtu83JBHDsyHzsdWFmz/s7eccmjivfCwv2hQ1PbrN5mpDuhYeaFh7AoGq0WCFB5zkSyJkgA8NfA
TYbZYSPOA4cKW0D9WxCVjKutGfVggu3OzzQd0rooj9Z1I5cZ5mq1DjZur/MXTaNOjjLxvq84GT5S
NAq1oU02ONuHj7I3fXnIagpSETiDaF+3X8MX5ONAmB9t8bRg5SrXIzylAIO8b4l4xd5NrUV1Cg8a
cjSHtE89+JZLvnIHVIZgPNz57uazGgJiADHaD5gwHVxmrpqEV2lUQeEQQs/1WU/JEN06QD7xRXs4
MQqx+XNbAnTiZx0RruOVOhjKC5GDBW0avm+v46D6NN4bGO1sOBpEbMD5sFYstkoIuXNppYCGPoOK
OGFRPWQvSQwa1UeMvKQnxyMRbl+GY9/YNtfUSE8lXYAyUod9swmiSHSej+nYuQY53P420R4UCdT/
gm4AzGbYPTN/Xi7FlzkfJaHXt/PtWEuk/rt8JdZNwLrmPPSgMnBRvYWvcnJA+/3/pfRYxYZFt3aQ
N/Ubg+bYFGnVxr4YV6X54fyOHn++vcf5yh+cewi9CnqMk9n9iocfN0vo2PCpnAX/PJMIX/ZJU8NP
oPSxzhT/crKOlK6JOjYw5BbxUg9hKCaKwrofbwK+Sttn4X52eNeXb805yDgKSSXiLXD8yZM33Yxn
1GOy48Jn9kf1QgoIxDSKZM6WEZ/IgUPouN26yLJpTu+xn9OPeW1vXYrLBn9O366qA7z/HkLuBr04
KP9AklVoQzl81RX/YGJrCHqGu4dQE+y2EarA6bRq1tma23VYMMpOoJ9ESfZIys1VK8nf4gVXV/5N
YRpXvx+21F5XMnEak1Z+6v+eq2ymBPCWvpWH3z3pE9LU6x8Q6TctrPoOmSCRQu8XKIeseZDOk+89
c0IJZ37WygDr2Fpx4Xg6j7BGY0lltTZprU1ujc6Wp7ZoTTqwddDUvu05uiV2Od/QJw6E+JwSC0s3
8ggotnVoXqMOJslqcEXtlG8XgKFOVvL9WcxBPrtOwg71A9rsZKpJFZf5Mj1ZYlt3jbFWKtl/O7Tt
oy7+4+ntw5hsilooNRAtuojuhqIoem4yhmw+Lw6g8RnrJvwpylFlC2rnRyymDb/rG55uEF8yeDL9
bnJSxoUKndhcDYjSVbjqHSEDqSLeXYzkfa20BZGRTKmiKGrYVgC5VLJYe846WhaZU9nxNl0OelBZ
YzJOuAcS6vMLVtt/kFDxpwem5q4pKU1VAmH8j2yQnGUEavOB+N5vMw1LBrexqXyKQGfl9Zv9ZeHq
i93PF10Pqd/xsJ6WCH6XHlaV4Ebcj9ROI2aESRUHlbqLL/TjJvmQ7fTDhY7MD34BjZ6rX53OfAta
eWwm970NaNN9f8G1c5arfYLhutZzWvABh1q42gMYmf6wkb798cJGGDbblh/EWpkqqRavgXCImNad
eGxPkfTIZWrR2z5v0pFtOpmWEJZNS3iqIWm3OQnkJ98V3N1VDYzajgj84CcsUqsWYR2bb5ZMtwWl
cwJCuohqCyJFMJGIRWEVSTUxHpWVqLIVkeuf9ZZfsskEXLkYfBM38TE5Ed+FXuz5sf1CGfRBLJCj
9OMDlAFcnL1uzJLfD7MuRoGl23SWgxHc87QtDa8WD45/vEr6zr/aFEcyeAMddCVHrshCPZFkAfyA
Z/qPUqaWYeeRArTCM3mHE0WGaf0kdgR9AhwJvO7VIki2oIyrqSZoDsw+EDDPe9+nyJxCPNtrMyq1
0A4YzNdyCJ4JaDw00q3FAu2r5XoKPMSvt3V0qs/MzO9SpCfFEvW0QKrWkT5b8PmZN0AR3UO5eOth
VHM+j2LPLxiyj8dNBBleWSYBuDvfdOIiB7b/XroiurkhcYXQfQwDAEPwn9R8Mu8uVTxEaik2hUVM
N9QTi8zrM9oXgOxPZ+uZo2M1VIf8r9QPz0otqEUAlc07FA6XKV2itqfDTI/Wckx0EWxnfimKFNMN
dU14Uv6tNhhW7NEcF0ms2i4O/WW5HdP7aUlTjR+jvfgmVOBBC3mBqGWmFFfijh5mryLZR/cXdqzf
zGo9N+Ja12WI0NsdfdjUIKm8jotOXIb5k2kSGZZpQ/1cLyCA7vgV4h8WGKOSO0TgwU3G9cFxLj+m
AP0NCUnaXd9Z5e0qG5N1PhVzc+GO6pfjiWtEcEvo1h8pQiqC3+EorGysBNnXNuxQlPl5n65dJ8Wa
iMhNi8mYRS4ht6yK58HuQVucg/dPyU91sFPndOGmkHSP1Vz4g/juvvJqhA/t5WmXW0rJnsefNtqW
kE0K5Cvqqr8y/kyIv5MlwDFM7TcXkpfssMviwMR0VGoKswpndeeYpiS2q7v5DUYiGllJq3y04xcl
3IiQBs0YkrBFf+HEDRqWi1+1X4xDw5qc8oaPkVGdVh5d8MuyyDAHn6HMR3rB0UztSijFPy1yjMaq
rHoxZZd0zMLqsR68B1ef/UiHWWLaT59ly0KOV4fQ1ap4TDbakKIVN4popc9adkeovrqyvsTmcTOK
GhK+0S4WXzVjPQCA24zOc4YxPm0+BLJ8YFK5oTG4GW+6nZ/piK9OXV1iyDAs0sdl4rigaHQ70wCb
u+e9HUnFTFLyiu3tvAwM/sZYiPME0rzm8MluvxUTVOu+kdGLysLznk5Lme/IIYoEPZdOgOIYkFQa
gPzSwodZL3p/PUnnY9Sw1ku0V8ZpOKFxNXzCPnqFNSAe0xOOKDKcKbID0EsP4x3i1PoKLa0uniJn
QKvaa7rFC/Tr7gesBdYmoqiB083Ew9uxsDKlTZJFpbzitYWUqq5hAwKoXRHjotshwEJpYWZehAkW
UXgKilwfCQIMFaidRsVXmmk4BVr9OGBJHQPolaqBEl3H//ecG1gurFJOw7pybpwDGuBcOcMc6zQc
hxUU1Yqlmm8p2nIGV2Kzq+XCBLw4puKqV7QvvCnKBoxfHZUOCjitAuMPZ/Sa825gHEiBzm3Dw9Pe
JKKgqAsIlcjy10jlsL/u1up7RS7wrSKfyccOgRv6FtVgxxmfwCVll4B7cjgjyws/GxjnQykEOau+
WA7UzhY0vbQQERWCw3uPy5iwUAN5Alvl/zB1KEO6VRqG4sUlK1sBeAXY+EmDqbYH3Htucq79oiW5
L+sI3ZHDpS5QjF78YypDvw0fRlmvksOyydYQh7nD312AUcy/4tQCdb9a3TL7eKH+I5kwIgwsBb4m
fX1BrgaX6xvsFHVpaqGYY0dFHRCOH952wtyMm+9kMXjjDDH47On/KWupQWkIXrLvAD7AlN1Jca8z
XzpcYwKO7Y2iIKxx1xdjqyJccYsFrRcrNs17D0TXq/ntxO78ofC9WW4iGk55yMJKPHIlNQGHMoHH
zNhE24vc4Q3AYedOAhT3B8MdfZ4Eu0nweV4UP7NTSHKso7/c5hBZaXCzliUuZTHyi48cBtaL/Lcq
evBuDR9zc+SfUUEIz3BSSNFYJmFDmDBO4bkOsvpywLL+fnyOkKbYhExlwD8gprfLIMVMKA411P1w
xosij+BiDh/LQECeuIa4SHC3gxTswsVwA5nlrVQLuAG3dtZFJ0YprJs6OnyYfLDzQHAnadocjR57
d5yJZyvMFxLOVhusu29cRQlIXTpTos8JtaKaAtiE4EQpBV19jZYmtEkfzo7ZznHGi0a/BAlbWq0v
HJmK+DVBRxXct2vS8d63ScM0w4jVQtKB24GAn56A7LQG3g431iN+ge7lERov6VfxUu97WVhqtuVH
QmTNbuKmAf0oQTVNzyAqfgsHTHisPn6E4vxmQUfz0zXfPv69J5+qAqrkNmNmCqzGGvrNgEKv1EGf
MohVTzslAT/7thtr/AiYgIkDYLaW+G0Nn0gjS9xZI7nCzE0pDlASbYG9qn7kHFuFPByNstnliZWy
Qhu6R0DAhBVBoFNPaBvZdumtg4NxEbp9eAMNPNsv7W1gdicyMr0N9oDYKVbxbk5bsU5Y+d5kB0Hb
gz35OyJWFZQ9wOlDdH07NOYiht1/0BhbRhEktbfuspyHFE/RNYP6owcZtruK39rVEiaKNJb9WqAy
XhLDNXrFqm1FTrg7u7YP3D1g1Nt9Od1s/g5L6ZALQ25MvXpe0WcKrEPfGXgkOWwztwxDalwX93Sx
DkwnroffDWt2NxTMDrFu9bVRZWwem8hDUo8ZCNzHgxxnLDjIGUJy3hScCZTtRsGVu/L5bpLGztev
VGSmT57hxO62Mdo68K7qsjAyL6mcK16BjsJQcHsDsNk7QNWCcJWRzipEGoFZcedun+WvExkBCFcx
kHAlH2jyTx+5sNR5NurjrXdDLwsgInv0cMq+8e3cqyFS+r70lgO8O8dw3rpwdlZeCZ/iHBsulQS4
6xNPb/5aB/I+iEiZtnr5VexTzKkm+3wHPcK5qtdcoIUDlcFRyf6ZHcPA3ucB2RYl7g+9daCPejZ9
GRRlz+/wtYdcq2Px2DJ9eNzLtKz63Je/a32hdcV0bLLg6NcO/Hf0joICwWZbdYeUfXi5RzDZFIjO
Qfql3uXppJ+61eBZyHeYEaf6FUg6+mNPBj7W9+AJUvzDgaK1BdNjByGlMLPm1GdNrwe1pt/SNO8c
aUQzuGHjy9bOurVxPIHcYnCW0GYbO9QZW/IgVkVwK7wQFNgEv9aQof6KGoDS/IqSPPfyQsio2i4G
rB8LPR4HL53XM72JiGHrTxQIR2a1juhrxVQv561fbQXULX5VTtN/wX6aSnQZLlCoXtGMsHGAHUpn
/Xbrmh7z6ODkj02hC5+/yOzJl354wIF259yFMtVlpvNgO2t51rj8gsEHdbZsIxQ2hAQ4/cngZeCW
fhGvW7QRw8YBapzZOsGRVfSTKg65myi5IB/KRx8m7CcJ9KLfxsyYu6l7aLIyRiQcM8h0ykojs5LV
qHarjg889uMUe7TwHcenVHLqP6vx8PBQphCTE/c1O4bYcdnlINo9Fiy7NflCQj6oMIjAXPkiqRwa
9HB+Kge31/hvaobeoyBPrhspGRIRva/tTuas0ABX/6Q1mgOuKbemUQKaghPL73rpeRBadXIKypXH
QHC0tFhvO4VBsgJtWSMVD8e6+v13pNQoMyuM0CzoF0sNMsZKUc8HS5TMwsIOgHSXyeCNIGZ52RHq
6bfLDrvkxxc5oYKxTxPRMIzXalsijtX22NcmH5WkHDaZ4LFaHqi6erWUBQQ0NEsWbup5ujssccjP
x9dXiv/7lKWQKo5ha+NqZYDgIaIfTu+xpfcyENNDqrE++gbtC1uoN1G7OucrCh022dBlCnelWxUw
I/bgC+NlIqhPiRLP8ybVL3jz1py4eRmkmdbjUrksBV83f7Gvn/YarmE8qMYajoSiR0y6gHKiejaZ
3cLZXC2jl3J/9b/LU3Gt6EcHt5caKb4X9oU/r7lXMJaj7rAz+tDWCk7N+Fq4ZMplJmSAEwrrFQqp
BZWGMsl/jRQ2q18Y9szIEaM2AJmpw/HRrTLt4dSFKRxVULygI21TBlrMqYN7uCi4TTbIUwKQeoTZ
wrFdURvlk+4aT4hKsuvFcMmCHv/t/gUZmHRXV/WwEueP9CtHLZqp+hlP3U+iTjhToGxy0KyCXqyw
pzSexqM+VudqfrbquidJphyw8CfpD9mRZ1E0E5m+8459Pdi0DU6ypRMAJIKPbZF9wJ++o282U0Ib
YGPODZwIsL2mHRYQMsRN3TuQ56wv1PVgRNUBFY5cZ6TkhpoMCoipiUFyOOa/S2ZfXSVevAYY3rYp
DB2WXInTFCuXDs+93Vx54pCbLI0YK9Mk8tFydXivEj3V/yby9wqecusDKTBmIxMtCg3MTD7wqOk/
Rqw1DCH4G3dYZZsnnP8v58AHPIN56ecfVBCjOUnGjenPapiON03zRZxsPOOio53ZxCZwlcNztg8S
8NVSc3V/r1m5KVHok++/3zJnTiZce3woTseWR/9obymKBJWsnkZP4CDimkWDHvU8oyv/qjU9RmcX
1tQpIRoXATc0yB8C3groMTlQlAj/VvOzGN4UkaXTI6k+TthPzJoTyedZbn6Cq8z2kIo4pcqo0ozG
+bJqxVbmf98Nr/8VpjQ1tEOoeZ/5pvsskOM7YZBGcTiYM8q6Rh7DRYJgl6COhEnYFxgdVaCDbkFo
6/mQZOTbYGFtDVX5RaZrm1HvGaxVZ6JNsbeZGW8Ei2OFEMMauHvq8QUcduURIqz2ZCU9x4GlH4l6
ta+C0jwW6/3tP6OunD5QFYujSSH4a/nz83nYAhEGSqhLM+7zk+KRanzobHs5srdKOiKOD7Mn0Ni4
rhvrnLvucVot/X+jAH7UAjlPR3zBWGr006ph/N6VwU2UZ0Uhlf4NyRrgBu/B57t3fH2SCE7skPdw
kCzz7FK60vcZRGoHhwuukZjrAvCgBgzsAtbjheljtBX1kwlWtrvtmiXFDoMWcRK//fXmJwMce6E+
sD2s4EOtngT26eUEgryLoOQd7Q6dg8lduBY2VA2obmyJg0jFkY3lRXI38I1ocncQxDSs80JDDNwc
umh9D1DA7HgmPTrH4J1K/4cSTyiL6Q7APZpJ9lPak+J6dEjVckk8xQl4mCLRpUxhdomU1diF7v96
W6rotKTunDnbEZO/ZL77ZD8/AeDBjrQk5j9dGrW+Ag7TvOvLEryotS/6YlyiPxcwlLIHCNOnyVkc
aYERI4p3rPjerkGzXhdor4KOEXfXFQY7oTbnELbWYweoi57AKNadS5GqYYTgmATN90UvIa/fKKZV
yShsTC3DyCIXp1ctX4VdqGWGFoTktsLk7Bp+vkvINzx+lMeERbNhJ0lQ2Ibj30v4a1ZSPb69k2Rl
oEzZAGN4mhs+FIAxlsJ5xB6KuMOL4vTyOwCJCRIh/fcx/2JnL5sAFfu9qVce2xhVoShPsWJrUU8x
8ylRivJUzQ1wXPQRiLSzUQbP+kIGJf0+VmmpKsE4uoGIXYI9DW+m5X1ULoKbMWZsBLGdu8+lhwYM
rX63Zh0hyA00fyhtp7V770OWM0gXIbrcCGNupzk4E1AZV3+isxMWzHr+ouLsBnHf/pDDMf7JIdUP
v5L9h8q2DIEN9rxhNvbasgJkm9H0lbKiiHDo63Z9a64gbY6dqZERWospUpj9VCeONbYyxEik1g8Q
TwFLLIV7XJgpjk8/wzXDkI62jBxq1ajQMXFc8e7r11Gve/DyyV3LwyEmEkosmJLafQjRVo1FN/o7
6uc+iNaK8+5ievSxrQ881EZ2ebnlYnPyOZRrUn67ZqCZZA8JQavwYw0nkUJVjJt262P9Rb6StShO
SJdwKBlC6Hcm9u86TIKC0Ocsq+MFFBtPn/W0HBfSvPJZKuGSw+Y4J6j+Gsh4v46E82RPmlIsyx/x
wWXAfAl6CnQ7fGGN2gzuzBnNY9Czf02dkv0j1Ev2fvrn/yGDwYkQ4gYH4gqma+PmaGcfoN7NkEqu
mDaublw/z8ZdFyNw0YBr1LKBn73FO4sOeYd4/yuddsHkd0xeApoGThAIolWrjS7I6LWwo2wEfnSW
C8ePjrM7A437gXUIBtSMGVr574XpUjP4JmcEHgYh6N7nf2TVv9z/cBobnbSny8FZXGx/nB5GRwTV
BjT4xhZKUHcoAXpoYowbk4kV3KUrKvFo8PUhiBV5+GwRmuEdgtG8oFcTLkNqBXZa5XP2oc/45Zix
Rrboz+uK8+86j5ar9Tj50oh94qMKPFjs4Zssmc+4uXxHolwnXydMqpAn0TgqINCF80da9e9ME2LQ
19PV6615ch/tz/hYg3qV+WaWJhNuq4v7Hy8nMTZ79eAtmn/UfIoCKox/H02/bYTjg+BvaFRsHSmz
dQPM1FYZ+/JwybIMCG2sr9v7OFbS5+AZArMHuFKYtYN0l1+9jxAdyaG/uhbnprdr6NG/cyAcAXlc
04ocdtyfCTzdtwM7Iy67NKBtbDusNswIg6pvlTtaRWkiNRfOV0RLSeY5jNSobo9bodukHfAKv1Ap
zEMxK/ZFVUp6mw3Ieny9WgwGZXbVTJE5HlTtoP5j7UViRq+79yUboc/k2UzL4oulF0BUAJshOnMb
VsTkPILhY8P3k/RqJjjS1mzYpSFEeoJ2n3R1of7ZBg32WpER1aB2oy414yvq+8ijWQtY7aR+T9Nc
eFlfqgrI2yLNjoSQzPiq6iayU9ItJgJOcx6y3UG2Gyt1SzGDOtTLoYNFmVtyFBOWdjIP6GeWOmS5
1a3wfvWbCF7eV9A6IP6thMiw1jOzcdWw94mUzWvsIiP7lZJqyjd2R9Vn+rGLef2MpFSk+UTYv87P
0WKua++krsLZpafw/NNGQa5m6QxG7yX1UE0XgDuo9AnSXS+AKF5HZ3ranml7nGIAKWVoA+MQS3IV
F+dhAkqPvSIj7IEt2OkDjjzLR96D2o1aMIpgx/4fn6gca4XIx3ej0iSrs0UK0jmjBk9j95kz3pzK
Wo6x2Rvc6f7PkQ6Undv2kYX6y7OMYYa1Nx7CalwiF5jdWfl0UBnUSr9m5IDPfR/g6J2jwU9n2uU5
95KoAEUdNn1V75GJZhXct0kp55NK1UGxToolfhG8ax70BCkKqiTlNWljDYAVDYrFeSUGr6GPseyD
JL4QRjxEj08DLUgarH9u3ep0X728IFK+QHjF10e+m8OA+jATuGLI8L4P42CvI9dpOH0RgpqUZ42o
hv79o5PHruEb5b86QtirxDOxjFm0Nto9FctyR3PTL3F4FY3EYMI/rWDgS5hUMgcs0Kz+orcCHJ5s
MuWOplSiZCEh3B6ZI91acK+ZRSJXULrPVym9UPUM0drRn4Iw1XixuTSebrIMK9/Y84bq0qlpSg1y
ubvAKmZyrRAYfb1yDBkVgNgzE+msBoEdmJjd1aYk8qLYixEvhDut72VNgXGErkclxKhpD3SM3OJS
8hVmoExBIISWxhseach6eubDfvMjl3EIK6hUeiBedbGRHjwDOvMGmPtWRg44Yju/mMTHsjltJTZt
5tmQBRMS0H25f4E3R6gttcYRw4sqRFICVgxixr5cSJmnqpOrR8gdjTnjzzOz+LSar82+mzPAZLqd
z2WO49fBGYTzmczXwLjR1yS3XJhf9KkJixQRquNlRgMEDfNUpQkXfv7amwkVP6p5phSYMNYr6s9c
H4yZz/dHBUbHtAB6HwZ1tmSIjO/zJukRYNwSRSsyZu7Tl03/NLM7orFbqJLv5rGezesdSSvFMSEU
03Izee9TuNYeU0WLyL29jqmXwPH0tXsJp3tACQen8HdqdPqf3wkjCud4SCjqPOurw44THNKHTt1j
FZHKyABKuJOP3h+jaPbvdLDfsg9svLKO8iaskf18kMouqC4orogc2gsvgbKPQ3eddydI18qEYJQa
C9vdK/HREXJIPWmW3nzcvES1COhuF28nzT6tWHluIzI8Z32rfL7CjQlUA3dSloHnAJYoILMxMlVE
j0v8O5BWrEZgFnt0k5YRQqZ1hV8nEg2T3FQmhHfSS27rMQIYHpacHXwKW36RVF47D6ypf9rRLVC8
1BSMx/LeEhrOMNK4FQlvGw5u5lK//sDx9U8N6odVr8K16HwXXubTz3qQQlsqp9fKNzeq8+7YvZLd
PanpTBZFSX7ckf6JiFDMdErVoFxkGeJ5rAdos7oZbOJduD1M4GCyTPYwEBu1gf/RJd4xmWOsVHsd
7S5AQd+Rbvo6n5wfVm4fl8YSwgw3fV8lKsKjjpZAsR/tQZ8QM/THi+llZiW03erVKpDAS4Qsz7Yh
5G9i60eqWBDwjYkvUxzl/17GUPHv5ZcOpQFbK4NslvSgSf3mwF/AvZgL1n667CV2mdWPnOaOBURI
yYPR3YWNc80ZyKe/PJqS9wzdBUdj5+w9sZWYsB5NjpuP8hFaiBO22ms0yp1JPB3kWNC0JGLFIh9q
8xfhjM3MmqEL7IR8uGKSlIShWuzCM/HUJ96OkYzMOz6nl4voBYjOPWrVPbExom592FPFIIw5k2Fk
xzEM5M18N/3NKZi2/O1Dj7IcTwR0u2G+Y07MHoFj5QghDY32rdyYsJw1cZoMAGTkKx3Blw1udvuL
GBYpc5qxKNLWCPEOy7h5yIg9HjCYC+xmJLMo49cjCLPDemU+AYY3ME5lvmrQb8xfmtU4Ohe3Vs93
Zxu7eTSZ6H4u9e4Ywdj7z3oScKt5grbU9Tmkz9Qnwu8YxdKTkjD2u+45yJwP+2oI/ch2rGXZ8Ap1
pkykrrAIF3exCX7ZNvWws7iNxfYWw+iKlCqkJ3zGoQLJIqC2AtfTXs7XZNQkuTijrxRgC46fuNzo
Y/pYO7CvX9O99tgnuueoZQM944bGPMpcMX8F2jLnNivFqv7fb58Hyk0ng6/ViArAkzi0q5W3d6Bt
F9lIiT4KUX2qjrleK9Moc/BuG3TO+qumJMHlTk2+VxGDVSZs0dVXmx698MhNyymg34iuvJdhQsng
ngVkN8WamM0oUJPe/V97Px0vzneX5PvYhx0UnwBVhNaQ+JohmK5I8TIiry596WQsbuehYZIWN312
YAkWQEO0GwNM6kRVauN8hDOJRrV2BJb4upJKLkPmQwRmEPSp/BCMUr/0sMKgY66RAsqqOWsYiz7K
aKw+7embRUj2lM8l0xCmGD6mCrlh/zFIyjHRT8XPG02KbezwslxcJzxMiFhEQW7AyrNaYosWHMHC
SNdHSyBy78++D+nALXNBIT7RC80gSI8KWmBX96c3g1iTYgGnDzhJKxkSLLPoAsH6ILeEGantmtQm
9FNScK7nAyg+CazilvCA2WltzQOZFMVlgVSKFgMeRwTxpvHR7JN37nwQj/VR7XbTd84yfsxHQrLb
q2J2pKNnSMc/TcMsYtmz4ardOLtaPL3GQM5icLeAHLVRBRqRirpZ5L6+mupfcHTgIdJFG0QjkyQO
NZCEYv1mPoHviFnLdR0tjHwzkcMzJi55hqW6f9fkBZakWFF5yZwRXdkorSaZrda/BcICQKHBiRIF
ybVo0L/jWSWDnN0SyQzY0ijs83MXbNz7Xzvgz5oxWQeOHv2xlMEHnW9n3rXRZbTkk1LZOPv7nE4G
fTt4xdSFJnjTNmQ0i7EdSUDerSfz53zbLGNxN49svatHAPEJ5q/Ut7EHxQUe3r4IVxxNBrSureBv
IkW9wM754cvKe//h5qW7P+kg4/KLoCqE+W2TPkteLst//Az0j2KGk9PzGcdn6foovkm+rSdMKol4
jH7UWxpcCkH20SL0t9FMZexxJKg5YcmaNZg1IrEE+97fk5p7B4L15SPNYbjvAvlEe6yp+aCANYmL
tiifsEFDGSbn76OZzhNWqqql0bmS1/ilCR8XHcfnYXDQH/Wg5u+Q38NeqohckC42jdx+DLcNpAkB
K3fgFQd+aV5eSzyNKrKSx+FKgZuCe+dxm9e0Rn3233g8pMXmi6NVGVDFMA8+YjyKEK5YxAUGf39A
2n9i+d1TERja9EkKN11gC6eP9KY0duX3eR6K/Rn6otM74qKx8TWqG8La19aKo5E+xjC0R7ad37lE
nfAAVneaXv2WRcrk2YvkyfbszVR+twxBcNMSTYjN5iw3yc5uM662jCtWztluWYSVmd/QmbMEuQDu
PebhFhUGR/QZCXb94GV4h5B5XzcSPko2c2xSDE4fQjHCqvY1AIMTHjmV1zEP5ewQtwQD8ToYSwct
c/CGBEKXU1NIO8sUr8dGlFPbA6UD4A/wQG+39h9R6M1j1pc5xotLLkyy0ULvm6hemHOFnVV2W5N4
+Ri8oUdrA07gwvBKNNNACPJuijD5Mraw043lkNz6a1DhJBdjXI1412tfgXAM6FiWZ7BqyYXjh95+
f23neDguSDkEnCnkBJr2zgy8utSaEjHAiHPHI3eL2wrYG6E6yp9YTnoaadaS7yTJHkW+AUo3EcWG
XQODxSY5b9x5zQ3bbY++Tc+2dLVs0YsD/tpoTyPHAJ8sAnSDEv3XKKG+Iva23U7dvWO/a5Yl2lUG
MKSW33iUnPCo3lnpCYvGee4xkAXV1tTrEOmpaUEYLS1LqQmHuLOqXvE/001dxW5TdrYdmuarJYMB
25UO3ucU0AfCTN42h60JuXVRgmGcS5Rkwrav4wYztdTq3je8LD/OJGFc3vZz2WcHDgoh5AGF39yJ
Vm4ELgf491f4cGu01PigVgaLQx72dS+7c2e7nAIwUpT5bEBs87fB6PrrA7h3F+HqUkg5pOHjy9e8
VNlxSSUuTMAJ64/i8tKXPXOGzRp2aaCYYkJAml9QRpZYWil8+gPhbLdETeT8mepVb9rhLIzGL8cS
3uHld5ggTz2vsVfSxHwRW+FccGEDid5K6SRiqsU+otkVVFdsP+Tayc4EnP+2i2m84zB+XsEqFf5w
6wcOBaen+zdhcbBDdrVYz2MzwfEvOj4jLciiu+EhP+LAOfy6LzexiJjACdBoL7HC2CDiulfvXZbs
FmqTTMPbE86ldXoAZgPmUXp+RdI4nhGvahUAu7HHfRGOnWvtmrW3uJ04anqIjUs3cnEumIyml+c/
zKSNzL4LbqSzs2YWgScPTJNZihd2MTNYdbey7LeAEhinJgsKPBZ+HUB+ZPoJ+LVxc2XqX8yxqnG7
9uQ128nxyvckektGkFngiuYSeCt2u1zl480bQ62d/J8AkcuCSeh9Edcx+xn6jyae1Y5rQSZI8laP
xBl5G8hCcrwaFp0CGqgFGdMIsE31etyz2YXxIoivzYlW0s2lLi4jwrgjhlq02znHSXaVom4I/ean
gW+GL3lFKrDj80eEXNZd+9VztClW1qKkTPJzq6y4tS1lVTqL/1+7Sc29o4PeINtuWDqRyeb9qwOm
yNMZ5t0McfjeanRNYYqu6vTKBHFyvsUyPjR237XiHFLE46H5gz6Re0GhW7LfxqQ6RCFlrp4yXFG9
pXoJMC5eDGZbrM/Av1qfctJ06fTtSRw2vhlDwfxqeHvRxo6DS+Nl7chp00ntc0EPb8eUxBoDxsi2
N/VJcMw91HPwfR0GD4PTx+rN0tpjKpw2Vfe35LUmrqHaSP1Cb6JDsDNL8x7DP1yL4oIqpy4Qe5la
nqai256OSKjKxjB03p8cWycJvjPuUDN7CxylM5cVvQGSfAaCH20FGI/4U8973Z3+GOOBAsKoLwfm
kD5KEayt8/ey4gVprmyXczdhc/tReOLrP6zUugDABls6BYFO7O3S8qsGGqORcTc2wU0jZtlfceql
ketM6oIwAEw6Un6d2ZraLzzsbquIE+Nef1X896XOXFOEnVrq6wjVDVWqNtIcZsoFCfrJnLxX89CV
CAdUPNooKerheKhUeCiuGMtm3tx79azpuFS+DJViUmNyII3qD2iHL02rAs5/lS3mw81PeubKdh61
qrnWh590j9TaV6JyatJBA6510ydLGiDxiDTMuOmvipB66mea09NrQboBpEoH/VayiqfOx6BAtjG1
TpB2glzaEUvF1qT3saw0vaSkjxc0Stj5aYJ2adSlwMD+ey3++PDfev02Nzz6fupQha1tJ6Y17aSW
4PskVUBa/kasBjvgIZ+iC+nt7n7FIljQbX9u+K8LH2iNfHBdjeAjlQ5DAkj+XUHhd2s/58V+mw+V
c1K9BEp7U7EmK+4yriV3RN8899Ewp6qbdrygVl20Z9UFStBI7PxctZaLaYyT4hYYLdh2CvFGCJM4
teF2+gFb7P4RLZI57txOkMR/V72ieJNNaDsgEFKXqrVGnbWLmvCAZD2NvnHplVQarFW1q8Yll2kF
AKwjXp9GdQUPLJEhUj8pAqhRJbw9FEWOWlT0HEzz+8iK9h1CHa6FbErjmFNLv4UNJ6lecym74vrO
b1D4u297o+r1t2VBOQG+gh4d3w3QrwFY0opNORrn3cp0eIa3I9pMxx7qTjnW7PM/FPbxHl3U0nMP
QM3yDPI8Wte+uDqiD+Rba8mBlL4mELY5NY9QRbx9X/9vpbZas3kA6xglUbw6AeQkZH0EmnCgrSOt
Zx3n/YXkX5S3+fmHoIjeD63dzCEj2PML5wTOsyroIShLu1Js6ZE4hjpTXppK+KvxRwdvgYesMrYq
3vqEa0wMHDKMzmpVwf6ZCb2ZFuOzq++B58adS9+qoryTwC4mUZFGXQ+FXEgbznrggwgSernqFNJC
PkWgocbzOaoxW9iZ1IdQ933MnznoowFV7TALGevde89ANKyQ192WSEyVMQDXjhZ1KDRbbwhpUS0O
/02yk3AsXbeoJGE6nSnkUOkByeFBNEm+OENKLFjfXKoWwBTIChYLcpsG2k9kd/FqpjdzDxXbqNa6
QrHLtKke/DhRj0J8xb7iqZBYiMEqnxEFDWHvqYeVX0cBJ0wnljFcZchdHT1AqVS87JKofX12eKQv
vubVMYjPQXdC0edZdaamfsHcgF96IUgjg41KOwWiXXZgHjN0IumkmJPDw3dMweBPE7eGiTKjlkMs
XE7d+0Q2I+ZX8VPYwAJZYIJ3SJpLEvy97hky+r9hRquqigKFdOHj5I3ohowyq2NcIQVHj0CO1Toi
gaBzZUBy1rQJgEVQYR2OUePKs0i/455/klmvldkiUvWjnK0ItF4n1l6RXoTw4D9vrMSddfS1Lvlv
b5KnZxDu0sMCXX+XfyxslRTf2RIFgT0GNzMhHthiGG8LpAB5mydQREZjdUiqlVE2jklVK5isWU3Q
fqINk9mpiEVXx+msfPyel9dmleWjeXd66vPQQQrOploS21UCRPY4ef2OBlMd5k0PtPtJUcftr9fp
6Sweqx/75Znb3xQi6I7P18F2q6IjTCPH6TFT+AJ/Y74rfR1M4NObzXmzgs2nAJMABmXzHmQDF3k+
R8v31uqSBaJ73CQSsz1iSxtaDvleAYyZ0hfWy9khJnFjplZuit2tz3EUkLp8TMOQb8EHobZ8/eTv
kd/H3xgeHTGQV99i2rfRbU0ctODWF1hzCULEwnPHGM56MbvpHvYQkSYWSnSc+zFq91okHhjpSj90
T1+DldtWcPTCL0LC9OV/cK8e59XX4JudXSxtGlbaAVi5mmIzlkFnW4b13C8GYbTrgYzC0HIIjjfk
mu3NFq/m+NWC2C3ufBiS+pBf8nGLgMxmFyxTpRDmCg8WYHFcm011BF/2PHkqq0Ofzk2Gg5UnfCk7
87VyXxGpPAEkyXmOyTS4TffHC6emvY5KnSJnxQOS3brzWsBoMYx6fxU7wqGqcfNLdoQ5zkvvhYfq
wMd7Jp7r3N5KY9symAK8ZAzBDZI0e6jLFhDLoFBZe97W6A8RH+GqluT7gjVR/2oTKvR+V/40Gk2q
RTiNx/d8gJfjVpfEQXfxuy/vQuh7omWrV+rk1ZhTacE1WTLGEls9VNe2XzM9fFjVaYk55fRZahxh
djxDmiam+/Eo+7hPUyYnucg8Xe9E6edP1qUa3TH427SsAhTp+sTzw6ATm/iZqCUMb7moHZskA4W8
hEnvJUotep0QdY4OUT9Gs0m1E/tKg6JZcrSz2lT0E+KC322mAPESAkKlSDFgnR3q4e1ZBkMuQzRa
OVma7IxQS/44kEgfSXSt51x4P6QLW0muj8qlPnt+E5Z7BwRXnNUhw/BSZ1aSfln59ZRwNvPM1LHk
1yzJXds2F54yH6gHVBBbZVq39ctm8o7AQSkfbWLlveAeqjtQHU9YF5McTYJNKJg2/CyQrHNKaTFN
ItpZkYNDIegYBur43q6JMDvVMOyHSdBx4+jTytnMVCsgLrwzmwYoqIADb2MoF/eaBOTZ1fB6FvC7
J0K+L7lq/Fztfo5yN7HFxPHezhPVLtuqju2P9P+VGonhDuH5m+A9gyrniFNPGU2Ex41gIP7E3JLk
hn60NH1OZLtRfeUsjV7XMf089iITFnjKSEC50uCDEeZlJtqmG0VqNdnUE5Sat30RHzIwp8dqqfdO
BHWnlenC+AFxf9HzzAQR1dhflf8WZXxKBhRkkYgeqEoQkGGLPMEcuaeopnapCm0KwU+puUZgIxW+
M2rLqh5WnjjGWSgsPnUWMUFzfiGeTeMc8Xe8yw1JZCbnUok4S3Emp1momurTJU9ZvGNHHFeqraaH
/D0tC/6g0nDeZQpG4NaYSucgC2haeajmuqxdwqxLT6mA6wbMPxN12m8YowUN5J1aeVc2PHa2voA/
qdipEx4WPO6DTVlEm4hBYD/WlLKnHnju14pPuL7kaIFHC6C9IGXxvOy5asv0WBCvTjvD70rBaNDw
VX9tSIGrWBWW+JweNztobF4h9Fvex7vmRTPuW7rW35KQ7+LciOdf/dkm0lm9ffyES4v0JTBY8qyR
KZOaRS95+hhcn8xewJFdcW8hPg17Yo3sp80MyBWzQO/73e0/JkDrE7LtS+HMpE3hZbdEHRagc/f2
DLJ7fZZ/4UdWk4H5kKvyI/fpFyq6Kcw86SUSvR1EliyCafE6ZzO0Vd5zzi/t0dUDKiIGeoQUdUlg
2RU9LVvfCBpcuiT6VheJ2l8e8BJzC4GxVC0HnTggYfiHOfN2OP5anm9ej7VgAc7QL0Vn10IB0wi6
tw7EPaBzHrnykbFzD0qZr5CNYIOyoQtWVOdK0ST+S8lnVxOAf/0PqSrCyffJnFdAWkQzZbHxQeNJ
oyJU9GkhOCiJzFJgd9lVsoKTUoL0dEl6zZ4gTyNwwG9RqbeHrw9cDdYOAvNEb64YxPMdJU+zayUa
iPpgcZUepIQSdpSVmpZkXr8CQzBsc9hNgi/VPIU27wu9gI09yhwgPz6zXi/yyQXuu323yK3ogf9z
GMEDW9gysNeh3bVRSOCeQC+9suQO/S8VLrt4fv9EF/O7kUikmxb3txqOLf9Vd/QIDT8gdGBCiN8q
1XcU5+v3/X6lwYL580zvnEQvTByY4HYlun+68wUzukRCLMHG1MKX9QSLQ8gDaXazwCbrvvnGaPdA
m+SFsf9PGqbWcBm9OVEkOXme8ZFm9bUhncFllYK6Eyo/opux1PpfqcHtKa1BBSVimwoPatnUp/Ts
RNl71V6IT7d82LNpO1VrFmUGx/lz/WhsNBqdb52qE71FyVJTCIcjwwUCt376Aee8j9l75jSQewTF
lSiGfXFINrZ9UliUjMwTWipx0ZwzUHL0AUl9WkL2bPbu2+MkELp8ahE3aA482RXGZrMiaj9eqLWT
H1sydB5wSI9wARWJXWCJVHaMzZKCCxlzRggTd/cu0uWuQ0O/Y5gFeESw0Q3ZrQWG4LrpwLleMT/6
f1OyZcBhsqJtO3SvrUrDar9xcP6Vd134siK8ZyBQ7r+XrYgAVAe1d3QkrOW/nh/mvqWdfdwn+/Tt
XUrzIBC2TI/OQc/4GU+LfrGaAas6D2cBehZ2YCz4BCE/W9q+zCGnP9WDYBhJ3ghSg+8nbPfP0noj
qvpOfK8HWwSA5Gx2RKpGsQwMvCHhCSsgbiGAWmoqNsrqXK8H5+MJSrJ7JDf3Cl/eEMbWCUMGdFZl
E8Op5tprP8i56tybrmHkWdnsBdtSw/Yk5cZn0ZWhcB5WHm6KT0ibvAx5uyUY0OR7BZZWPCHrRovV
r7hmirEs5Ymr2CjRmZ1SkLdysIqsTPoNS0Uf0gSIQIWcsMJTcLMgBtKPG2FeqzpQHicWqZlGG00F
8fMs/r9voVLP5A7vukSuYctSDSti7SRC12gqAFtS/8L88kKBDwbftDrU7Cwls28fbzXhLx3ZAJAy
LxhvWo6yKqyZ2iXcOXouJ5Hgj6YjozUGTWhLULlQFh66pKnaw6uGy4+PBh0nSxt/y2q4xplB0XRc
jA1pGsROX8Z58WYYdltxm5oIaSTBMvA2sOsUH9haI21WS8DYCnYNYV458HspB+v77916CoLtNy7C
a3Yh7fp2GlEuORTkTts88Y9XSFCMVoUKsKYRbFYdSMm/12aGzCiAMBHIrnwg8FLQG1CUcYAXzV2x
1CH3O+QclR4nK9agjRAKtxlG96XLVpLxB+hQ3xwhu7c+NQ/tPoaFimw5/07yyQGiCx9hhOnIq3sq
nMgPg3WdWfTDheLpVFdvC4uSjQOyqKHbZ0Qgde2gR7yo6E8wtMxFs4Q26Bgd1YJVHm6h85E6xSo1
+x+OwF3uL1IAlsMwe+PK9Y1FYw8RVhwgMA7lNu8kmYqh5ONUYvoRzfpNxEXNCYpK/QnP5+Yhc256
wEVydB2K38V+ff0KBDv7V1IyE1P7Yj9iiGu7LcVj7FshxAXwvfIduTmDOrY8TvcMNuuZZMJR4xAb
1JXhfdAYHkcNQcHbze1w60WGdPz2BXixZCtMVCwVkgO3Ky4U+VTTWc/XIQwYou1Mo8ECkWs8FHNM
GDvtERCUSc/yq6ScZSRuRgWPGEpaGe2wXbTKZ7ugyg5GbaInn/kRdFiHQzItfgx5aRhCKeispYku
5YzxyseZpQbXNjMxdLF3joFOB3c1NqK6fTsyi/2F32lULqozegm5P60oR8PJrHdHyq4vt914Z7VA
r0XJ6tyLu8TGXGDMyDo7d1OOB+6AZJyKDcndoxDUF7p6xQuvQkClUlUpl9hzwK0Q41tSqT8iXJlg
wwrmAvBaozGM0ctYrG6/2hqYBFMaMlnkvyDai2/biiUYX98NQoI8KGsOzkWJMmaWRd9xff4uy4y6
V8omg+9fq8wbdlJVvt2N2/PCPYxJ+rMTDoPgErHHVllsyZ6AgS8vRi/XBc3kcN5ucmJmlRC+tTwi
TyafZq60XzJFFBZwPmASsTLXfE3vVoPEDAFTflwN0/wWLwRfIlFYa2SVTt+MG7nAmWpdP5cExeQ+
wCsNaiOvBlC15gZrHBZhrlTu46ezdKIyDAdve6XIMVui6skJ+E451tBD4/9r8MnkEbqMJD+PQ3nQ
9N+bL5uYNFi0ctHWClGCQKYruUPeH2oUntyWlOYIsVciO+T7Fmt40QzvnDl7hcGfuQ15rmemAuE0
vHgUO7drVT9nGdSowrQrc5z2wIvAL6iCVUan2DElvlZeUOG+YxzNukZ0DM2BBEDeSRi2TB5AlDPC
s9tZekxalB0yeqqr61/1EXMJU3iu27XRllu8qCHiOt0b9xY5uPkjMxtfCPxfLB7jrM7a33xV2mD7
aZ8Pf4CSWJs121EtCCxZl9SLc1CSPFnjsHkQPiRNsGUqmRCJ7BGcPxLK8QvQ5GALHXfdvRe7Pjhs
ce5MzEaQOQ+L128mgCmPjCjUHxWPr/ogUignScThIUOY3GdQySe7VID7MMyG++GL0iUbh67cS+HL
ZoxIDC7GWP2jBWM2diCEI5ypz09/YPdVd9PJWLq3tzLIpyiVnSFAFN/fiTolRWVk5PiMeSXjBilm
ca5aeF+KpVyl3h50xOg3A83cWljZEblzUdDyWjq/Bjb/xZOB/vZ4BAPZJT/eq3tqaLBd774bSdrb
NrWOjNzgpxNk0ohsqWO0zm4XoXwQKcfrI60YuoWerHM7ZJqXOdkQr+wFMLPv49QJyXH+To+U9MX1
P1uTVGX2fJ4CcVFnzX9exCkuPqbMWzOPJvl/gf/4nR5km4cU073GfmdMerFK50Niq5ujiemK9pJK
GHY00j9Fu/m9Qw6U5q0g5YPNqhn+kjYzQgtmI9Tu0B6leHiPjRKOHOuXEAW2KT4cRUXJa3IRwo9Y
QUEIyzkd7MultLH7+u8D2ZNh7GsMGWbTpeVjlVmeUkUdtkTUd3G7qjIHCbaWfJHWqUF2j+3RacNO
vfiAEjcKKmF3cbqM9EZ+luomJ2Kkyw/jyjP19uF9E5jSLHUS7NZwAsmh3UBPT7bugGLsAZIeGiEX
Awq0YfiHBmiPSDr2ExXdbF2ePjhqh2XaWELhERhMXFgMAGvvGZA+Ect5d35/EFxbX/3iC/trRWvv
v+WjMH+u7UlTiXBjGPc66OgkDZ8PrLKEw9CdYQM/4NqEqWb/lHEWRodBlNZgov7yK9gSi3IJet9g
aMdn8Um9QH1fln4jwVsS1NNy/b81OIowsnJ50WhjQRUJml4FGWxu94wriQs7+r9vlIUgloTkHZNc
QI829/9/lTdZhQo/3ZzE/AZACp/IJxynBC5wXqEzqtKM3yF0f5UIpscGUKg/P+llXHHjcJ6vLjnv
axDZKyStapkaVA5B4N5Nhj6I7mRifpC45Q0Wu4qqmXlcQmgHPwww0Zap7dLZPMFHKXb+MRSh1k4z
ujWsWHNYV0lbYVCvUeTQZq0YuwzA62y2y6QHkbiD8RzzEL61HbbQgvwGLulcx4smNebDiGaI36Ln
1V4TrSg85+iCwYlAMBuRk0pQmuYUWdDCqWicjOshalUbHP56nV2Jz8qCrUBVHwzE5Ni1tOZB3H+A
Pqu8cQ/3QiU2LK1oB295z8AnfxM6TAbl2H1dqATQ1+F7Q1E9oYnd3agGm4mEpfaeceWUercs/26H
Cfi6jxb2xljuCE2TfOUThszJIXuO0XnqyVqjPGrEtfeuST8IAr/YLrx3G2UXAy9nTcmbZ7QGLvqt
nuoZCDmb6x2mQShcHus8/cG9lUdVkbmWCQ+7nrzUbbYIqnR9G2XeMC4tAXTaNA7O54kwCWgNINsi
uFowhtpzTq6wRs50vH2Hq7Aq04ItfmJTwV34Z5i/2f9M7JQgQloJNLZeqrAgJrRj1say3fcFkvEi
yp6m7e6iUy4gXMrzw/UJYqGRrQ5FyBqvWuQrHGHvXCF+QH7qfaoZaWBf53UQCsUxnMWrgNMQu52x
wyPMA4cVb5CQHbivXP1DFisU3G5gGyNeOtTuWD+MXhvXQYCMkBbY7e2Wh8PsWRfiD5RV9DQFP6wb
btB1hj94mSIfip2wNsCaj7RU0T+FjUgKNsmbNqiq/uB3qq2Xkr6ZpBx7PYsndTl5gUWLuXYvHP6l
Zj+z6r0M6Jx6pgpHukbRz28/5MaD1O1RHXE8JV9+Zp/IuSABpGH1aO59jCPXbCo12IC22dP+ssgR
xDbA4YSivpD7HwTkOEHdC4GzY+r3jZbM4UbFT4sLoMK5OwBtaev1ZISh/oGgX2QxghtkN9hL+2t3
DU0HYXqLY5xxB3vj606Ez4aXCHSFT+ZdIf4kpx9PfcRKivIpQKrjFc0Ocibqn84Y3qnpxgWnlswa
qWjjRfkB3b2zHUNTSZ+LPhKagGjWNWL8KnMzELzcg9pCXELswdNuOzKav+c95cPTdLzqW1CpS/sh
Dg924euKbjHboE+wzGCcpdUbkQzr4X8KVml7cdCtWOe3Ne0whHyEktE9m/E69NRulUfPcvsRji4f
yAvyR8dIp0DgA2qZ4nzTuCLQl2wrs8Pzfe60t4jyDCixrSjMPqWkNZYVMSGkWZj+7LMq6aEebL2m
C3EoSaonlihIj0P6O8vJjxfOphzSuzUDcdR3KT4B8iWJH51U55Mxa7IoMwQdzOofVbPWzlw/QzGU
O9EwtAs/sTNWckvsLlP1K+OajnecefhC9ECHcVKoJmkWk8b700XInUB8Wo3vIXqgJ/2kolism4mp
y7ynswHC9CnX/Gra+9YVgJBAC6RvjMr7mfYzxviXAHG81jC/zgEfi9m7ujMsXLN7pUu6OapkZRgy
pUniZuVE98lolYeqMCAUaR1FY6Mo6ZH4yy3YCfZQaTDsyfDMSbJCFXIPPYQb263oHb+rho81SF8F
LGzughX5JjdBT16OvsFALSdVJP3tP75LkdDhPmrdD/xwxRs4TmM0XXC2sShdBMcs4dgS8kpXVk1x
NhdjIS5h4HK6yy4BqoPtpbLkg45y8QXDZot/sq+cVFt3L/Axme82HRoruvUvHSfPnpzSut4hILjt
PAUqbmhUDtAoeLce59rpsem3N2yQZcWAig+kpo3Q2Z+Zr3WFfgyROEH5Mxv8hsBX9+AgZ2qoFU80
I9phRy6EoypcEIQj5CH0nD/tyw0KwgWl9NU45Yf6l40Y+trwaQEITy20JN4M/uIW9q3/mRIGu0zc
b3NvxZGBQPdFQR4O1zOWxQtSJk+V20TwY2TXgwYMyrWwG9CcI/pUgRTYNarAEMaIQTAQOJZoKOSO
jd4MKaMtfiL0GUSX33J2BvHMrpUE5LZRolH1H5ZUDiSL2/rCzV8Ikt+v/N69EZNzfXRaYxXL+nVY
Mq/gqs9KQz9jWyJQH9vdWh8X2bvu1W67XfXagJ9AhIea100VRlnqjzk6f9R8vy5GoizFnwZNYhmS
uJ5GoWKSwilj0svh1EojEOOj4OcMPkAk16oRUKgmBbKUiRbTirNJT5FjdyQXDzkLZOWrHt8Sbg8s
zEWYzaLL4uADVjQUPH/eEJIaDyfUzeTdLAUStrhwGTMYxVci94kVvmM5sI2THxuZpofjndUxzc71
c04edkvD+4owIz8tPKSk7pgOWbOR+akjVw171FEujKfZTp1ZUJKqTzyL3BSaAorpDuND3dAK5AG7
7+LvtbnEoi8N3ylqTLoCpLjxL5S6SJztMEWZq5dhnO+aC+u4JhXaDElUA71Uop+peXZ4s4QSPyKz
fR7fOt+McD9PsWkr/3ISA2DAXxjeqAR0Tw8DqGYBfE/ViA3/Aey+p/d4NE3rrDQWal+MWoL/rDNj
8M2dxe37aMB6iVSRhtDvSpg546yHTAqblKzalNr+Yi01MWD/Bv3ld16tPVqTuKe4LxG5GApMs0gV
+9ipFowjM6gDHP0qG2AB/FDYYlkAKfUcnexzEYvtQ8k6D7P5L136czjYqcszH5PALVZcaAlAOp9h
20++/hj59TRnY+3JF38zCxbvx5nldrX70TRXWqT6KoY/o+YjrCBWR9wFxe/7JF6rNUkAIGeCZFA2
JM+CyiRRY9CYmlNpA+d8L1TG+XdSteaDc6xdh0qJbyg0Uo7XUT/mxGgeMD8TJX9UMCzueQAiXg0n
f9ptuA3653BPhAdAyWLMV7Fw+yT4zWjzqrAo4Oor/H9HJcIQUS7AxEBC4DDvjwrOSO/CzkPBRUgD
Sn2plJGTXC3W31lNkYPRKZFs8Y8E35DlmEyxEma2ldHJzkPQGPmTaXhs8hgjrkkRJPbvJ6xvQK8/
WC8bSTZWmZMO2usvhKCVT8CV6fZvwb/dRhQmT/rHcarsA8fxZZfOKXO+cnEpBQwvg+IzseiCzjo5
MYDmarpoPmUc85qE5WMh2u144DGl+rJjbQfX1hZUZajmCF4as3aVlh1DM62oJmcCCfdD+Kp1bYbA
ycRp1QN5dytnFrusUxEoYtxKfC2vadYt2FkdbtnDgJtidb0HjDdXGyrXn5MH4nd2jdHmEhFOMP7O
fmeOAxKWDVtt/7PFZ3jwfFt3jlM7P9aqqiWCPjADl6emHMN7AjusjPcu1BQ39AMM8vOpPROd+YA/
xdXvvvLd+0So5LPe6w+OebTvJ0gbXYoOLCSbDb3ALzj/27/iiAwvewVHbZ9YOWz3CkMqULf4b2Bu
zCsjX6h8qt5TapEzXxoxpa5hEVd1ejc9x/gsq4cRlKb5TkLjjF8Vc+gf4I3ohGwlpYDlDGoTmFpw
c+B3GJD5mWK+ecEmTvZZ+egLvwi+zTIYKzRc1hUOkXOqiQ3ieTOfxnc1cF99Wr0p8w4XUnp2tQ0s
wsp8INWlYnVre8gtBeM9wXNb+O9StXSUyvkJ8tdu7OTwNr0bOI8bP12vqsXCFpLMPVP/U3F2Gvit
D7hlhNyK1WkBuMOdklc2W2eVQdtRIp/QK8zzu+cKXYFLsNpPHh7K9zcsf+myPEmYqAbBMTIN3IEv
ljTyBfc8a3wY4m4S3dCtPAw0a1z1zK5wo6kHmXxv8OUiaXX+hTb6dFEr+KH9RGeysyBbae82v8s5
lQvBqo/CY4hsNL3NIa52o2pXaJ4k/kphpcE47DAIrwRdHDEj7nc3nNl7hdbqZ/2F7WnTKIjJWhav
ouuHi0MC2DhLekJjce7qDSb6CiawK34DIDXHhNoyIc42m1VdN2mbRYjFLcnGY//vJf+5e3re++WV
B2LLT1mWtsOLLtkJ8Yc1ahmvQWPArU8tornT2BtD7iiBXVAAKLB1wDoh3pdeyTwJxsxmW56uPsKj
jQgfIia5h+RBzKT06et6KrZyWygB1tCrHZoRs1ku51Et/Mi7NfPHuTeLOW3qWE4eIjIgSv2s97Re
pFpZzHc96pvJsMNYQTmLb1N6MSvnvjnh8rOrLo7A0Y25jJxALOp0YITSkdGfx16C/KnberVSDVlp
Pi4hLMIGhCMHAyasJVSWZX3pP49Xol1iju4mpsOL81gn4yET5YbQn1YktbroPkgyY/Rul/qKjnAK
GRS89F6xauJesBNmSTdbYUWQI4LG0mbbDUSHhiHfEuPnWNxReg+5UEbeBMfwyBZxC5G3ZnT/zbFX
w+wo4mzm5+OlYc0nvdU0mb/HQG6YQRVm7nsa2SDzTiNa1rf3E2yNgXMMD+FZbxevrl0fIqkdE9Ng
EYR6/EO2nTBU1+U3ED//BZpSS6YV64goupC9s3lMpHnLl5YY3u8Jk/b4Q7vkiy7YRE+0dqY4u5Vu
LIH3K5YRptOZ2CNek2GcNgYShRXZhCF6IswtD/HUkOmBFrQMHDLpciBh93e5J5ao39/LySC2IJ0C
CuFce1Xxzl2KDUYaHGNf08XRAWIA356mXO+yI5TQwvAIpUNavfFgyJy4jzRBMi/Yzgjioc8tYD99
jwbtujoYXiE3yD647aJCOJDADtEjW6j5MrdG/nSmC3nEoYQXfwdeE9v4FipZjlQ0BTOVb/Dytmzc
Lf2y/XyfzxSLlWqwK9trUhLWmEphNVM7gJe+1LsdUBZFPPuJZLtE/livBOn+mt0EIp/rra4WXDAS
pySWSIjniOcmhvWuRAzAcFG1+HfGmpxJrw0d7n4bkKus6SmOu4/xA91fLx63ONlSobCryx1b7OWI
Awti4iIBXqLTtFaF29hDHgEPf9qosXHZzEHImfLVuRZoNKqIlOAJ5qGyybU1UW07EmDcQxSbhgKF
J0dmGyLAtPmQ2M6mP3w5tvCuJ3RnlKwYLx5cwl02Y75JuozM5uz3XaQWflimgyjPoSsRRvwJSkHB
dqAPjn8LhckqsaJW7LSn0Im0sXyMYL05NwBcXA/npBEztcyuKGAZUmH3OAujyDOMz8kgsxYgHSGJ
4L+p57wWYof4URwDUbcpxSZ2NnUTXVLGeO8t6+Rsvb3r0P5a2rSLtU2u2r0KDu/b4E0KYeU/1Yp5
aPlbyYsesshkMPScs6ymgJvcESPYSPTS9HLxOXQhmFYiO2nHbOVXVsTsc94hx/I765s8dd0kKu8y
2sYN8Xfl04+zWVE+Rrwre3k2COvS7UHcH4v6nxrJZ68gPChDLu3lprv+fGrP+dtElCIWkL226XAG
J0uVVRBiyHEICF/d9mQ3vN61nuG1DiPSfDrE4jbTP878o0DQxbJ030aIXKZ4LjqsMjf1/CGeU//C
NqdL02qak9qOUqGaDy4qcrzKX0wnKeBYDDsKII0o4DXYwsUGAh9Fq5+gOfSrI2LRL15tKqsD4W6E
EGdZL+FrGQuWmlstyyHABCvdHH6oD23elqzF6NTAlQrmUStLMCMNu1V2B4wCcQTtejpWTC3uHs3s
6QslrGDSakxFS6as3UUf+H8ap4Kl/TPo93oVrIcQ6SYPpYO9WhuP+GvpIRzEvu9R1Qe8D5DghryJ
P8p+Onen3MbM8xGDchk8yIzHAvi/0XbWQ4dzaE2tER03/jwtDZ74gdncZxdxd/imzqms6wRTyxf8
Hvhvo81UbWQkBWCKEhUrlgvQdHVd4oA/u8PEZ420shiuHuFXh5JdTXTdg3zqWOaJGjviZ+0XDx7W
w8Cyv654yRN+8D1yGX6xD1epZ+l8SCyVXrvUqeTNHhGbT9FPD1dDl4EqN1dh+ZL4x7oIvOiEZIno
N6wCKlE9BLVzvU3XfzITawF4E2em/SjrHE9zT+UPjxI8KNViEZyirdG6uOt365zsZD7cj44zgWC6
cWPyEBQc5qfbfxr1QgZYTAH068YaihgEjpqqJz336Wrr7Y5/tz8cEfbYmvZWX3N/wh+94P+lHI/V
80LGy+bgCbsIlQHAJWwUs5fJJmgduVvoJ+GOT4/MaPBMRgllUnPU53J+Pcm41e1HPmCMQ4lw1R/P
wQp+TNsZ+SFRs/qjyQhLlTOe/YRuyLv2OcuP50OY2UbN9hriVmI4vtu4FY+/OCF9y37ZmWIp9zjn
6nu+TNoZ4pLc/Ql5+iBmjRJ0vx/0eNUvJ0jKx8RHRpkxlUO5M5BTvMwr6tN63eG4JM5qU9pudiBG
gwjhGBq/svCUsbjOiODI/YDhk4N/TyX4G1hjwVUqR60npYksHx9oK5+D0MBZc0y7CpFeRcEm1Cjv
31Orye2wzMCYfP5veUqYOPzzuAXEVMHz7S25ltcIau95xmVPVwhWFKt3zSn0g3un56g55drXHAUl
lCz4Hdf7nCdrdIy8o2aF+sLVViNQL6zq7EZBfbJhtwTYiyIEI7hJYtVMuIUdD8SLNK5JQjEwgTyH
yjc8/AmR+8DOr5VW24sCOrr8l/+o1NZh8ZL7iBX0sqE7BPCyD9yJckm8KNofw5singvLj+WSSF15
PRvAoVFLL1Boo6dk3ZHOFrlrZvZwliiSthqq3WVY1k/a/fTIQAi1+az1F8L8VUk5SzvXSVw2ZMeR
76TlG4gESSJZpflIpcT52622l9WZK5igjo/pdn4Fe/LNaqbpAGWc63QIKNuzLHrPKN7oLlY9eSwq
9AiMw+anWUoPlcuLikWfzuUZVHZL2rDDG6hOxqDfocjBd7HKZvr7mcK5uZqAmovwWvduyQIdoC2L
JHWL801pjEuvFJ6EfVAcPuSoYEryzFz35RKuLlFOOiuHn6dh7SOvGwUV2nbjYyzIzh/zFr6Mk8zj
031lD8paYYxcAUl6gfFeRSB6VbeHFXD4bTb4jIjpXOJbKitA31vLH4nPNYTTorSd28o9GXAaGBSY
5drPtax1DGdBF63r2AzpiG4tv5ehifQ6HbR2oKE9eoWZHyyrwmDvyF+tvH2ovEZzsj6WiOL2dtuG
X66gUukY+pirXs6craQHLVSeco5DUUGgSMa+cs7jOjCzzYgXpem6MVezyiNdM0rnr0E04hhnCu0g
hmbzgKKQz97SQQuoYVzr6yM/g5vad6uFZrEApmEiWJ7j6iTqfeRaYp2E8SdGYIjdREolOKrBkggX
bbQX84qlEOUVsvfexdH2HhqRwHQQ9gzXj76cuVwa8C0KxDlRL8xkSJS7JlaSthhRmHz6zgg9+BBH
m5yR96ABVEOpFMiR6VzXzZaE4tyhZpL587MMikTd+quDsCW0C4ieOqd01q9ZJlhAyw/2fL1Fr6yZ
hc2sf0oyG2WlKLKLit67M4+A0KjiZHUK39dTRhLMXq+I616JJI1uvi/fv0exQtgWqI1igJ+sHPds
PNhXsbkzJR53I5P/ago1nASQXfsOeGIqYdTrcfTtGIw1Z5NX4cy2TPA5NcYteCpNE+URWxhjId/U
HDWigp3uVPVbJh7/lihVq0n6pUOyGsKc4huwRj/46TRSixJHP6qK7v5fC3GZcLfqibty+gA5hHas
xU+hhevJ5E4xrK8FiJNjVxp8mJjO/vsA2GC+ptS0laTtZpHyEFCBhdXjD4kQob2kvzjSsfCxfdif
KZnRY+xecdmaDvrhLoc+UQFhSi0meBBzzmTGLKxkiO41BSJYDY+pqvKA5FPMryzQziMKHM7Z54Lx
v+K/VU98y2jSGUtvWi1EWSYuKpE1VR8485iuJHaWaZBfq4BvzMBnvGkfq0SlwS5m0TpN+JNAySiX
GcwG60Jp2aBXsph+iyJYYOa1YzBoMppIcD3mSCBkt7fABIgIUqiBkwfyNFrw38PoB9Ty351QuFED
pKuyIj5+IH1uO/ZR/E7Mano0ObhpSFMCzN/wIT1/SMSdifqrZMtpRUWclWI8dICmdsCN39vr2USJ
CtAJP0LE9juxPzQjO4DW59iV/M3wnst8bIgL44MV3Jw4UdMnBertXmqvRJ50z6+sAfAnLQY8KN7h
HcAjkD72bG2MUFTuzoImY44mh/hdCKC/5qPyew+XgF9QkXurDq0IjpRDUP+AFHiMLB6Mr+xbrMGz
F7lkByu/rEe0XcKoBAiJq/mG0/I5ebAOa4SmtOLsVfwKeHgROx79m337rDhbyHdmju1xSCmE2neX
XuyfiOsI71ULIjMXpDyrttfuRu/pJvwSqTSHUFVC5D6QX1vCyNLYE1krSfLiyNIiVuKSzjDk88nV
2ScL9NY2kyTAq4EuMaWqQ3f+7u2wSZ5zL7Nb/p34MjkDuWwU+aKLn9JrAjrZAGUuvOdLQlMR+dDI
ky6UZTMx2//3cp2UDSmZ0d0rVEfchv8R/TRZiVrtVl6iZGPbyrcAIu6TnTsDhy/ZQPetVmq8A054
xn+DabcW/Hq1LC+uRcW+0+FG9BKFFjiGpdXEvkEfmxpAZfc4sdlSZCOEpzDynB7YLIR0ubRanVe3
1OW8yXVaR4ICyPbY5Hnmq1+xSkaRBDa9Fotc+zJCcZipFoto7DRtHc4YnAV4hN4A55P86Hw6F7AB
Xf5iVQtz9JeI8F0KH9oiR+U6mNZYinf8AYSuBi1Y7hpZu34lfymFgys2yuR6XSVj9lzoGSxqx+ii
bjgT6NssPoOkYC0OgpkW3mxr9W1LiqZsy3s6qUkqb68vLz9D6VAAzL80HV793HPpipHg1SGciO3S
8y19hjhmx/26zSVv/y/HQv/VfMSbFG3WZKC+xK8O2v0GrbYhI9UyTam73JgCHD78KH1Fs4me4PNV
oU7dqJ6d8oh2MmbdYOLjUBh7IhejbqKaHmqPZRPo3I4BL3c6sT+w0qLMxWJPJoOfOAIKiVQbfYeQ
CS04mguYW2kGJpLi3HPkr/5L+eiEN12VeorCnKwkXW4Em3YxzqCzOSRJOGBBRnJ4XcmZUoBfR+z2
k4FF16b6k825mwGGrUmm/xUfN9SuIxEzrHQRJNb1l7SzUY5lLK8k437lnY2jvKAlWwn5KfuMjlTv
HWghQqqPQfGqD7OyvALEK/L5VDZ40VKgut5/FugulzNC6qJnA81A14jKxe554LCHga3jcCy+TjK9
za6PHBgUBko2elF76LRnIM2SFbfDuWyZUWFCDpDTN4G0k/Bl9SE9aq30waJRO1fj9SViBtoeVOtG
OHCsIoagC4+E6HwOsXYk6v5ufccpK1dfE/WJ3MIbkbX67zFD2lNAKzMLgCFiS1A3yWEqW3Fau/I2
1oS0rKUfG3SaCczEzKBIguVwN5r8j/19vzFsIVGe4ULGrD9cIq28yASYwQpUHPXcm1zM3Y9ExAGd
u2y1Bn+V6jzi0oNKhz8Dw0bMLUZu5NC+nVnout1Y21cavT7/H/UpFPpnMJG/RQOp1bUZZ0PORNdy
oN9lqdrWwOy5CR/P64w3T/18bmrG0bvRS1Fe7SH28osUF99vIrlh7Gwm/La7Hmq80+EeQDAMeFwb
sOZnsnt52ZV3qNWnD+rhhcZNtpzvP/eEGWPNCXbfwvZGEsTnnmR3ZaI2HCsP2QGZZzfgHg2l/Kys
TSgVenuQCUA5M5obaDynnsgWOZRnWSyWHVR0q7Yp2O48srT7NsA3WzpARD+r6/AOYSntGJosC3i3
15ERs+Cjr3PoPmgaDT2S4/HAid4deSRojjyOWtudaLtz6zQsQUNJqEG+GCg/aaYcfOvB59pO24MI
E4hDn6RFwlMYO/5k5PBT0iaqwsv9z6kQJHX6hAAcZrv3wFu9pwsu55BLT/A5zktdUi6DUoPIqA2A
InItaRy+7KD+14/QQjtQ1RB3zqnWxMlc8eugAaF7L1LcJz0gZXZSrlnWFjFjRCDjAEmAIFk7pimZ
Mfkr4s10CwxDGXatwAuqcVWzsGYwPZWIfOK71bwgLnAm3bgySGAhQel2k10x3zf/xgYIP3LvLt2O
Hp3ZtC9KM3EsavDCrA9zTsRclclfw9jwgPDQfas6pHsXEBh9Hm0PPitNRzWiBWC5HKw2tj9ssuoh
Vwb48W+KJkJbj+KLrgvLSL/3LxNDSm0+aIeCar57bXfIxTFL8IHdNFg2JzLTJpVZ7VL2rAbm2MJT
AC+1WVGAT0DRxt266QppZ3aVlMKzEdaoE72NiIXhfcBC8k0i/7CKFWLqxvd8XKyTqNj+Ky5WXuaT
5aM/AKCC4C/e8XXKu2fseM2t8c8uBTUahbBtR+g29bM8vmiDOpUNf+tv3Q4LeW646Kpx2Fh3uGOu
KVT8p+DR9nuq6khJEDYrYWAAbHGEPdh3ee2u/IS+3HETKBVDQ5LtQxhD5Jl38FAym7tbtBhF9oul
aLCGWdvACKiBxSWzhKQpgu32rt89Pw9nuiNxY5uKfLfZKyZd/UhcG/BSdyfrHv6vSdZVVtTtovNt
BJ9xpmG5Ym6RH5irRjvIo3Mt4S1FRr7l9Gq0VP6cEiihoKIMcAIh0NX0uqP8Yfh9IPkGDXCl3gUR
N/zxlT6Vk+NzwSsVslDpkujEQsZ8ElKAEQAgjg3QUBMpdV3ziqHQDZFHbe+gOyC2A100ct4BQMTH
NchSbsavlZbT6pbYOYcBHH5tgSLiDeVw8d5m5GFkmEwYCEVLhEF+eavF5vwQziEn1U0be1fywKFf
ZnrxUE2sTP2WXvnJ9eew4bEmtQTOvix4JQOpvFpsI2+5rJ9Su1vXHO0l2rVgtFrof+bsP7Ei9h5c
SXyWNvGmh7C1kuDZ06xrFQZajJQb0a4hyiZJGOa625ukeq6s0YpniVECcdmE/5y4lY9TUbkp8j2H
XSBC8mUrCsG10/nUE/xBH30rC37jFrIGlLEoF7kJ1q6av5HXnw67pDAf+3m4O6s47ETqaBzJFXMj
fxR0OOpDiWNEmhrL6B73ITGGdutPdq1OQ0xuneBVH7z3PNgCClsgIzlJXANaOMOXE0rm+Kj4Tbhx
DK8qTC+voUzxsSr1He74a+D5cA8cLWoBR+nvwg4f1LPBHkqLZRKTi77ftuz3dmx5tZoQ7zMrPrTp
UyYOBpTMvkw/eK011m0Y63dOwhzxb1qQP1d0zZJe8j3tMouNXgI61UmbO0C5YTnNU+qPPWvOdTg4
fCtQeZJXNDEF+EQY4X6/K2j+JkGfYJbrpLZGd0i2PrjrSgZKcmhEzSsOW1DBYFH8LAAeYtrX3Krw
69ubQVeyqqiUgEM87D4C2TnURvZJD5Cslo/nPh24WKrr1o8kZd0lKqT6f7fi/bUVBwT3UHQqwhQ+
FTCqkJG+Jt/TMZVzKo3BxDTFZTlh9Y/ZjIIdw1sr4xMMliWguLSuk7yn8kXYs6DAl8EzoL4sQs+f
UgyKCiwvanUB1xCWoarS3Ns/HcDkpoh9A7Yzoqa5gutR6Y+V1hi4tPQ4sYVW0H6L8dMeM4/akImt
oNklodoBR8R0maNhlSmzqRxGyK+MY8yi3778rhpPX3GmBQI4S6rShWhPJRuDPpY6AHwukbMeszqF
lUL/9QyUmsSSWTnhGXNDuwjHcf4RgJwVxWkLutuRMXloNmpbqLEFroY0o3sydwTQUcr8Qg+B9I4J
fWekPGOyFSEzuxAmV8EPmun4/cY+pQN3x0vMptL+fwvFRMdgEStNbHQNPcR7nmal7C/gXXFCFPF6
ycXl50HLBF9KaBHORZoxhxeIgky4MVD9bxBle7O67/kt/LTyMaGXclFqGhgvvbOA69R+WjW7jCwj
pfY1k2TLcOvMK61Sw9Uoe6iF+p515DflKOagGJzW12eKw+1+pLQwQSdlVS1h8ji6z8OkZ7xUAUOP
uEsVYpLDlfOSJjNHzmm7TtVjUeRXKD0QCWG55P7hxY/I1KwxngJ7/I3FYuYTFZ4MosTWejnDDhp4
rji0+JxJi7h0g9rNrQruuGMTSZ8Rj3Mi/06/eWbMOwHUeFh/d7JHlf+msiqM2dA5r3oMhD99IEJ7
LvLI4eqhAPYoIV2Q9d6xsjV9GoxSUmTHbCW7Z/Bhst6YCRr4t9Tfg0b0i9yLJr4Ly1ECv/UXXRkc
hWqecPmQw0NXmyxXc0IyR5zsgsQM0TkVzPtrDFzqKvIb7qUGXo850v/lXi+4fdfAEEXuFmCUsN70
nxWDc6RWJoGJfm7ZfU1+hoP05qUOViyZFq+VZ0okjrp4JeFPzgDVB6RFEF+NYMcwUWRdPs+EIE9W
Qqx8S4T0zyC7lEHg/XLlSyv3rG7uMkkVi+oeCGJOmiK1P4PVOYN4VWcuAosZXC5RxSQdFtB9GIFd
v86fEz2ZEZLCVnaBH8Z3rlxoqTIGXA4R5RqxlSFZxfpFT+srzZAJ4OxrG25DVYn4C3IVY0Hl1kVZ
pSTV1WEqATU0xa1lhOU9GVApF4uRLfF196u6qB4thah10MgjtKyWapVLCk6OfuujpRCBngY6MNYY
CaOp/tL2E3mpL/swem59u14QYXuwck36cGJxQPu8/Pq+vVHsspF+rsYJZAzqNkM1xv1Ib/aOXgJY
P1VCz5Q2uhGbh7cp/AXUCwz6hljSYgox4diCJTJb8O7NgTlKnAzV4BhcQSXbb8/++I7Lx1yxGYuV
0pKF2qtsAamA0I9/BETZjen3P8SdZuD47rFfRIhhP5hw4+ESbsbVVN4yTc6qxdnwIASXSOhR5E0w
z43/BQAzSU38TnPbkwFbhWoTcvoBJCjZENHnfJOj5OsI+vdJpsf3rNQ9f7Hzj8vytQ22Rp/Ru4VB
2sFo58us5YOIXjMkqvOehZGe+80DvAi7qw5TKBFJ82dz4e/G4BDYNmb8FDtAOKbb6pkTrRpIolly
OSTzUJN6tn7x8NYWnaJhRSBg5KYH9h2nsu5Vcm0kriZK3sUC8mq3XcRfg0/ftAaCFP5RQVHaoext
MDtGWo6xzeSbxX4sFYjLTgF/9WNVGILhqEUh5XpXscBMvzfG8F15GsAM1iq5R59XXIBoVzo0Sdzr
N9kwxl3jI1z7QiXOYaC6BQnhrYtXalQxsODwdjhhzqYx7VsXLmRvuifTWKGlclxTvMSZvPIZ/vGn
crbjvcjsHAQQ1SsEttncbaGZrXhFw+9C0ENA+Nw0iFuyHfo8DPE4ySshRcq/pQHRQkPjS4wKaoj2
ZZ3ZhZtLz8qdptFBgoe8vbQXq/jE2LHc3kB/yFj9VlJgqPDrEkL1BQIszPBjq6EnBaDUcx3oiL9s
Q3fTWAeDcEfrRG0yQpxvxug4k+Z40K5MbSobK5fieFtAkx7wFmvPphKKfVGXhQgmfWw0icRdj2Zv
2YNLe7iciThmq4IYuHPSKjEFcPqtw7xY0t59mz2a68se9x4oQn3QNzEERIotdaRsBdO9JxPbtPzB
vy7eNsdTPVDc8yCUhtmJhhSJ2dcpMHr2ISwN5aKowuI4jCfyysPRzIiOgdHfT47Q1CzhyOz6DBIb
slRBI0FjkOE9kYpuSwuDHgT3/HRaQYWQEjrDj2fOCp4vepgZ77QrK8NhKwsKoBIgJzfO448C8bVl
dgiT2D2KXYrpd3TgrfNidx0VYhqpmc987HSEACjU7tExQC2PGhW3UPyo5xIdMLYsmMxGZ3pSRrSx
R5JR+WrJ6uh0M3Qf78ATC26EKtxvABNX8cp/sDPWJs+8kSbsOAD/hHSu9mQU2hzyYAh/T2Olh5Qt
SyFzPsawFFKyZC+5XN+Lz1PQl0Avs9PQwfEgxBvXcMsSYioABTsYlBM3AvvrPv2bm/94Vkfcb5bb
pq5+TPkeBURSi5R3h7ezaVOHu4UWJEp+E5k4z4Zc66Jvcqq6hD0hK/IrSpNsbyE+Myr1XBvsV2vB
z22cGDkVsm3X9/NB6IoxLNxLhuQ/x7AjxDQWJXoWT35NY3AiNWCKD/DlDueJfig7aUs+5lTU+Ukl
2ZeS6Upn6WK741NFitamjb4JTwlWLPmsSKxwaiga4AAs8igdvRtptkNq6MfobGre6oKwFDG9wij9
psYwwkgfRbMZ0/bgjBUEOKWHCI8yho8fPKiS7iKk9kGfqp2DU7DAzPlM0uR1Ns0gAg+sJ4kvMI8t
LPSCRWRXvDIAjJItsSQQU8qijpN/cMeT9xyF8U5SfKNm6N0CgKVEVtxKnt8mXouDC0YNPVsSvWzO
WFpsJDeyMA/Xd1klj7gBtCBWWQ7KPxLeqTqE5Id5wIF2I18Xujz69ypc8wCa/5if2YbcRDn0UavN
qEp1rZfSMLwLosE/y5ra3P/TcsAouzKz++/eT8RHe7BIxBbr68KjJ3fsZ66aQXZQH3FVZqBM+CaC
/uUii7/KKCa654HN7trHt1FK2FYKgi8K6uV+vX+md+uzeazutcI2cWxlQuiaZrSZhnlmCw9Sgdbi
xSx9F0fqBeFBcFAGKefKb8K4MhMMOEAbHjZH4YSBA/NWWj+5hRmbizgWa3GZQ8lO8V2Kb/9+WXzL
Skfk48+lDH+F9uLVU3E/tOVzl64Cbt0jmrwxQ+XI6dAEe0bmN/38e2znwwk+3C1rDppUscF1WzzO
KJj/ihR+Vb7wSMwAbUBS/KpqVOqpPHuXh80Ze8x38GSqyAL+hUlX3RPvy5JttJvlgJunnhS/BdtG
L/J4iscbIsaPLy9x1JlaazxREfV8WpXwFUJte2BjEOMIeH9Faxqq441kvzNqCciFnpO5rOZwKOMx
C6DYmrnJZgcCoriPWKmLhgBEeOae1BJ416S+5ju/5dngeYCEOe013zCDKvV2S8sCFlOaKCUV4sAK
D+KUPWVjemHkbdtALF09MfvH99VKhmuIaQWl7FR//J+5cnZKt+IJUfvsQe+iyasoXpVb5AOtty0u
LPxS8UtIv1pNm75QaRAgRLYB6zfhKTTIOtmSOdu3bQrh2fzQhPnj4jOpEXu5fD2Gnd15Wx9G2pf2
hiJgb1Q3XLwvPg5OxNGg4CIxqG1lwy968z+uGiljvBm3zI0dq1vRtIodhjSpjgHfSt6WFAto3rd1
qnT6zDdiSyCHAywsAABqXxT5Pyj08HDAOidFWeNb/uRpXXhHe5kK60n2RjSrKA1tyU+foC1rRX4D
Szi08gt8IqzDHfkLCs8j1hb2Fh+cLT/057qX5MHZsIWb50SQ6LlIj7Ox9ZnEVZPt9Tt9IhKzfzMD
6bzqZl40erN0uYgzQTH1V6WbS7d7PQxVJxOqWV4ZD7Fx9sOdHqxQsUOcxaD7LuwJSHqC2I/kyfd0
Mnd0zJYj6Lhvb0xF0sJUbA2rXribJAeRdyn5Rh8e4bjm/kEb4hCPWCTOtSI/9HQZI/uldCUy8UMp
cLazR37UtzytsfnMLDwB80TqXD2vN7BkSVWtXgkSZzHZsBGJgGn3OsvtEONBkJHBlU3C7QrJwV4u
XNqpq387/ls0os1OCrOjwd/Z+aSNnTpALw7bOKgOx7410qxj5Yvs/TUPDzvXVRFtEOHRoAL/97ri
L7APp8lgdVC0Hnz0F66wQc5xaF9saulepAZ8oihu+/eZh7WDh+0ELktDRQnhWhgqESyW19OfP/Nw
rU3gPGuEi3bZq8Dlo/KiuwzF/At3R3YwSXsVkcNmYmAF83VM8NYNJm2UJdbfDQLvQuDw9Ay5aB1w
912jkwYzkYqpZEm+4CRiBH+kEJ3YpoUOKhRyflHWAEVyTcAx7IRAhfJKd2Uv567zAcvOrCErOEFq
AOP6q4s3emHQTkm4GpdOIco330TfmeZJR0tHWNCAbeJcGhDlRzytLswYtXhJVohjthQY4AgPhMYp
B8YX6b0l/1IcQljfPkntT64sk06si2V+Lo57ivzv/uhFsSDPnYzPdBYPAyth7biIYXahiKa/Pio0
OkiLZ7rBMeSr0OMjveo+qRzgV83E2Ws3REqMIJYux+sGvJ3FQldEqYkUTc/ntyo6ihFgV0UY5Hph
dt9DuJzyy3XkEYSk3qcl15SawvMJOE3I7IzZOkh0pH7OymnGwE1xNTHhJba1J86UyUkwr64ka7X+
y82oiTyNy3oIeAh1nUpQd7rItjquL536JT7CKksMhVIiEdicOKby80wUQKmWj5KOny4NcGxhKyTC
e14BTB/yzgyMj1cmmZ9MLmcu2NNHHnPeFhEVu2C+6OmBHe71IJ1I2oPMv6cquxnmS8ULccd3VqwI
NLQriymsPZfNdD9kX9vomWvTDicksoK0rW1W+//soc7eY+seWPRL8mlOClLj7Z/lZIltxi8A3HY/
EiL49cfEVqa0fEIhbwdzx/becPCTQIlJrPC7X4BKNIKn1hcgV0/bCOoNk2xkFG/pGuZ+S1QAMc17
aW8V0x+GP1ceF7+o1phmPfLUlvHV2yqT7m51mz0kGHOAAmz6G9Ux0CVY0wDaG2pjDlIDuaxVRVn2
HZ+f0+MichgaiidRK1voanErBEQsjEP3YbDtQlvZei+KlKWpGihmjxsPcB11mPgkn2ptotwHv2hu
DtaE/7x1r1nMSoQvqigFnH94K7ML0NB6ZF6OUEMoLy+odYMeWujRnjHs1hpYJIo3eYfHqBpFmicl
k2XhBf/W8sQFzgE84YgpzpPSbo2GT/Bl5Y6mLR6k/5+WaIpJbephCTMbDQbYe7XLwI5YAjOAY+z9
PCeIZV1PtwNpv0CnjWMBHn9YtWTkhRiK6hx//Ct3mUv6SQ5Y9pP+HI32O9HmGCa+uKX+/HHPkxef
G2xzEoLuSblFz6L/JbJYyR09y/eY+PliX0M8zBFRdeTjFTIWs9nlCn1OsYhdpV73gAZjP/RpL9mG
8B5hOdUNRPYleFSDkDSjAfLK9ZM501EQ40yCOunGVxDdclnBberU1DWPdlptgTWHULDWD/JFF/Do
OHHWATcGP+qHbJKdROYqD99RJi0gL0WUvDff3PkwLYEE7+HlQdC5dLu6Msm1rNElv0fSvBJuZWWN
bkgb3XpSfKMxcacFe7eYdP39vtGcy+aLUaY7MiLajWnhtZ3yzJDSxchcSdphASCPKaH3mddoD8Yb
wx8EB8oyuDDTJC3H5B5fWALn5Q/u8bwSMKIoM1XObc5NozuFMxeqsfOwOERPx6p48BVs8STRL3m1
n75Tc2te19ijNAfpKkDSHZSU7kvB/Eh5L65qRabO7tHF5RK9+j9rG3/ejvQBOiBNUzB3Mur1WedQ
0PJr6NPbVN+hOhWSAScO4Ukmk5aRf6hcsotFwORB3UB8Gio+i8KbZRX/DZNwQ8mdywoQTdfJqqFb
Am7I1dxkEQoYTOSjchfUdVwIPKF2RqpI9xsanVVFaOqx5zuKMUFnFHPRJOxubHR4RgOn6M76Y3VJ
rl78HzhgaPstNT1ahnOx7jBWJnYu+t1CQiTsxHZ+F/8swuXTwNiMK948Vg4TGdzYGkcP49HdXAwy
Sln+W6NbdDeWHL71iH6UTYlvDMX4Tm5VhpwXqZypZ8f9OAXOvudlhxclbZTAr8pIe9tZ6HyiIz1n
NF4VeKhD7brFe4cbah0zEwIee1GHqc9HvtXlWd3Hfk2FJVG7EFehY9FC3i8V1kfSmAMkJWv3LAno
IMX7o61Ixxz9dZ123JU5IvTWcbxzBNXwMrityQ3XPUxn5EGlnRLBVj2tAMi7bZI4IUuOeBiwW+Hz
I9JXFbKoiwRoj+kLGd01+ZQ0TP3NazgQfNduhMaEslXTr4bkwySrHvYK2+Ph3VCGXJvoHFltX9Np
EqhDtos4lR1W+8btDJINQjInhyoTJ7kQ9XVOPoLts8/sJCglr97wzGKghcjkU4+4r3AZcEF7AUoB
bwH+I6ykFv71JVg1H9v8ALIvwZ95V4Xfog4EL8SDF8v8atUtsEPtz+iyZOTbcoZhPUulTdzaLHSk
TXaU8WnAaB9xSYqZWkvAmsF9A1oZHZyty/n+siCxxBJ9SjdYx6TcdPqKCt9TMB4z6kOy8Uirbebd
q7QMpxx6aX1dtVoxQ4FKRpnzmRfKfZAQrhyUkbAK933EQ7Eid2j4FOQLnXVuaG+y4cHG2zgtniai
x/wSBCcs1MuBfDliHgWw6E5v2KarO7iLP/td7I/IlOhT9ALWOOMzuHio1987GkrQISa10FGCJRp+
N3iEI8nE4l+8WMbIzpbBrAIFo9uI8Ri4QddUr/HaxbQEHYkOBylebbM150UPYk19g4JWevk3BQGX
BHcR64lltMxbKvz0TJbUMgYUHyO/obu+RdyUR+WfK1a/Vb5T91lfcHqz7fzZ52CdGE9zZBGIF8Ie
+gvXi5ybqjVpa/Uh2Zd468UANQEmOxdVdd69zbab/s4QXLpl8gOLiMwNwTzt8Z+bR1MfQNvs/9/O
hTIFrsXklIBkhSXGFD3+05YxGQAmbOfmWIRBxS1Eb9yzDGbkbNOidCXW098yo4vxmgAOsTpT6qgw
F99fVWaEfOPkA3Ay/J1LIzpILaalU4X/sQ9vZ7ENe6ALx4lmWaDfQci9j8RtAxfBmD6UBURXzKVk
+2H1fRTUgtaBZYR9ye+K+JJ83yf5TeyKe1RTkp+plR46PZHKa49iL/mPpCAhJoJClOTuheUgWkWd
VGfFDrmX1cFjHuxcs0Imwx7w8QxfmacbNI2Cak4A3mdf5UgoXoddMKqOqc+XsyQ+bNFSR37aRuOV
u5J2Ok6S/hTXCScFRwSrMrVEHtV4NDyk+vUJe6xLK9AbxbsSHvjNbyCbtSY0qNh+miAxGQlU6SG6
u3j8GgMZBWnqCTfyCtIbPPOI9LrFSzwFF4g4w8FjPi8Bc8MGGjTFTnx87k6i4AdgMQo5wdPa7RX1
AUSSIowXy1JJfECJXstJAzAdUsJn14+NY8wn5Aq5d5k6Sb98YF2YrIkG8QpYNvs3OkksWIoF6fLf
at3O5Q3vBpFgwk5B6AVyNo1L8jFpaT63ddmliVM7z2vxqtn+9pwZoD4U4iJonU5lCj/leTW3elf0
91Jb5M/Y8GONEQHpJzSIj6V1LGEdCtc0GQgE79laW7buHx0xqGLV37KFBthUM9RGJGqJQ0gmzXwh
1hNZU7jw9Irkl4ZdedcvEHTkVzK6NyjZsLpEfLc4nnwwomtDecsgT9qenKk26porza84WNdnbzhf
KA5ACDTnwTuw2jvXBmYM2/9ajlph0gc1ebfDqtckZIehkojkGPS5l/xC1/gCwhZBkrretAucs6cj
0IhQrRNCqwacsnntkCy820Xf7O2VrG0WsnFwcC3LwTadDoUEhk89yJDHYJIw1C+e1cCuDmtzGKYb
TksjdTJOZJpf+PslOpDr7K3hQ6Tq/o9HderbfGM7bP0Cv2wvNGvXduufSmZFwJuseEORAHze05vN
9ff+g/MiTZQLre5QYeXk5ITmG1VlHDM2jPcNcyoPMje454Aio3zn5OGhwVm6f2onzRJw2lXl7uWN
8zL2JNxwRVm18DBjOGnzpKXaL6htZXbuF2GDmpFrKXTk/fbAfqI07Xgd3rMIj7GOBVruItN4BKH4
xdDMvIz4aMX/v9f3KTW4BA3LQTFisYFwW4Vk906/RDvcVAGkWk42F37WXVq/r45/0euEZGHE5TOx
WBThEM6ol7eDiv58rVYO/UDWqTKPJb9/6ORDOUcw4chw2PEsbtPEgaAVJy2sHD54DX/dQJ4FHAEu
sk30JUUTb4hfoZSElNDJhS7y4+D2Wat87I6UM8iXCVTA0qqXoWwbMIPWEMYkUy2fC9b+1aEiAyFQ
w1vvOJFVHf+6VKMXYUqDknIygEyGkSTVNYyKG4rfCBRfHIZrqDju8qah41SwDg13iOT6C2MJgufv
shbuLktazf6Pcc+nfSWc1dxffaemiAM9eCJTvvWVtxo86sG62Z5Ox5/3cbxfbDlW6gIQWbUbQ9wv
9uIR31aBrj/cs2lC7p/tNDKuMcJ5hyg2COzCKAUWjRqY6mJGCDhLaeICSjCRCN36GAYNFDbo9CrG
0Qm/7OUhMLyC8r/mklHjZIPgHUEb5UF1Yis6ZYvznuP3CtiuGSW9UUaF2Tzc+8mGSJNyClpdZG2X
83/+VTjEHcoW4fl7toljG+hkVIdyRyyfJgKxWkwj88zX/gAqVZjrcm2+mFWwqLY3qdpj2ESKarn1
3CHUVw06aXvD68w4q1X4KY0cKBvOJdDfiNEzqhcGfsuoD7KZkRDE/Yj8szS7qaHMA5XPm0rohhwG
ZfVLoX8nhEwy/gSsbNocgOeJY+IFhpPsguya7zqNZllukqb+vBJuFMTzTRu4LQZswZFDBIjW+SEs
Y1FbdDRJMjHspO3emY+CGwfi81lG4/ZHZaTs9nYX77PsZr9F+CvGfdjHXQIufH6whEbKjB9/eick
AqjiWtUX1aIEe2VQMH9YRaE7LzJwVXjZgNNaR7VLMINSRIoIs7TVgOnR26Tue/5OKK79aoo6CDZN
30pfRQo3mrVbxtC6HBVGTv8xF+qy7y7w6gF35kSBJA6oLq7KCVZmJnNYydcCyz4waaSFAe5y8aLM
zzkg2Kc5ya9hu+8EPbH7Zf6sy15aLiYIEnz3Dlt21ZU277nvRHbn0oT7hTbGZi78fJ5OOGfPV4c2
QHbz2c38iyr0/e1m4T9B5Uyv7MQt3aKNRgbwWd6Gp6zy1QVD1FniOTdd944546+KwO2IxdoOo5Cx
ateXm70wZ7kS/xuG8I6Y3iIgfDekcgamfVM7MV6/+3vLq5ebHJ+vDl3YUmSeJkGi7UXn03qz2P7V
sJ+8vn528/31rgrrT2kQRooApBSAOD4vAldpP6IV8uc+48Cb4DiwAwoGvPC9mXs65Jfr0sf5at1G
AJqGrHxKCvbPPcrNukBQ0dx+ovtFBJ9zgiXvUa6Y1n1wXHzXGW/Fn06Rn8zden9GvkCn+/HCBi+d
VsdC8Ttkq9YI5e1tTcDlsisBB6WAeUgghZ9oOnm841Apk18hLyeLGouxlKP7fBNLRfzDRe61D2ZE
lSlMOqKvdHh+C+relQez0BYeVxFFSJeimzrouDgDPpCvC1xMjxSpf6HBJrzgWa24/Unc6etQsPef
X/JMbpI4ppFJUEyyFAeB+smEoeJwTpgdRyhUvQOECEu7mGPBR1OCREMZFjGoTjvtEwvR1QIVFgFg
PZantpnF77wdpVXZSCFsmLdRV3F5o3tsXpy5unoCal1B90wpLXOnxda/BDgighRhqpKHjEc5WT7D
LKAUf07AOVZIJgwJazl8ox44ZFg2j3qf1OzdCWfWD3iuBWaOvRe7xGJQ0MJkaQ9Qhw0i0dGP6F2n
dHuhGlGgXGtwafM8TUApACF+LsZ8F00GdqOCD5+KvqYYjyFgkgudWwZ4mC55rzxPdUt7wKpZrCG0
CsoBy29TKLSBysFyVNJ2l2GZG7W4/l0/uMPiaJVpM22UliTEqSXke1uijDzT9k+pRQRJQL1d1sNv
wVa6DXCrR7y44CttT7mX8244HayCifK6kmlix6IHZ7tJBq+FU9457L+OCLXXwPAv5JFWzKyrW+JX
fLcSuLZu+H39+YcUSWGLJHwPgfKrXLsRJcQHmvs0MVmBFYtK5sVEBaUnna4ufe3Dz3KPlshA1xsK
6xlNI3kILPcUL8yCsKI0kC39ThXHCBtFVYMilYgZCopyNPZ5exBk9wYXPgUHTA+jImDVrTyrtNzY
CSPPxKD6ncbj6bO9FyAH9nZzEWc9Z+Fb+eyRfvA3hoKMYoOe2XxUBOQtx3WyEmpyZ9XMWetHD1Vq
ubHb9raXDfDo5TE657worTvku6Pit3NJT7dTXK7aMIZhgMfJf6AC/dm3o2iKjM/Q+77UrNpsn2sd
hXJR5I2+DcO8kLbcy4LlSWBPQJpCHPvNRAfm0X81UmRfyKYBp0Qeo1vgmT+Y+t1ooWzajNDBvXOs
sOG/3OhH+ImkhMDAMg18Ll5gVLVVNDhzVbqgEtp15vQYHvW2FnrMy0orl4sB8SGsXqLLLA9/qcou
taZ62lmuL9DkWHiZXhaM7DmrkSMkW1LvaFRM/vxgIx5G64vnFAHiLW3hFXj9wXX8X/aUszbOvODf
DMqfWd7LlwB12cqWXU4AjPO2YUFxRtfh71JDMDNQaGyiYGVWv5tO5CfdHzmpjQwZXnjonyb3W73R
XupCHq2xD0yyDCGuetwlg0XvQoF+IN4/jQdCtzuDxzsrgrN8WNrUrRqzc8CDtfMaIpNzk2t3mf8y
oQusxR5fKKwhBngHvKE0PUOKN7Pf/vlh+rbjnid0LuELL2dUERQmi0almtJ0ST+l+gyLSoN4TFzj
77QY/z6wchwggzhXoIyQH6MFpX2kG0sNolO3EvoyrVeYXWcWpRz8RyWrssxgd4pVqZHTFXmJUhMN
B0lrYXhO7YAjbRjKqs0RQLNR+q0HyvzdRYUvyxUhCf6oxArZc0yf3gkG2MyYRwlszGq7ZoP5iBX5
78hma6gT3Pp2DntVEYxSWN3BzL0dVxzex11gAZNICuzlv3P/tEl9wHKJTykPzVltapFVA/HIIZus
0kM3BuqzgaauwCSXTu6SdiFV9xUIJkEEl/pmdYeyu9Y3to54pszeK4hsaGgEBNm4ElFRETYltQX8
4ISiJbKw/2rb8Zqlr0XSs4XDw8Y0NZQITal11sDJHRGEdoVNXqgF9Ll8tDK/QH5N5KekuBzB4F3w
a8HWbIffaxTDoariWOerydF3LxnCHAG+lwh5PfVBgiZM7F2nx6pXvVQsjqIm4kyB8oU7i95wFaNv
LuHukiMDvWYiJyYDH61MHhNCOSIhPy2WY+r2Hd7dUX664rLc8NPFgk+wjiSofD2UdXUFQMEcU4rM
a1ZbqpnleYtNbbMYB29IROMO3fjUXC/8R+s8XbSuJ2vAJx/1tFvR474jYUgEYur2FBlPUt2HU5yu
DsKWklKopCNIAKQJkwFQY6odWvIvkiwxPxRAmGuxVlfdEGOj3/OI+ftL4ZoUWvfxqSMCiy53boeV
7swUiaCMn4gDmRrSusXhBzf4PxL4RkVyCajDuoT7IMVRoDaaHQbhxQtTgWRD9RHyHvritq+JSPOH
zyqArBfGSzbTr+Wepi2H14WOroxuD81lOhickgEbbyZoAUJmu4h0ZITqWH1V+SLcHaFOJvhPQo12
pMB5JvcUM5XRfOo1acLQLaJ4hC7N0fz0dGK0R5zMoVBayHhG77zWZlhMh8mMDR1+KkLLwVglyRh2
O9GPkdnyvsNGBNOCeLok5xhV3Oa8pegpjzz8XmvqsZneTCPDYPvD2aJ2ge7DPdwEsFTkyTCuWcHy
0PB2mvqSsDZh8NeFLUuwahFM64oTWDRvJBFMYeImeQkytnO3YUyebeUqNCKxhgwLz56LMfy+E+ab
FhHNvuoyqlYuFuZfLimkIl0Gw8F1u6G9dOyo4/9keQY3USxSY97meuFsuw5Ptz9uKmQBQYRxXJt6
HP3Jmb+k9C6ZC4STjZAAOxlNOHFhZxXiEfWGSVISD+SXr+WflewiCC/Mv1cRTl9qVpf7nuQmlM1R
U4iAltV+MaaxanO8OoREqsC8CsKbqMEBXEQUh+PZ40wJ4z8lp2l2adGV2zB1qoWjEt2PbY2NLE28
UtgYbIvGZagzKukLOcLPulbQF/iy2K0mIXaD0sC/e5Hq/O4qNFQq7MUgLWt/w1NHFgmpI7NZYc55
aJA/qALELuHLM6XWTJHqhuEMS9ndZbaNg5rRse75bfYupMuDAlcxMVB4A/f81HVyd6gYEMUSNAlh
MMvgg2F7SLjp2ZmOT3J4x7Q77+C0qVeNY1x1o4jlAIKJfNKCO7e9KSHMUm1Fm55WcWxqE4YEljkc
FUGW+lpCfVfjkmzQzQjzCoOckpIBrTghkg+siX4kFMewTJuVw+TlsLFhkMAWeN/TPWw2o3AklhuP
k9jxiVKLls9skdbXajgz8F3Z8Kz7BGCykfNxTZ5sVlMDY370R6UAFFVWXasuRjhBo+VwmxuyB7DI
uKZWC9ORDsz/BGSqcJkHj4Ed7DwbjIMsdCG3zKwB17QfjmjMU/BAFqzdPX+Eb3Cg/c1589e24Xnc
7YVGR3Dwl/9iodsguHVJp65f5VGHPQ16ROcvxcChZVPL01qaO0Jze71B2xPQnF5Lpp+Evnu0cF18
Ak4wVmd5ogqNkR3z8AlpPVMmKx0xc0ZuGXEJCi4GHmFu0+VfwLW2nI3TzrmxG4BlGbB1tUml/QY2
Y+ik3cPxDuw2z/ANwmO+kGfWD73vlWTlm6Wafpd9i7piFoM3hwi9ZtVF4cr4+7WzSNZJ0JLIFcoP
3BKn76K/AWJXEf5oM3UtZMzTPTntYPqTVsjwDznEyHk2hudNppJ0O5uYhom6qyZofqP7xveYVYUO
CO8zMnufkfYE/T86i0mhLIu3W3Vqb4hVoMvjT4nuJFL0JQJT9zAZCQkDV7kXdAqsV0e31flkJh7P
B20VwQDWUV07PoIMSSq/TqzTIeA/R9vEtFtxj0B85FwTdjODci74tEsI3voYtwmXcyNzq2WY4mb5
7zvDTJkwg4yH7GU+oieiCZ0VXmfPNmqqv5PKQaYOiQSeKiBsGsjOsU6zjGfl+z4k98op1spfJveV
pEwjlNvgiHE+ldJG9OC3DLQk1sRB71XCbAiCeP8uPKU4cDSBzi3x/dRxXALcIAp36krKulF4aToy
XeE9ZINDu1aRhu9u8os9T8vaOHHBtf63sIlYvWMFGhJp/7aA1d0RnOp5kzTYw9PaUJalnic86Nta
GuUhKtIR9sN4lYLVeYJ/7WAdQ5FJYLJyGlraAh+Aze7jfgttqKndC8eb8k31b2QCNFSQrAH7hSX/
hG1Ueph9MzIzyGhE1brS2/eTlViBhW16GhnKbeg2dxgqC2wKAp0GSWlw0fsJdRv4KZG7HdkF7BA4
1r1JuHHMuBk0B4kZl7U7cLz3d3f4ilFHkNMWhIDmm0sxVg+JGW4P8dNPFE/29KQV9budlNsEelIX
CY2GmEj1q5BLo59vDHhLeT7EU39toa5AmFX4Kb5eFinQIwQKKmzSspXBy0F3c9Nu26RLN5D7IvOS
YO+dlG8b0RrRWQJxtiKRapi5D0aVPqrTWfF07adFlT4UO5IYJPaGdo+OaoQtSElDy8LQS7/xpe+i
lSHgbyGIjMAvm+bonxP79bunVZnX6oaigQZXzsErKYhB9TXjWV6e4iLGkDwx92alQvF8LJJnBkqE
WM1wyvjkTfhZ5hKI/iKTjsHUU+lel23gLV4sr29TxT2TjKuz4/222mPNodjFYM1N2rR8Gbbxs1ZP
ZOR6lW1OIh8jwA7L2mSjhnthjoE9bgf5YZYYG1m3sFliKae8kzjgY6OdzlEbGMcYlpTJ+Y9rXIQJ
K7UpHPJ2V1PdjVVUwFms+W0uIRnhPm1TkFXxRjrCH5ft37y64sO8/Ndu4MuFxQ65lm7u0+BlmY5v
EZ7AO12apwN9sb53mqMXWBgrbHdJtDIstuTpR6A7iD9l0CWBnkWOm7XfliezrhymbUS6Ib9iHIuh
NGB2Uo0UaAT6Emhi/eTIfnLmXUJsOh6l1I22XAf+C6gZMw71TrcyMdIi3ZMmMxrsgHdJl0GTlf69
fOxhn7CDIYKVbWb67SEaOJRdHsU4plbmI+Gj3yHI3PIaO4xWbehlcyREc52iJnyydCWith/m7Fg9
v+9SuDFt9gooEu0OhLdjHQipAjaU9nq8vDNVEmds2rAQIZrwsLQShJtWUnzVXy+w2BaB/RoYWS21
U9ywLWsjs8KhURHpgNXcJjMTqYR+guyAlRmeFao2F7cD660oFV7G8Qnx32rMLh9Zf4oDJRHc3zbR
olYdl/Jto+aX4HcUL5xJOc+1nSRnJk4dvZ/BbcQ1qvReDFRtNI1JnyqXPR2y8KywniAcC3g/nnHF
Vpjv3HERuGY7PbT1JTuG4kKkalHo494DhLGTriq+J1Mew+l09jyJuXiAblmAVZx4tC3RFshZh5RH
1dr5Y3ivuDzM4SWfqyUMagnprz/PLh2fbWG3VHtXK3+Oz0LLlTaqyxz8PtL+RA4jcR8j+9Er5jOu
Xqc3vbb4N4Z8BgBLUmIF68hOiBrFP9yGfGAJPnoWf8DAXJ6Tr0AXoDGVqyjFqvPlsoumjO7ug8No
JQiSmfP2l5xrbWZSS67rrYBQRElCmaThBqTPxA8Ed2HN8bISXYYATkBtv6JYl8B1+fhU9LXncH5l
MGJxjo7S9wW4XxHZK0A8P0a46SKnFNASlYyiXoDcx2Y30qZuZM/XwNhqQxVAsXsekGvyTuC4eURe
M7MiZJNl+e4/fqUWtNKKoYeScSGLB1gVH31jUzMDYeQXTruqAwfWTi3kCIWjGHAthx6XjdRNehC1
9wr9x4Stp5UUXK9LZsWmfP5BorpJpafUHysdwuyC8u7G55V5qaQ24BhhqSPeiUOdP659GCRbwBgu
Lvefnz6kmH0AbLZwhZK3epOo2aNch2XJAjQm2gN1Pq9OSLIYcSBjccxoYV+o30XX9ZbwJpGWEQmg
dn6qf8RON728qJkpS5NVJky+zVTf8dGFS63g8RPJoOjQILOtnVCH5Rc2zZEykhfATHvMvNjmn8Dy
XuBiBWET65clxjqrW04RH+xPtxy1pZyOVaOgiZdEgy8g6hkBltT04U0TbiCqjGSNELbMrjXwFs8M
AkMfJWXXW9J5QqYd3OPKHj8s3plqt1SmSn2Ty198u9mZD7/ZrSOkaioBRf9r9a5ST+2UkcGZFFLr
zG8Y9qlwoPJmA35IDKYo/qBjNKCBTO+1Z96YFDKlHClxkoYyvQpn8SNNt50X3dMKhZI1aFNWs9Hr
ca40EoKQFhOd4pzg01X7DAJ3/RTPzvEjAsi21G4bbc3lytvDqJXHyK03SP0gFK9i1tKK6sAje6eP
JnSFSw50m/XqnfHic++ttpfIZe21BUU81zTTmzVDGv9ZaaTZsaHGiXL73oa/ed6s2uLClS3H7tTt
x7p9DYUA+9apda4oLFUkzNrtJQm9SC6QfRMElCL7fFcaI5birRzW4rUEGvkoDYoY8aTQC70QuaMk
2XTuuIZ8/KrzrrYbQKnx+XZ/qdCIGPtgAxW324UT/Hh2uoT00e3ekYGuyeVQ097PHD92/94dzBWP
jJUQ+4N/lVwrAExar8cBc9HkB5gwXkt8QmiXt83nbCzbjxSRYpzzjzcD19UOCrn8HPgaHAHReJx4
6VKOtM0DzCkDPk+/p6XVDB8LX7DfWXytod4X6jXPqRiiYgCNSRXZmZ8fT7HkehbNE9owgZGx3svj
8mQb845wrPvvGqG9Xg/oSUB9mcBagP7sFGc6fRu7BlEHemglGJhjohYqiWyrXbJbnDBDtgQYaCI5
EfE4ZmP1vaRmmC/uSmx8y9t7E6sH/Hj57aXvtOy5iB+Tlbfo+O7UHBA/nuRBoNOVeLi6TGCXEDEL
XIYmuyfHL9/YvnntYfaem3MV97LZ3pSBOhOL5y8WZTS1p9e9iBlbHpGIKqA/l7ZtT/QLw0yeXuVl
3MG8HYyxsHqO4wKuIPtMTgxEPhBN6mVfNO1JSUbowzKGNfuTGV5r3W1eXNzdzeqkDZ3Xq3PimXpI
MJgT/LJeU0m8Pq0PWgJETFQgUaxEqmjAbtqtKwdWmHlzva0rpt8dY+rubSAMEmdXEjT3eCsXiBnM
VC2mV/qfxN9pnfT8jAizGv2aCHXLKNfwPytQ29dkwQVOebBMGpkP1l2WO6MoZvjqBbE+UIHyowF5
e998UuS0Drz24HdSxDtzUhvDkcp4fWtgOn7u+Ev8YLpKxCJFUt8ZiIKzU5zKwP907lbCzBm7DcaH
5bz2td05/hb4k6U8AfkFWLoA8ze0hL7Gil7w8ZqaBK8uMMkwQyZ99QoxbnkkyW6LecM6TTQoq8R6
nSkJ2giu+iaOE7mMm8St0E5Uhg5ZxmdikoH44yVvBgzOv96Q0XuvAV2HHCV3Fmx/8DBO5lN+l56Q
7ntRtsCZXRYoHvC8eQm/vySgs5XL2nq3ieu2sDBscPayDIWn6Xv90ZJkEy5COQ7mupW2yUZd890Z
kLXNA9MsURBrrhqcA9X9D7JqxPypRDRkNof3rwiO51GpWGhfAhjJFm+9X3LOBldKjmGVMB2WbA7R
GdY2ad2nrlPDVBOZmkumDDNQTd0YFtapRjJDtjf3Ab4TjradsnA/VjANoZKgUs1IMvNse3x5x5ix
1iKI8n9NmXfvGqykBMlFhwmEpxc08ZSS46/HJ4DHS+nF8KLENpwITHcp4Z00bjL3BSs3yeEXzvR4
TzE3OSWRUh0H6CpWTFcmItqe1TfrBLSLBdu6dTaGhpxdX67sFeoAhMQpANteP3OZYFnoaLxdy63g
JzngGXldXqQ7/JL6wPeAu99usRvtxBmMQq3G4TbfxcFVIyRgkkhJSrJNz3Gm5oYVL1TkLgiTlLLC
yqEVx+nvqGa0BlAVu8mwksNF6k262qcXISpoXR312ZBf7mJiF2tTMiRqh1Y1zG0Jzt2cBhZPzIGT
qjOWFzHoqGs6Y07mfbD0DxTmr7YQt+e19xb4iaWKAgf5kx1no+qSE1FLK94Gc4VNp6KvEU6b9t5F
q0W73SsEgAlVaOs9voB0DvOivbrkX5QKEeyWOrsCZSiMnsKusPJWtB14DnEUi/JpR3EtGxFXIbXz
thxBbXg0nBKHmSpO/ekLCsTxq/vNcwRyG/s+P4jIYpDxvgbg/3nZPOw96mmjueNiNn/vSDc48ChH
6DcQAguO5z53glF1cgg1q1q4CQz8Wcszekwb5OVeBKpoi6EEY5zdeEFruW/CWbydOnLvCU1RvAql
Wg3WhcLu0e0Q4mo2vG18/HV4OScywMg+Dwmzwq+HUzbaYK2YhhCgJd+LHnoFs8bzGVJ98RkpTCPP
1YPsqTEQyupEIsg5gUfpLOYr1tJ12kgQura+xJx2tYD3uQopq15mrEOTAuo0gu34PRZPzT2KvUqd
wFx0e9Q2eGb3yNecOrDf1CPUZTWgQr3cP8ghhycF1HIIIVcSESHqaeyX8ZigRE4mpo2nZQPSqQMn
Ge7WFPIUoIrUpf1sJBwGE9RdvhBR49WFoDMH1yXobXfS9NDU/fJYXg3PE6U2NHYMC3GAuUZkxSy8
r+/LVduc7oFKBc4BBDYckfmk9Xiwix0QwJ7XPVltXNsWGoSIkrroYCsUDP43ck+D1X16VGAVF5xM
Qte4ycTIIV1M6k34u4+l+FjqAGVZofDlp5ADo1MVlVf+cxmyD8/IdLTuz1XsIVafLD8gCGRaIbxo
kJ5kBqIBkb3/20TOPBCkgM2LuFRX0TZtRBDP3LrgfJWOM2SFkJRM49FmnF8ghd9Ksmj9DRrAUG0z
jN4tS6pznT+mz/l8r0S6wGvJ32iEJZcqd14gUmJQUHQTKAVb+gEloRJmwzUAz4T7yFT9yIvY73q+
bdgYDdU6aRkMahex03N5aZqbS8znMd1akRUedGNgC15DOLen5nSdVgioazYIzoRoXH4c6Xvx9hMQ
na35gYrf5W94xoCCbNHE6eb1BTYemLBpmhl+lK16GiIbbERmj1LBIqSpMeqHcEBzUkC08fThsBR7
Lw6qEoyDFbg4PdQwhrHAWdEFycBP82WyRLqC+d83AyMAP2Foo2LBNQPSBG/b1i3nqfRfS0Te1JUL
MQ9r9BzmlPzSZehk5QH6Oh29Ea0I/nLtDLxtk8iAS8F7YehlnTpKqsi608WH7+s9FiM45u2SIhzk
iOaNQmVIrZfQbT+pcd7jm6YySCZwZQIIoP+US5IycgomH2MkY5Jws/FtqoMJlRcHt6Zw6LwPBaOi
3hFayN9YzVFF+OvNLEL/LAGWeNhG7ckRSZyMHc5O8itM+XqCZnrTOkzP1PPCvRxw/rXtZK2tKKs8
cLs5fb9tbQRowUUvBb2BV6bAT3ZpYHmxZ2qoSzpaHZyd7tda1y73NIosJ/wTpYRvjh2Zea4+c4h8
EFUpyVc3Vtky8kSaGUEdXQ+rCUC7aBhOmw2rjmeebvvb7/qvcKb9NuTmaiJRVUtJtVr1UVZy3by7
rC9277529wl638EYWthA4qx2JvRjxcR8XDT2MEO6sBQO8+jtr3FsnI+27zNM1vP1m7D8uCh5x4Wj
ZBkxpbs/kuFQHBJ1xRerC12gWKfR9JtJJO7ula7BSWujhnVFFUmI/ba4Oyz10AIb91VjVWhMUsmF
onpTZKhSNc/y7h780B/Ig3deEjp1xFIWiTYFp1CrX43NtU/F27zu8k9vgx9OYL4dFEsaPu/TsjcK
Mrp04JZ0YhNN3i5PYZHGbpuxTeaPMiv/UWthJhknAEEDCmHsO+COxcFAkywEkuBKOANH9mKvPZRJ
32UjkFWyjk2Br6HCBAb5NRPMA0s986E1Ba/MDi77FJRyq+fFXilHs8vrnte7wzL6R6nqz8sF2Tlz
MnIWUjYU+FBkPrMxoJ4VwjtV2C2dFUXXElC7E/RDUtQdmwOucrFJpK7cWK5U0lfivSFOwLmQ7WHe
Bej7SmkTWksOg7j6LBpAWUz8Si3Gtg6h26Or3ZaE3C7DtM8wSSwPbpCCgYEr14PmPuqyILNGghWb
TZrDmeHExGcAFT7rAXxDMGt3Ml8CbEKlbPX/vMP3PSviRUkxvm8S0/oJNhXu0f5aRZ0MpBEtYbo8
R3cEYW7emrTNMsZHbYYBAQCN5bueFgC6BqO2rDDaj5QYeSOpelaejN5i9GHJRU+aUjz8i8/snHa0
/vSFL0l9XqaaWubVoPB3iPldyNHn9cc61mEqP600x+m5Nzu1MGU1Z6dQkN2yMrGNwSPxrqHdElAl
ZZ6PamGRLPr7SYZCoCcH7smMTKIOQ4GubsXqrNFhZ60A7vDNzqjTj4mB1ZX8T8J+Mt/JhfNYPlPI
QyNMVQ3Cts9T6uR6DoUS3vYT4PjzPqmG1/OXxx1eUCEhtaIrLQ/12+ES7C1hXViuke8OWt2+yB5V
sgMLX0uZ5g+1U3sS+rGqxyjiJz3nOV8kekgBOk8Q/6/hH8Ck8cXJE2RJFVksTgrN+0FWByMEw6In
pP/BgdW7RclmPPwGPFmo097YqyWMQa2DjeXYeuYha9tZcVstacRtmgr7Q0EDASVhWmNzDHh6WQd1
ZjOY9AuP9t7GcZmgUlyneGIV5N+LsWgFyiKyGSc1Yy39FG5TGJSFfnZ2eAkpwSqV2XbNIOLtROKu
Pp52rrtQkf359BfYV2h7AifxA16Ghlzo1QNrBFra3oRdQL3gduI5JQj6XUxJtRV8wFg10pEoQmnb
vLk1uOeM11x2FZf6pwukQSx0Mwoyu563o4m20pSpzUts6m5X2F+19rmTMDU1kQlez3NZw2cu6NhG
UNkBN9Qg837kUg5+fBPv9llf6U6Cy7yreXfQPkTMX17dm2evyF2ukjEteTt6Kto2KSjhgQJbYC9J
H1egLaPqvpsb/OlWbmzGOJqGHPINXuvvK6eU6XmhOml5nkOqw9hblp4XmENH+cIi52Za+TafAuSs
1kP3/4P+PGr1Asf4zXMKxGv5UN+Mb1awJ8y451NTbCsu4m2OrKMjGjioAHSrzF8ZXHTQjqXf1TTF
2snIjQbcl678ssh0olXUOQTl1MD8RGPFFU2wgSRD9z5Oen877khclxbyS1D0y3XUhqJYq0bs8p1f
KpIhRa0pjDOQo2Yxu3UQAX5ib6whqGSWxlZ8fkFEqSFiyJyZbQuammpBrNof7hUTq6itKbfRcuC2
BZMX7x7bjkB1Xzz3HaMpxsDux1PDxIEfskHSu0DPcipkVM97pCiKkkwpBY4kAZX76MaqTp5ELZw8
JrWV6dGhQ2A4b81H1IERFNiNVP670xbmOubCd3wBXinst1PQ6jTOkSR70rfzvY6a7RIeD/HA/+Lj
mrYkEcd7mKHz1TwzZYKc5Mro4pvsni8whzvEZCJaRPZcSfq29tijSv31P9KH2jjU/C96czRr9YGm
sQdUwGB0Rdpl5ldQnfBC5O4G8txuHL+VWRC/M7pF/AVBlLP0E5JAGdMqNC/9wXosnIvamjKLP7x+
61mUgVlXdrc5nIRB3fcMezKMjlsPQPEX5viZ2comOMT11ObpTmYfOJ1lItBpdKw8YRpiajHQr8Up
zbEiuHue7QGmR1HV1hqCMcL9J+qdveHDyIzpIM2FOoe1vPwaER2D3nnzLmOT9jJcmsWtsFWYDVQG
POd1Bva2NGj0N1wD90e2SEXQLvLFej93fVHPXv/MDLzcvFTg/qGClQkRnFSWGZqp03igWC1YKkcD
yMQRq2yMtWIGi4MNg4lZhGpHgpXx2Z6z/YRwOUnweTjyHDoy4Ga8Xew+83M18cQcNrHiwlDP4YrK
ofZKDzczQuOcS7w4iLnVkGdBqRVqnZ335jCCyaixPJNVBR91u+qqSYt7FJDKg2Fy6J2hGGDcVnsb
AFaWI/aYUH2Ko5+Sp5IhCTfTOoHRStl4zWedTmLsL0nqujt0LTVUehsfkVEu3Aem61Ql54sPe2o2
A67Ou/lCKzH2rJckSWDUnqEmrEHfFqC029K7+1TnxGbQs6kAkMs7NDQsC3eYw3Fx/zy8tt28Dyyu
tqhWMxroi54V1K+94queLpwv1krvjrkmJzImVdmTPcs60Z0+agQtfO1mJ/PWAJlSz1WhS9Dh2xfR
4jbw3aYgdLepTi5Y+G9UBjTTHoHGs2dlccQDLFKIMWoPBesetbINmkW5kqa05J5NvFT4rGk9XShV
FNoWuFayoYJgRksWEF8DUWxpVhjPyDRizN679rrEkHsG/a46yztAaaS7rrujJkof389djJAvlKyC
RYlKt0CtnQxKqIU34nN1fsNUubKNQ8Km2EYx4qYgTEKvrBAkbeWXAtUTdlgLcYou7VFE+woxcSjV
BeV22YD+3ImQsOthr9I8MlBHym3vq/ZleN8UEHt+QN39f38N8wf1wfA9/nYDe4hKs5/eIbrRF++4
FdCtUrSXptLNsnLGKMnuxE1o1LkMgH6Lta1dVWQ4YDed/QYn1vP1PTtdznmuyvG7u403YgHZi45r
J0kZRMamZnd/D4Y0q465SiyFDT1JdLf08fziCo8ybNjorlIIzevFNc90pfM3+k/n2JA7wfDdgWBg
PBv3Gdsc5HcWjB/OTZJlGsBOhfTjz7DSMQxQVSC/r6XE+qBqXjsB3fT0ldCkO3voqgmLDEfx3iXg
Fdl8zxXCa4SkQJTa39QhTB41tHbhCQs4oKSfmZ0Kls5uNampOffZbnfSChSqQa0WDMqkAPXIJCBi
Sx5uagzbiiQLfVvhCG9Dnv4ZQ4V95Zr2WXz7ADCSOAL+9BJFnBih4+JQWB7wmg2ROyn7qTcd1xLm
WlTRc6eXoUJtw5NqN8bWV159L3sqiqjI6RXDEScR2Ko20FKf4VHDg53k8AodK+0cJmkGYkJGqHeS
0JMn9pRdF4SUInF3jzYR5DJAkcc2DHtrCGUeyCw7BQiik9ig1Zr2MM0hCVPnXQ2J1UKzTNwY+8oO
WxfuWmP7ouacrw9tsmVV6tN3Jg3jaisfTXCMW8zKo/RZutR5xIreygmmJaBB8do18ZQJjwXc8ELQ
rTGqw4R70/Bpc2c3EkTjz0OOtcsG00yH65A30yoe+38v/B88L/dXKC2lk7Fj7+WpE84bdUb+jEeH
7S76bfYTDUT764Z0yOnmcODcAwCzpWQIsFP7P2OHyZhbh3VnVcP1pXt2iXctIeTXKCydOgKJK+dv
nz/UYrSk8sM42/+4KzB8VDz8Ncx/xvsEVilnnTlZZSoFWFdCgts4waNU7NFrLNNb7VsHRwlY5l7l
4R5gzwgWzLcxVETjM+N6FV1rmLQ2jzJ4GiQyr5rgctse13dlbf1VRiWxv0rXqQICZa6SBrrVmN1M
98nIv/qjEkXMbtkQQSLQieCQbiF/wLhZxiBPPUWsP7r16dZGSmAFEb7ivt8kUx1jd64GCyFW88ri
CcdGOc9g69lNmW8tz/HSaQgC8nROSzoyCLlokA90nBEMZX9ybgTcj6OJIXZsMzjMpegfj4CrEiOr
PbcXVkx/GvuJ7fJ8OCTDdcMyswPuk6kfmmFv1gblfh0ldNwJEadc6LSAX6u4V47kUpg3i6lv7SsM
aaXu0JDlDunCWU2D3mapBPXG9OOtWbsAeeci/hyKj3PJpJgHkJQ+oFAuayPSujYqQPR80dMlDXux
bLnHMN/aMRLUsAn/SNNEwlhAVCuRuP/aWt/RpwQQXWV8bcgCLEHIaBSnLWnR1JYC72KlgJB8lYwp
kQ7Q30cjfZWCLO+8ehEv7Z/ZEAX6RcRlx5zc3OH6CLvCGDvhzs8X28/N22tUhLT23yUloSQD3gr6
Xb22IQ/m1zUxr+p+ee9udnO6VvjFeMtqhOnA4g2DvCfco4YPBc7KbH9uUR80cD+fr7HVM7CV82+q
6Psx2mqqphl0DwW1w1soTDr3kVfBZreW9nKVONJbTAOIA7lUwNqCyUhhR0rlZQr0E8j7xRAGZYrc
j3s0aDknGAn2ZefREZTwArukxo+mISIwjTMros7sBRMghImo6klf0QIRHEEXW7CsfKFHabDn8mQ6
1NagQ90A6UDvFp3KX2eE/SsvOZBZI5NRL5xrwq6qwCFVqtoizZFm7yILbWfSJGeBqITJZz2e0YvY
CfmpkgRC8Cfuj7jTSqq2VuvZ1U7i8F4KtGa2namd38IPCClVmehRnFXwC2CY3Dtf1SqJL/H6l/Ui
1FC5Zv7OrNjpQO/jnQvjrPJlv2lHrYEPWX4ntf8N4QEgFnuDj8D/x3nN+JW6dBRuJQ/TvnlVn+0Q
EqebhWgb4Egsty8tzhz0Q4osSreyvikVc+lS2HidlnvIUn1ktdPX5SY0BvqktgxTfu77mtOk1oy5
sWBmEGHLzWW3NnWPs6J+8pSTu0CtlYJ0XaHdtC+UEo6k9kUhCC7kLWpu3mNiDi1aJI5T94zKqMzk
A1UtnOg6vnUo5FlIk8xpgiTS0814Gj3UxLBzf1aN7E4H+XLrndnc4ygdi4RVtMFrpp2Hs+8cH1bu
sE4Mc9XeXScd4olmJrHZV+CdHFPkpb7Y0LoTzzCrG1Yy36+GeSXa2T79yVNy0OvO7HmzjqWo/u6j
PslnbxF+yAFyxHya8WCvtITS1DH4ELvT+tmMD1o3xxOCpaMv5ZFAM+VXR85h5nAGXIbcW01sVcR7
7Q3PEth50DXKEnBNiKXtBm0NY6eEd0MbhA+073/MoXFPf8s1QDFECO39z80YENFq9/hVsZrK08V7
99kjnVItCfaBw0bFooTX7oHocIhIx396sqKf9ciqumdeVbufolSnABPJ/My/WmueFvtckoJZYolo
LiJ2TO72OAlsMf6tzGKPoc50W56mP1f+YYmCZvu9Vcmib6H74kJSOxPux4aeIUf2VEiPmlCIjdOu
MDMHJwc1ubZieY25tfBktOm7H5xVOm7MV3EVdmNJ26F3p8l7y8PxqfItgqv9q0FwOt2fiv/QomlO
waIFKKTcMuPzLGLn6LTpnwAZZZUS2PE5C9o0NtXIfNlYD+wEABJWKGkzChbFxaMCPPfiw7Zp/Au/
iUjklHjR4G+lQubG3RmDCzBVz2ICVMvIrtVTD5GkSBrSUaeKjFbWQdDrDAkDGdPHlr2SHJIaU82G
CqRv0XShnjhvrxsWVZKpAm4Dp2fpJUCctn5JFmkWf3k3F/TV2TXD7X72OYiAh+zi8pend7aJLufr
KZg0O6NekGXL4DGSYXDyPYrhnRJcY7c7cTSKN2x5wSyr1rvDenSl8hksJNGIqBnZ4GxsuI57Wbdb
rFUaUcn7ZU6fpjf/qowWbkQ2LFAgC5wff3IpWU1abdn4jbWunTN8X6keCya/rjo1/36cvzSl4qXV
vV/dcRykKPN9FPU7J9TkGwoh1EfesWpApZO/kZcLle/9dv8bGwyBk/+bvvD+kjK6DNVtyf/4EIBc
NrlpwXzp8OSKQZaEFQQJQW/kzlqARDKWq+hz6DBuEBzPO1A2l6ZVlF78KuPllps1wtf4Nc3eYChH
Hf0jFubU/w+SvlYLGrVSh9UyCcn78uYVLxmtU5w3uCuBq88bP/jq8pcE4xTcAQmCRdBCQX+JitXI
OzNJYhoj0JnRVs3sCjI7DgOmYiu9RdL+ynt7jkNAy/Z0p1uRP5bXGLeqYtIlLoTGrBZaUpPHLnxu
a356P2ovX6wSxvYU8E+9uRkI6bc9igPflBK7+mKpir/GKvotqjnya5oLJFxm5QlVQEWYSP5fWL76
gh6Ch+ClAZ4Pu8X+cSjIFnt4xuM5mVNGXADUZ8P/lC3odFMVZ8CL/mxWNVkESg23RcTSDuGoFwQA
+khukE4x27Nz4j3mkOLyokZT17ghsgd0sRO/5lZGH9vwzmu5Xi/zRADsD7e2hSwEocVt5G40NVDP
KKYTNynyxvOPqlau9t1mGayL4SjICdSOMNmFgJ+PCs25W/LbTeQiwUCJrRz4Os05dR/h7/CTZ4Ii
YoBVpS/JOqLQaIyUJtMR9VbyfF1gtEBIxEEaKQUtLMtFLKYi5t5EdMjEL53XBCksKDqOB9ZKtrKQ
y7qEiru5oRO4IXlamTUFjd6oU+kURNr5cd0yPy8l199oDwg+RgjFp3Kjcuh57GDP5B/GHzB7ynCF
qqlqwd+CFBXOEv+tQuInG8FLyJ5sq4P+Iubu8SfZidu25ZiUS1lim59D1ogU2CtpUfTVMoe51VdR
XkiRKcudhJx843FQqy6UEuDIAWZhhP6TEq2M1AHpXh+PoYa7j7bS7i7A1+X81sOIITQY63SgyvXn
eiI1hFTw1fKy7QR1ZkuBk8NmFThAwU7PD1JokljmXn9xXbv3vauewpHOnKK5MJMUmZ/TEiuYDL+F
DJIMno/5QWOxN5Td/N0hoawQ5utNOspJiP3QqXv8YocQDvahOQu69+4xsbnM/FDXlF42ChtycdQs
Sg6BIPmVMJQWx8wPsWo1FiM9fyYtqwyisCDuV5NfvzCv0I3eaJM5j84f881wSk1l0rA1mvWD+JxC
owQTKWknSR7x/hgAJpnvp8Z7FOhixRqPrCwZ+Wx4Rc3SYmPzef7aY+LUnaaH3ZaGbmHnksURlkN1
iKBbi1aRL9z6ovALtIgSPXYqqLya0Sj39JPiemQXUkocfsrJETRf/0YDbmAFNxmLzi1PafVaTFKg
3wK/ywQnvBhoOGtefmyJhAZe7YuhJIMT3dZIv6HXArvefQPF7aYVej3lEeHTxBVaMEB6+ZEiF52f
4SIKhLOEWZVx5EWW/YDjGhLq2YabF+ZdH7sF6gD6eR2IliCkoCOM8e0hAXcF5XQtr+CLm+a2bB2+
tt2Pm9pHLshsvc8T8w5r57nlEQUoAEblLkzVWezU4piCZrFqm0+DKQ2CI+bKEhTDX/noX/h/hzvd
3hDiBFbpV8b2YX1f0kFuDIxJ6nXIBiigwVlABpq29rxh5ICIibhul+ntjzC24bgkDKUVa8oaQBCK
PaferNOxZcnHycIbBzNh2il5D69caXuiuzC7wKPZxt6weBP5f7lmAu7abETA4fcijPACfXex4pGo
vqw+2S5kGl25WG9LyYRkbowuYXBBDkZw8h9TQ7JySTYGMiKKF5V67v4RPDFcKGYdRjAvUNADx/of
vBSa2HY8Kakv8zdNoLIYftAlLYXjfiH1jiD9iZYmpYxTn6LLKUN6c7w7S6sLmrCCruhwq6GxzpFv
K2tS2FNsJHEiXLHaKdRv7g7LC/VTf+RlbyLUvZ3K8l2LWhjxe6B7QtWDxXuBiTMaqPGBbuIpNSdS
dkZ2olClDVO9316jp5O3NI9wyvBC0B5bnVbA14uEvG8g4DJFjwOAQxPe9TK7iyrX6toP6rZlysDj
LG4hMlM1DfZbQXQTYNQ58MZGSqtxbUtQKnJGK1hkNVGBh7rlKMjy4JJ5DID8u6IlEYcdv6m1+sDl
VUlB5rbyDT61aBwrCaPagrX/Qa6lArzkjA2lsd26Oi65TG+a96SOVnCrEC02eYwq0/GjKdMyhvIC
dWAy9dpeGLcNQd/T1p6ioy2KAIxq0nSWtNRRRmGIkXnkiZp4OCYFoexy9a2imsfCBFmvuGQjzvOf
YB5WMztrMh7oGT7KUs+Z+TZozyb3N7sYpHd4Y5+Fh2AnjqFIl2V+XeR3eGJoQ96lgor+FN/1nMw+
qkkesD/vYBT3lFYfDeHw+QecncrbtAjjq5Aq8aFKlaSCawtlX2XMS+hYlFomloNLbjrLO6VbDYfE
riE+itQw26l9dFNHCvRFdeUTWeOiUNk3YyrBH6jfmwL40liAMiFcSWyhg6f5i3JUOb3V6dukJRlj
8lQhKHnZEGzo725yYsd5oBmQLi5G2rmkPwyXmaioYVEgBCDGjyEmNXG5ZzwX80c97AZwPg0IHEHo
R4kDH/ePjYFRqJmB2F40/f32j3WqibINYOw3ZjZr9I0kFvbsCvz4L15IHFa67x3NOWAuhQxlyBX5
l5suYN3P3uD4/VLD3/nbsqyPiKjPxKCAsUG15RgInaVmBTD5QPm0m0EISfmzGz+6NC7xYVPmMWQe
uTEDEDqhGm6M3HjAPF0fQKPAEgbB+vSFRl9QWDh3VpNAc0HZ025SMytQ19THyxjN2C/TIEed8qqS
k+5ORzGA89yi1sRsIkGELvn09rSNgCyInrVtaBL75UNcT5B83pTzsM/1VFovMZ2AW+YIhqpigm6w
4FCUAk3t1jqN+YWWLOFgZK+NwzE1d6bOANK/w+vueNA7hkHpmreTmCr/eGiUEjzcth9I7HJK4mmf
qzHCguUq3lFtctp9Zvio51LUHjETkprizUM9DoOPbE8m5tfqGfDZbhVPbWM4lzAgXHlVcC2llCUH
xUfQXK8124ggvSxC/YnCS5vnNxNx2oeQOfb5xBoQzrcKrdi8XaP/R3TV4kDr2+hcA8/i4w2Ve+Pf
q4igx+9XMTc4QpnSzu0qCRn7PeOGBiAJUiZ3O1HI3n1fUK0wew3DedfXfBO5pvtZchl0fJ0fz1jO
p7X9CQA6977eyB6ueluCAY+YyGexL3cS3Yd3qks/Wh29En+PTphIsUEIr8OkFv4AiD9UH8AXBd0g
hX/L35g/oWufFUmCqV0bxP3aCst58VH+PAw4CO8KzvTWukUgtw2+rZMf3bMwu/9aAvuN6bSm28zT
MiZIli5Fmj8KwhuQTd0Z96rFIgWZBwnZCcNnrOBoDbzENHbXkiZLSQB9kr+oo3s/bJJ/x5Qc6Zag
YRNML0ytp275SuAeaX9pHSGj4lWWzfte2BOJJA7iGZh0X6kkcjH2sNqFv7C22M8HSfeVSHGBVtt8
miY2T2/3iFexVtcx9jFC05jyQlaDwOkm1fdki2IuK3ETmNQhROkJ8UGmve0z2/fvhCHg8JZ8K7ua
FZjk9iS7gjCxCQbONDh5RlKzoTm0BWPAoDSsKng/RoOKecZ8En0K9/XlKaaikKlwnOODqfyJMNOJ
N4PiCMuM2/jNGeND+lJUVQzTsEZ4K6VrPlEOpgOjxX8gf6W9Q6GwSl43tEoeFil3YWa15ZeTe+JT
MHLf8L2d6SEGk3uuqovSSi9O1rf/7u0VZqBC4zlJxWlLo8hgtlfkIdKHn0Ghuv/0ZA/GMRLPdkSA
8S6WyMeAd8MmqFh7M2nXzqAYBkbZpc0aXRdUGmU/mOCI5egmf3+bYEPQAO7qwSdAbC0oi/83ui3L
Ym24DoOQMUzGD2IyQbgq05c4MqynJa3s9Exq6n1vD1+O2RBmipVw8ldjQxes4Ea82bOscIcCCcCD
dqQ3q4IAWqjDKkf19HK6hU+kDRzzFByctlnuHJkpie51abknq64uT65r/KIfeHnT9Wh06WPR8osS
u4sU/MgTvSFBUJwSkpZDVYYCnYnOII6BVnfqYXBl4nneFbVafIQDMfJBglqfMwxWBXlP/uNSFurC
i95lXeN6Uf3ieinq1WE5GSIKZMTJksfd+HgDkAw/8TGVHka0JpJ/Vt58jC/f2sy/NBYxzqRPBTm6
KTcaavyIoS6UETN+yPOfcNNylqJbt+JPAaZOWlPpwp6J2mPgkPZyXY/xrKrLtt4zCJ5g2JV83yLl
nHVulvyLBYn8XkWRuz9bYZksLlpHUOWWOIFxfw+awVndtRdJugXV6WukSvqp3Hi1coMVkKEnIBx0
T10HMW3bMZLFedAHmuz9Gyc0kWPSIhqqvMLW5TIaZnni5bplwPrdfOLOB3upUj33n9Q0Q9xYyDDp
x4UdkwuVO3+rLOMcLZtNvaaDln7foTt1BEI5h1Ty+V73s3ZFWI4mxK1f6m2gp6OnCyF57ytmGhAY
mIY3TavvRuzcTuqVpDlVm5NeASKvmfHLYMxGsUrZgSWgb6StzR77FRa2pAo/djLKbJEwEQsJXeaI
krL1UFPVwy8wpVP51I3zPAmb4C7Vtt5CuTbMzaLgVf0IZmO6ENl0EpY1v52OaCRjuXlHJnnyLOt8
bXxebU7WHa1j6Ld1yJ/PMQDprQqH7ea63G+CftvjgJvgneaOvvwiBJHH9iO3WxxrEEHZf399y0dI
0EtIR8XbYVQtbx4fzUOMr9/z8TmXiHLEK2fJnP1n37y8saQ7xoPwuflYFH1uS2+NxTlog9QqnY/h
VqK/nD0Ml9ESuKUf7G0/QDClebY9ThWQuejTfin6LHhJ5to0U78S6GMzCMMGuH1KMMP1BcDk0wHg
JGq8cY+IbeH1nr95v4pB4gEvFZ1gizCsR3v7y94PQhFbaQX+IfLV20NwqwS+oOaRBPg0ltnEXi96
Zw9X5amINakfSn9gUkuyuvuTXVTtcDuP1gZ3Cibtl4yjE4kSlXMM6uWJaaYZLioASPRpYyGmafmj
giVPryBsnj3kbneVoh3NEoYKFzuzkZ0VegWkH1NDDSV0fe0w7xgDlYPMSmgKfklPBhSOc8vMLn3F
LpYpEdsDKqPznzfN8cxALWJuqk6Ko+I9sS7R4hsPN6ZvbDMF8af0igKMybOtRma7UfoTAwKV4Fpi
W2A8EDOcN15WLCQnTb//kZA8pNpq+m5760K+IIBvcjRg89GnyQ7+tHsS7jqWYr/Izc7BC4GQ0CE5
Zf79uWqQMcNZkC4tn2wFz10pn5aFMpkBHnBNGLuHc+6cE7I2NCTH1Ig9mtH4o83N19auxmYQyw0S
ewo0A3bYeVisPBs4Bnx1/8NrP5bVMc3XP9e27xdL8dVLwikkoQTTmBzL3ulsTbgcGUXmRLyG2qUF
zsWR7QzcQVo96Emt6EsmSOYgqf9mVHfZnHPk2FmiA5ZRB4/nZ/gTzYN/z2b4/W1gNu2ElyVz3p3B
bVuFD4nMA7/DkntL2a2OylDkmbRQWyIU/TnF4U7nG7lO4SIpmyiFKJ8WV77YRoXx6X9fMxbP3s8u
P3RSfuMaTjISJM5WMgVIFN96a2THMtKl8GqIjcneOCEW86p216to1UY9NBLSWqSQ1an2B+s1dXoU
Hmij6Gd9jQ90cqedr9ciXBP769uzv/hgG6pqMoQhAetXta7Y6m72AG0UsMz+T6dLJXvrnZLWnS/H
y+rlqg8YFKWwvENZJ4L3gQdmHXHTjKGTBx79nRQJJ1OiMlIeRAfilcdOphJSnboUkPauuupyaqqW
wPURKhgUxcK34QjxE6ydiHH7+f/oWqMl/WlKcDmb2DkZdJuopxWO2+3jMdbBjsOE5hKJ+xQakKym
HsRCQ/k4zUBYE/2vCOOrJy8C7zM+RZXRgsD3ffgDvHXZWIcfIN9Gp1CQf1JlpjklYx8DUbd+nuE/
33bHVVg2dpLVzZa1Bt+8LK+PqTNoIJEZTN5oz0hV+meM1l0b3V8TN6W2fvUUuXgxhtOojAZ6ezX8
3FFNvw/86E24EiWB5vH24SLEaja0FN/jkxb3Ju7FjIwAhxYgj7Q5VAy+L84v/Ou2k2JEmIfqFRVu
JkLgSV2G9zZEuAyNsdjkv1HWJqFjn53SMugyYjvP1s71xoeDQXrk5aWpXQiGcSd66ZOMdsAui+h4
+ZLZ52CgXLvcp1toVMbcQ4Tj5whFbbbAt85ZQiOYQPRafhqDChjl+kAu22Vnz/ji+fizX+aMwKXM
qWxAIKIQOthJqXr4mBG5Anpcqe2PTkLy1AfC8aLoC/60DYQ4fZej67p7wYtY3Zv3eRyWVWlsloC6
zmctCYoFjMUGqpKP5iubfFS6sh2Hp9BWlFEO/lnouz/gkOuXld2XS4/M2ji2fKIdW9+lOvVVlsEv
PbP/0tLFFguruvBIA47eUXP9yR3+5OdCnmKpyV5QJAjusU2ep2nw4xX8JlxTpp/vHnvGpnUmmZnI
XfSA7SXybgETbel8Fu5+llCoBadFfwtFOUxUvg4JNQdahcLhvCnkCVXwWQKZXoojhW6+L0Q3j9oy
Au+kcngH8gitdlKVJ8jVEBCqcrrkK1ay1vI0OpbfU7EB09D/o2BcQUmmkJVupEqM/YrClBhCRM6P
XJrQyEoOySESeR24hbJ00y7qffwELAsEvSTBhPN+t9iulVdd9TIrM8Gfjff3DJ1Sfk5jrClJtokv
wr0qSAdY5zOfK6AMgnK+vn2SP6lWqyYarxyFsS5YtwLTR4/cXI94YF1/aMAkmeA/ch6kZTuyDf6u
5DX6LW8RCTzaCwH2OdW/Gqj8jaL6Jd5Nr5TFqELJSgCvNnmnnx/ixh7Yyzs28jdAiT2/RucPTWtc
TsY7XK21v58+hUAU4weW8Sns9bFzshZX8KtE88lM7NmFaDejKxD5qaCRNge3GYI8wtUfbDuNiVTQ
ZNwPWrN5wamfWrQKqPr2YkkJIzEixNpMQi83RratPf/xGWNEHsefyOwmOrMTG0Y35atJYWRZ+yvv
QsP0tKNGviBxVIoDe7dQ0q4z6JhXKPGU+j2B1U5PZiNSeIy0OpYy80DradtzFx5yFYwfbwZ1uUFN
oZHJQEp7f+g0yoBeYG9dJwlq8FSJaiLrA78QF+pTuznil1UM4+Sc/+MVCzuq1GfjAkdF1L1u9Wm0
3rqdZXSxJS/a7NyxIToTlxq0SqKbWR3dEriCAt+14izwXbRd3o7lMp6YymQ6svZJPU0cv4aJBaRl
sODkziNwgAduYPSG21gS5xhga4At1ohijZD7w0cvmGkIvayXmFlNVN6/W0LfbR4qoJH/cwsmofzX
WdJO2mfZPris1DrcUuqpZJ8vS1L8Lp+E4At+IGGq5yOU3+2s8c6QSYIEmzmppYiCJAkRGTIsPn/a
BvUe+94dgCyDlHBGaME10Os2IeafAp9et+oartuhpdkDb8RRMbE2lpGrxvk8BDOLxCWvAD9XfHAp
CdKTvmusg+LVTxg+Dpp9j4tHNj7UXeKuZPLCpdeSWVGGH01ntu7VAQ7XguuvE9ReQ7TZ5AOA4hX+
nW92hO5syFKiGeyJEzNnDDSpqAJL38BYJVgF92xWHkvFFshTI50if/jLZqqa+o5IaruCm+mY0PGM
LvxhAip9QNs096dE9XE+BLjnLnStVpYn399jd/oSzsRTBKsvzfQAu9CutnOkNz0LVGTNgL09DKJQ
lZmaBFDfzI10SNkT0xsRU0Gvk1Bvkvca1q48yKUxbKfndAkCOzXU6FEBFChod4hMFVQL9I1VRPhs
RFAwnHf7HV+4byJVfaa+GcAmhC7uJA5JjqyyOT2dxGpyqJqdkioFe4JVAZRpcnKqcwnPbWsABwFG
mt/ObpT4RTnWbKHA3b0MiOrl6SLJxrVYmFVZW59+dGRNVi5WkSE+pmIZn/6Uhhl+OA+H/kGfLJ+w
Qeoq3KsMTpsAqBds+qsX0GvQ+kwjnXrxQBs+IxtYrCo7/UmUtI9r/UU0wlftHHmGu7DHI13rqGdJ
G+uqCji23/m5Ime5abtZjfP0IqFRg+//dem4enNwGzfAakSPE6WH3bCYE9QuMtezOO5kpavXCjph
JXJcNqiGqapGYG+87BXMNbHGWn3HBs4WsMGNQCRlM5Y6Z24ZF8oIHwSAyXNO/k9IAsPI3quPT496
iSruL/H8OhVwoL5yhnKX7Yy7+Qe/NNZ2F2FQKuURVdL686pkjwQZ5NNHUiA8q+YSn5hLD9a6gTwb
PVRlOlu36qUSTFYmQN5kGLPNDnnGuhvZLu5hr474BAwRp+ux3pgE+7jSJxo4+znTM5WB5dYQd3r0
DeCDon6klW3T6wUkFgl3BASlTEQIYNLBprwbZjrvmLmMn/ar09gy3gBxBijY4Omr1Is3LMwzvsyB
WMzlFL1FfMEOKy/w59HeKyDKmzwlnh/ICAUOpmcbc3gBMRh+CH6V9syKXsBpGmMMQIHyrkStLlaD
WxQBYdH4jbtrpPXPq7bkcRAOcpaAC9HoSNij+U38jUnHbcfU2APDM2ZqSA3cbSbQmRIkGN3cV8z1
w83Hmp8SAGHGFzfKlbC3f8dO2qIxbnLewulYL8Af/1uPLwjsgvRXfmmoZLjV87whWWvmTVMYed4Y
3aXDJDB29plny4b2a7kXJBVlwN5S0UE/a+bCjgQshPsU9rvXpyToN7gtpgi1paAgnU/sxE9D6U/c
BHt6mtS1pG88AkjwgjdyBv6ux7Ngj6+iQtnsrZagj296uV+l6sixTaMJ2JHENJVT5TK68BTTwgvW
TQpEstPNS0mgUepvUvoE6cYCBN77kMlfuRgYyl6sKCxZNVHcyZcmMFUuzsBfQNHn579a7K7lcA9g
+IBzcw3vYoJURZ0z4d7prO1j+bquf3a67yE5O4/qnohSmY+4k2oFfEypMCsMN6GXrIK3uzu/CUKt
LY/j6ObAoPs6T76mT3FAcBQnxxzQPAn09GKAbbixsArbGAU9HcOAbkm8q8UMk1/aqYhwle7xBNry
RXUHvFa6RUcxrY8juI/Ud51rBzG257PtgJ2zGZwZ6kkNB9amH9z12CrRh3I5l/nIeasRTYu7YcOL
hT+40cZ+fptNPUOUxTMuZKPfSlY9ZhLy/A4OBf9ygtp4dl7YbNIpI9G9P7mOdwWPQhQHVQR5wWKm
cEgtW31GhMQB94Gt3t6kQ59Z58ULp/1y54BzyGaLH8fqU/kSZGErPz707/q+X0RwB9e9ACW8oiFO
/Cbr71CrGPtcJ68DCeToCMgr5S4XhwWzw+lhXFPWhDt+X0WV4r+GqFGQbpgauqQDRBsueTXwTNfj
YQf9raD0UCvSVk6AeC3odGUYVJ4xGf014RsyRqyrNVKUhrxaBXXdRCDRhWbzwpRyjF/buomxqpcu
RT0+ite17MYO+ebkxXPk9BL0DnHx1XBvk7Wbdo/JdqwiyyTi45t8ZUi5kIUGkyAPmgTb8vkpWZR5
IzHtWx+wn/6y5diF6FRCeN0Nl3vKUe0IiQAF8rjHUiAuim0CFYzrX08Y47goVD2T/MSz8z8F7uOn
/wQf7nQLzHDbFyYkhTgFI/b7ZqlNeaDx7lgj0b7L10GTFrnxlKLRUupthCaKllqcu1xby7Ti+ore
am2d2foLoerAssJqEQA/c5uYWXQSNnVNLVXsLpEI7Ju0elzSp2zce/KcD40Ta6tVjLzPINcS/FRi
2zKV6sWIeI5zJndKrhoQY2Z70/jFCXpa2KVPIwB38nxMeTwNWJaUjrmIg1jC7cWx5Bks8oSS5ZgY
6hcQ4vKyncnIgx9NLIDUzCCUCmyMH3j2EvTlZUXdnOkCH4bei4zyfehGLgGGrnBnSPyIFw3oKs9U
3CUqDXFOjTDfg+Jr9IWczKBAIzLjkGTTZ00yvN7sZygbFqkABUbPEKnbfBJH1XpSpyV5T3Dssd4F
dOit54w3MpMfoAd47Chz+5AY//RsjOd6O/9VJo7aRTplLrxF9KWa/5UvHxTG4gYl2zfsZYwgxi1U
H5lgEB4L/bwDn8EqZUrW0o7YmSyuIml/pxnn5LUco67iGwN16Aw3a1ilbmEmVHecCeA9onmGsxtq
2T+SRgJVclKK1PqUeh83DenWKHPFNV0cgeQ90kEpt+X24jYW8tL64pmYpqx9bdV31VHp/Cup1DAZ
zhSQpeWQv5uZcEv4wygSyLmxrXHLVf8rGoXnc/wNHw4ocoim4riYMS0faQKP/TLXBumJlzzvsCSz
0DoAQEOM5DD+pe/u9QEB44DfBuvyEgFAxRlDMMiYMM6tlNKMTSVNk5zHgffWJ46k6XzH+Nh72JQm
7CZnUpO+0r+ehlfQQJUQYjjsa2lwWilT7tGad06Wm+MitEGeP5Rd4CAO2YwfYJ6jtF/Ollt0MFya
HKgzz69vS+Sj657Qm4NgTuFbU6ewHfiB1nvGX9mRf+2w5Gtl7aSDuHvpccpMyYrWEgPG72IjWQk1
sT91ozqob0MwRx0VAqEm0wzMr2g3C4SmaomDQLnOBj3t3kPvL6dWBY/h3ITrSievhLilfiWIjrkl
YnU5XXeCe5i3p0jgjxWDtVY3oXqqwSRclyDgx3OY7Xe4cd1EtDs6sTr7RrxjIMihtm5826T9xkcw
yVvGwqnxt6mzd6Xd1ScBaKyRm95wAbXWtZt9lfwnjVbazwtftOnEBhjX5N5l1/KwqnuwgErWRVE1
nyNcGf7ZYmr9znaFhCLC7KVy9k4IRUZL+d70CWqurLo/EqcjOCXKEYv4jSb13vE1dVzDudoq59Yy
usYwMVf5yGLEj3878wvM+xpv4mCXj62EXhJr825lzPjy7dkY2o7wbqf51QSmG4Xd4Xgm+TXaV0ot
o471/ANlNWoGbmva7i7J99x5ukqWidtyumvmjyso1SE4JLQxB8v0tW+sfyLPs4isidHYxjY4Z6HW
Zh6Cr5TBypO9I7T1pSiCIh0iiI//CJ+3NUWb4iiSxi+LFu7UaZ08zzehijNJ1xGe+3UFkstyxRch
YWVEeLVwwE/0o5kNZURM/RxLDEcH8QSbNY4ft4tSOocXWF3QEstYysyHcQyEgNHrL1UNBzwsT8Jy
SaEh6uQz+/RDrCDWaPAKHKQkoKD9xOAq6Y/FhyAyZPpSP6FKm7VgE5y93MOSSXTXHmZASKfsrxt3
WW0ld0OAkc9geR0liXZGIVIcEhPzQl7qZ0Z4XRjn61VuxOFPk1SAln4HWEPG00ExPe6Mji2LT/1u
UmiL542sShltX4fK0m5o1Uiw3vX+IyfKk9lzkETzpiKR5r+GqOKMzGhW3tbssFp+Z9nD2KsEMByl
XPa5ezU73H334WdBziB9Yr41abhx54zZi8E0gKWuGIRJMdZdiDsRvCrE3YxOfkvr0mAPM0Uaj0/C
u+AcaokSqlSuSlNRo3+uNtrXzTrYoKNteNdyQCvjezLfSxs2oNT4IIvNSSN3mgWcgQNLPL+oJMEi
ObZwD7fpOrB7aCUyX0dO6nbiOn8ELrXogz0mmanDzVpm6k6lrfoDMYUVgB7lviNmUa4V5Vk5hdkE
Pgim3q/SRdawpq4sWXgeZwELVY25O1g5PSi3O2xrNynCYp+WM06TNWCaGrxQhXmwVErlO/alshQZ
/0vlqHBCuOBJos8tLdKn0rBaBXKrLPMWj9LjEnjYt5xCk1cWkDqsTjMf/rEsO5s8mCh99rC2QjQV
EMPmdkSi1rnoVifqTvlKL3mxL3/WHUMJtBdohqp8C7VlXuq5OgOGY1JbnQlhzvmfNP5NLeTviA0Q
D0ozGyz0FHCjIjWSbqJ7U1nFQXRiRYmC8X2uAk+mpTEu7pMjmtTyRTZ881r4318gYKVFlIVx4Y2M
hxJzP+nXm5c85dbmFF07nM+Tz3mzzbCPFqipjDy7ptacX+qOmLCPZi9URk0ryDq7o+zXh6Jf2ZcA
9BYmuShvtwwiQdayzBkRnQWIXkpwlPGJTObVNQlXSDbllRChNe/TAbofXIpWIAooTwRxwJmy4yrb
pAtRRrJs80pIDgeZnvSmUk8l7UHAgzvMhVSNdI4XraoxmU+Nreuzze0ky0IasJK1OBstqEXUbyKf
7mpmJhaYPV2YKRGEWvsm9X6yD2BNQFVUePvCl4WIx8LREj8BZEpkc9oXHdt+iIoEIBlSCbTJj6/0
wuf7BbURyL2F5cuVYfiNQKhoZqTR/XBCB5boUWtH75tKS68iF3WJlTp/K4AvAndp+n8eiE08XBAK
xVP+TnnNVLzIqdJy1NDyT0T4DOm4qqA3exUzrz7kiGcTY9czwV2wjZDhZCFVSYP3MlPYDQu61dMe
0jBJaNfr2W0FRogHX3B53PineY6yrEVzNhboQA9P+YMCROwAT8ZcxkA/gbsrstqdWT0yMiHBksP7
Zj5dPAJTjKbw0EHJGKja91PxbwM0V8H/ph16eiRWCYzyX0My3nfxSczbWex3YtQx6tfhMA2zuMJ4
b5aWXuLUGZYjA3RIiAOTGhmZ8IA0or8v+Sw5tDOwswWam3l6O+pqpSlmkzhnpA+7JOpLw5dHZYq6
hzdSRUj9LXp+rY/BramlEJWFrxmjSiuNhRxcYQjsogqTk2fUNL3M0/NXluPHEaOSXk8zPlA04FyH
OjuIIOtpyLft/5YJfQX2W+sAoijCVv+KIwTYodbjug0LtZEyoxfENDpITIA+aJR3WXkAp1elHfLK
xqGjgqD2CIQAxmlI2Ohl3nFW3TOChby6msdVaBsJHxReGpsRRhwSWJ34s4Zjq9NjA53sp89qIbBJ
4fVmNKVDY43HvWX0zkJG7dmNkB5Y4HSeZsb8aNm4GirzJXMAUtOxT/uNVt1zd01RgLffHY0x8L0b
VpiUg3ggldT+plAHs/MHdsNyDSajWtmkDSw9WvOS7IatV2y7W0CsktN1g5ZQFSi6mmBzCnjvlBlc
jIxg/lmAfasAmguUUd8S2qB8kPei2Of/B9bdL5bvmauSlXwDpMHWY+wOxegz9CpzOs4hiiZPAuu2
SS18OK+tiXS8pqMNDzUmHPtXPR8EJFPd0wWhkXkr2fNoWkobCX0xzqgW7TElYM3eYwFFRlc0vcED
o4TAbyPoMX74mfHUXTUIb/VzgMChXjI3DelGkVrPwJVtBHCsqyHag231L9rbBsKufOJmpmS7Yf30
dnTTn8+FOAFQzuGFzMySI+vZa2btegRHo/P+5dgXt3kJoHZVe+n4XvZlId1Lo47uznd7P+V8I0I3
TyVrO1mRobwWTT9b+wylFEl6cIpiA52jBATxYUFcW9KBp4ztGs+YAetyfQkqua4z9DrvGBF/MQOM
LK9HA3yC3bRB3LIAQlJC7Px53dlPfCYh1UFPNbEMIITUHUnLh58bsH/tNagh/ecAXbzKSqi4rh6T
AlZB0JfXZnIzKZPbPKzgG8HLT0O0LPPjHIAFD+Uaec86NolLUUstWlxf/Kys+wpVJcZEdzHDzfe4
32+SN+7Cb7YxdlX+nqIarB0uih2ElZ5I3C8IcL/5NImv2tkJQUmcUx96Yjfsl7rSdP++fp4rs4rp
OkBolY29qs3UpelJu+gmICtf+MjZRETUVm2Mi5kQbsIyezBg2H2f4ZLMmQNwm/lRDr8Ybfwfz6bs
osWOfjo6YZwyN98oSQZGnyROyEP4l0A3sXm2OAf5ZF4IelskYSQZi2QCSL/2BdopfjJoKh1sg5nI
KcIzVu3Q13/z4nfRcAu1qnfnGyJkul+Y4WXLUlYpowMs2NP5af2PcPS+E63J/7ckPpfV4bCtsm3T
slj/8E48ypDdTM6/Agok99aYRtjHJIYSnvXFJjEUopBq7bGfiphHKHaqeDw1pks2i2zSsubrzDKs
HlTqfRVmK8gVzzOIqc1tmFtbLVkaMQUwrruNVorv8WtF/fKmLCXCj9QqhbmmRQoDxCX/AiroH0AQ
c++gRfB6f5xaXR+OWcAMUcuIw8RrTCP/3d20l5Rq5bGA88xruaYkt17ar3M1z5KxrjOkVKmYCa6L
Q0K3z6hOZclM1FuEH9O7WMtwemvRjnw+ch6LTcvLBKQIvEMWvAReltF8TYO3tT9g8IzkizNKLw4q
RkwKLyw3C6A65VFBc1pFwz7auMHElUgAM8fIHx3u94LyA/1fGgDuI2iSu09b3rXnip5p/O5CZ4QZ
cJVkHa01EVs2EzvObskQh1WWs5AC2uAuqlQMYxtxSLXy0guW+uzRv5yMSVFmqJGnK66gFx6nDT/y
eeWV/3ZtCfFU7tC7Xc8wxR4JBdx1sipho7555AgxgY4/evvEdax2YSoSHtHcmy8LrSVnHbcNFj85
rNMyjdXYADZqiS/Q7PLUklBdsHC+C0nl9C2LMnkJJVr2hMBmTWM+YVjjoj7fVqUBa7YMtOi8UC4x
IGbUEtfk6OAvf8yXoAWw69lI5U07VdhZCT1e6dO3EvKl+tOHW4EuTnEUjeVZ76RKiqX46WWGAMLG
f6puyBKeC4QvXaGQG/Rafu1FKJ3tmyfuIC4AvWB0oi62Gwq7+CJ73AKABT+p5GkbMYuwcoUblVvt
27brdwa0ht1i0gH0LJNqm5SOMg2CFhDjXofM46g0T62NmubivoDvAUIXmHETx4KANdD50R9dLopj
JRTzeS1hLH6/xYIZkuhHcuSK75mfaS8u0+r1++43pAfRewCkkQjYnGqeCr7wjlOYHJL2LpXW3bZJ
Gz1nRYNGPrBC8vQ0k/LAfNc8hcOKV2nttNYXsauQgjkE4idvDA8WcrpifDX92LZUPivi3CNhnZB0
4VwWO0S+mgY9m4qEgSREPF9LzYNoaN4JdK/OxHSACfsXOG4+mEuXn49LnsCCcTavOeSyKJqoLglD
D/eqayudUliEuisLKKpWvANCwOlCQot6GffxVdp2MrybnfigFbROoEdovtDph7CPPTXW2dwsth0w
iQU02rKOX3yogbo2iS6qs6f87zQwn/sAQifLRkEC9Q0C9pE1PN6F/4Zrh4V3Vp2+rT9KFVfZ/sJs
X6FaVaiiy35rD7ACmP1f/IHYUVSmMjadWfiA/n7KyT6bUNnh3Yx3Y6tD49M3u8sZA8e2G1sWnlMj
VJay4PtzMAgulD+Ak4mCkD8I1igRv3LIvYuJmp/8AwP261+FUAXq6tVMLEiHK2Ys7LuLGPqYZ1nG
6UlX1fMhwwS6bFl9yuEdOmXxNcR79p19nSc5ZAvDD/k5oOr1lrPwBh+ckF7yANI50rewoKuaBCPg
y3xLsfHd7pirdHwtz6jXLxYGgo0vNGzqA4osqNTAiXEJFDSSTH++OY/fySWDNp1t7rkYcQbTAb7s
US3ZKIdt349wIzQRB27DVWr7bMViXqcr4R3lnKfANiYZ6D0+F3DpaSPv8anuFSHjL/cP/wCEKE19
nmlhjb/Cos2EOLRkCIO6MuFN13Y/z56i3o9rbKs4+P62NU8sAzwPdwhD00deZA3jmDQHFQSQ9SbE
qriPz1Er4tHDdwje2PdCuDsHeKFoAR3K2fsFKnxKJ/Al9+ZmLzdZZ5jgq0yLBVhhERGkRPwsApMO
UjpYzulGo3A5O1Kzue6NZ3kZFdgIho6mvWR2K8ew0cVrlMI1GK1ms0t5Gj4tEWTF56k4aNP3/76K
ZAQobj2+x4pOLYBlhPFeKNJB1SP4i3Lsmcyo0r1e0OBqFzSUVk8jEzg3b8ZDQV9qNQ1AINBg7Uky
WqiBc7vu4d4cUuROP87RccVI2SMk7PVKIVHD5QAw3nZrsK51lNNOV9GR3STs5NKseaIMNNPTDIZR
bUGcQ1ZfNkBNEUlxhOKn3/yeHji+695wqImKYubqUyelTJ/a1m/EniB2OZKf/M8vNRTIn6hYMVXu
WamK6WnhF2SOrp/V6anbYIU3AEStd9wVP7Bfq5oVtBiaUBzdbBC+D8hxnXHWJstnvzvs++hmpc5/
lZg7dEb0MDE5sYCtStlwXv/5OWSnE/UIsLdcyjKiVCkyY9F3j8SHE/zvVyOiaGMJoNJ0Qgo0RQic
g73lGbb1IgANJlHYdQs+TW3/m3gdrEKFod/5R9U2MoAXmIVcjUTb+5f2DKuMNLfIbScfZoxf5LE9
bhW7tXjESlx2vD4Zw5P+CcIUSnvrp3Gl88Mi+qO5BYcxaauWtSPTEZJBwHAuabDpNLHwjQVaRyqX
SWAhFCo7jQKjpB7CWnBjyB+dstSxmrvvYKJ3zktBedRrG79/98ICAbAyja7A+eOsbrnykV5fo+Cg
iFqz/ADMjsp9GTfXb8ARrqzAjyoXk98Wr+Fnumaf1gyI1Qwd7usQxz/MJeybQ+heHLAnpS+iw9Fo
u5VcmzNIgdWpFowv1skkbHsH9b/SgIBkF15HCXejCO1bjw+cpBVyabRNSloo2NWReYypEAggkA4k
jy5kMfj5mUx7jwfHPvSCDKRIe+kJPk/lgH7LaMxyvtLhwVd7x9eOCkQ8lsDDxxbs0kowuZnPUrW9
ieosIGczdQQLDfj9PMaojoUf0PJ+ukReWUUJ2sK2v9VpgCCLADd1KyEQTllCx6vyu6XWIoMUB5pI
PB/fznX7VnIRLHGxPU3uXYAjwbL0boBlBK7iyQoIqudTabvZBMQbfp+E6tVv+hDczQjoIeJHvj9w
6q+QvaGaw/+5qAi1B+pHnTiNaO1zGMTfa5JYM3xnELD25HRXO5F1pu/6KmiVDEqC6V2WeywP2KP7
szLYxGDJStocFMup+HFK14DcaoSJZUprg1/pY9XvxcgFAOrevX3XRqP/8zd7YCB9Z7qOmf2CaUpw
tfmYyS3CByaENFabdJzTLJd8l80QvnzptPoNm1/FjR/1xGURm5j9T7Ed5/yOsrgyzKUVszcQab3r
idDYiLBFYE/AZEepuNG0goxvF9wL/wYw3ydYR4O/jlkFKwCNnrrtGfMpEIERfF4PXPUPYeef2mZc
9L+Op3hA+VMEp0B22sRMhX1sWGFgf5KyKkiz0PNEjIKqXCYprq9SJScWhjL9GV22usuZg1HPyUic
pXck445sha+xAOUSNbCUrk3VPPyWOKSQNNZBjSOluKsmXRSN+G0FOlqHUShnpZTZdcLsFDTUFo0X
675qKg8eX/BCvULpb3+h6a/NPXetax7KhyigdokjGhj0VEXxp98jh7t0VV9N+eva37UC1UKcsuxI
i6JNBv0+bt4Nk8i/soo0DGJM2XdmmGGWXPDKs8vhFFK3Wvvjn0XBJ7OsGQp5/SkM5Vg04/teLsy9
lZi0uUCmJAbSjPqrhfmafMw+XQPYD9pBJY56QBQi18qoFmj5e0tJhlpp/RobZpF7f7OzUVwcjZrG
cjFCKg1yWUVhh4TJpV1/oOmzCwQTtil9RugUaGQqxyhcHMuiLsBEiyGn2y+PYe5b31X96ph3Aj6n
tiJpsQ/eDr9JU7fNXg9LMKQlA1zUKo6a87PVvrNmK1x1BVOPI2XFVfFaZw6vRJR8V/WfLkq5380L
t5lN/+h+uiAwgle7m8jfB4qpbfwEeivoKtq7j7eAqq5wTW/ShId39RQHTkVs0uWb6QHz8VC8pT3k
dXGZHKn+yJ+h3IIu82lMXwePEqen6otFyLob8ge1JCMe16qXvPIWftcXZ31L+TbLaPhnnMzPUAWQ
tf/QlbcutfiSkkK1SrNmPxorAeinozCfaTx/217nRLpbmmukr09Plcz9ahcczPss0K2cgsH2WC6b
r5qGRcqd/Ih4Qfnodg+XtpvTIYdEJcrucydIYSJcLnk+CbHO2tiGVytXhW4DQvHDMt2cH+4CCyYP
J2oWD7AvBMt6cAUfmp/s0f5EgiuT/obtgJVkupwaJ08jzg7b+krQete7VlxFnnL81xyZon5tzYij
p57xwiM+kZxS6xd+59gsVrzfaqLSfEsweyek2QAX94z2W7DddbX1NUonDIE9c/0b3lt+ATdRaUWu
SYuskk13Els4M8LZadvuT1lRwrzeXxXfG2PAj7cCvwx5yGoLWeex7Af9/7o6c1V8GyuaI/VdZc+D
SlJzb2w9niwwEdFlmtWoN3Wl0kCI3f5g3cQZZopGQ8GAVxxklJ/hW2D+Pya/6PKpHe1Pr3xcYSpW
KTUCmc7Y2bZZEl2ncWjmDFhgxQxJchkZF9lew3PNDJ8CiuJA3HDFCYt3EG+4nEn7pKKSLgssEvwf
PsSlo6MTX8uL+9qmtmier+EJBtieu1hvjW27DPRG+79s21DU0T7i2UlfrnwLls29fs00S4EoQOzG
3pDp5DCbpaS8yxfSjwlA9PKDT0sXyA2kk9EAh0GJKdSYGinElEYDeLzppI0BLJtvtqy9EdeWoz4T
AdzC0YmFOe2bp50BPYEO6PT+JlDI/6OEWfGBzLUZbaQCgKSMn0RQqow9jaa5skfY5FTc9ofnXoYJ
kd1OsoVLO1fSmHLKobpS+bB2Qk+Cbpq/a2MmG9isQgX3XHLZJO8TqtiCDEs4qBVqvSPDjJaPef+x
DggnSyUacbbZsHvBpCngLS9gTTGO4kirvvL6uQGv0Jv2DlO60DjF9ZqX+coxLrkFnGIsc0RPIKh0
NQT7cSg0mKE14QSYPRv99h7Uczgd3lh9ZFWGLpxc0AoSy0OCXAWS9WdW7cjrDmcX+kbAmkWHwQdz
0PpuMLE/e98PAIQh2z8NhLEK7nlVrgUju0P16C4sc5pzMs2Esgx+bgTRX1v0xYibOqpO4uhfgbAi
Bac8sS4PRcv4lt/CtQsEowSAZFs3RsHmAAvjSpmdq7x1ZkSZimsXPWqiLrZ1TDxO2sYfw5RifPMG
NHqcqqfUr232F0Ea0f+cLNka1YikioqdJ6/NwH8fpMwkvaeZZSu1Vx6vjRt+BI7as5U6B/HribZ4
zUMIVb6VQl+fKeM49CdFGaM/hepd8LvBVSc6jjDgGVj1/4s5L/ABIOPNIARfPEuuR55/3+1BCujx
mZHeeEhmV0PwEevle3gZM9fXRsXx+o5rjIVZ4JYW4+etA9/nTSATiQNpHGseprXq+J2gv0Qi0cJt
hsOqdoCGigWhy/qMS4emeAUjljWmgUlU22oyVh/RCp/kaV+llyzU7KeXUM+FfxZbDGQbtFxXSw4f
3ea5RpWdmur3Pd/y6ixC5rihdSRx7slf/NydiRhJhwIuQGo1Ab/bgALuXrj7n7pfvIYlUEhFRvlO
pU3rorcOyYXXkYo6XVqn7vZ99ilXxg7c5zNhuSCW4COlAHSj4OD0dEuORXDzdYAO/XqiRV4ofWmU
FQ4CVgDnPjIpYBwrIwbo+HruVs4KlM1qqL7OClU6iGqwvyL7WhyvcSTYIpmrPOjr9CWe2HwFwAex
k0ZKpcg0h0+7QWECf6XqMmWPe3KQvw7qtwfuo2yl7bn3pEXFkKZOPC9QtPaq14voMiKQybMSrzj1
QynRxbHpoe8yCekzJYPw11fGnnEeDKTIhgcJHVru454tZg1180ERgwo7naEgbJzDB1mS7EWGlXwr
dFiK4p1NoKUzJVRNp9jYecFiF0ans878GZqcsBQymeNezariXvtK++5b64WlaVkxZYAm9U9/UKs5
/gTCYgq2KlCVO3mfjETy/hcCv7kI8fEBT/ls3BSnTQqR8iwxBH669xE4uvsnqwdtm4cjdOwc1NDB
4dyftZeNVPfIWxQE7puIAtQtVNWVrWbBI1hd4Dvob8OtymWT6/ERozBSSj1F2NfpUPfjzJMVNyp7
mUmIFBlUD6fytEFvEiXD57iyI071fINrXBuaghDBhwDauc9SEqQFG2BxRuadjBf7KkLyV61FSKch
CXb2CPKTUAzLJoleKAadfcHW7joNEBR4K3QvBHPjhlOQDt9TPskMBHcf6fnGdj2dsm87VfpxgzAL
NDe6AoQ4YggGL4tWDOu5KEmmdwkt4BHby2Ieolqzj1mBKoTv2BX+fq+mJ4jfSX62eoTuKrBcTPHD
gZsw+CDyUeOyhs7//n+rfFF5M2j8SOdkSC6RC1PzcGM9hpsgQMlWem0uIYYG5LK1Gt2XU7fvldiB
vaRo+U0UcjwvzYMkLkECXPFz/9qgkDYq8YRUUIJplWI3zPr+w990EtPMTucOFMcW11XViGVaitc9
E6Iyx9gOjB39CucMCxh/SwqibDi7WRIJCsNxTBlz4gAuTHd/bc5VHqOPtiLujm62YRO7HETlERYo
ko5ww1dSbIYZWT7+Gm/1BxHVCNJH8gIXnv12P10x3Vu+hHmi28qlJRV8QhE/5vXdTcIJuwGiJbyP
nVBjybpyJuqV1a4Fh2GvyNJ7XwA8o4BLTNJOlVLDv8szL7w+bLkOWYCnc5968FfDTf6xfv6zDUnA
MtAnGEx/HYFn5hcWUCwyeCy9fvEtviZET6/Ukizeq1upcCoSPdO17tIdfkjZKETJtnii2c5f7Pxm
OMVkK0tBTIDXMxqRJIpYSzzxX2YB1zNscyW8P2ho6XHIlRvTwkl2/WwZMPWbMhmb8nTRWJjyFZQY
dgbQMYBC5yoXItgcqt2qExJKuory1xAl+eYAcVNIjpUqXTdoNIhv7ec/MmiC6rYbQ+T8Zqg+JEvJ
s5jlBFBrg0h6D5cKpF005jM/VBvqwcLfFOUW/975jR+G/YGnwtRPuvDLVWyjuNlP9lB88QE7Y/rl
eMqfyq6O18UBJ9EN7IlLH8jKFkTc49Jt1xAU6oP9RjDdGX/nY72jY87OvbahCGKL8XpR2cpQJKHM
RJnLwBm5sdurv0TbYX/EtmpIWf+Tbk4HsVQ4+Vkx6rMezjUXZYELWu1BLiUkiFSyBPaLyiJOMdWt
QvQQExPbV/lehlcub0BtiJ2wkgp2jqluPniizB0qIQCvLE8yyU0yhLKf/TC8ZNRJsPgSNaCctTWO
5INsfEaGhL0sPuLuQyHL2P/7Rp14Bi+nBsWRULXrEkF1BVHjDrUxJiEs5m3+ooB/ZLowlXIy0d6N
+NVtfJJRnvxVtoz4U5XMEF7ZjqNaWgmjGuf2Rdxrj4uHzBhFtpIh+mMJZhOHBB4cMpXJqG5jOxuA
M2HW0Fj87D0/sFE8uq9EuOPRDJyX+DsIqleSpNtIyvIvW/yhgAY9158fyc5C+C2aUYgA+RugY0tq
jbZ7F09vmClREPYI/ZzTEFl/DybfQd0c17ewxfYU1SIqe7g23ddDlHte1h4dKb1odgiw3OPxBvbv
z0nH7Cft8VWPnarmCDSkgfnziKqEMORqDCQCAhl0P2b1pAGCaFiezUR5UM8B20w8GLlP1izr+rz8
LE2HADtpINYFAYYlxlvpzm7QPrxBEEBnuUbbUYII1GpbaKvbgmbj7HSj9Rniz+Z1G1xCM33MmCLK
9a03A3hYcS3qjaM4aoemAuqbBC2FmCgJv9iwFv009UwdNphb1nBC2wLBe5Zi9+shJYeb5TfWVIIK
rnoICkcXZpkuASJRFKIBDygSX+c0hjFWE550laAG/tEzJTMFqI0zMMJf/U3uMJ73SAhXexZg6ZxQ
x2Xp8LfGJO3L/48IPPNxbCdWQdp7We2R406Zvo3RYPYHTBeLHNztafbBdmkH5PhgFWtnTI6CmGW1
3g2tPQJROFv5Y32Z5xyn0I58IZ/4QKa2LlyKzVf4Vwg5+9phj4JZeK2CXqhMWhtJRoYVJyIqfvyz
C4dgIDbj+VlyX61YgjpntHdQnc6Gf0rCNDxKuaMmw87EZYz2Q0mwNwxT41AkXoj8AQvGBEx9AjG2
2MFUqbsuya3P1oFrZ/Q+odK9dGYTHy8snZl4LUfsW/AnxvuUqEtxcnJvaoz84sBFM4nr27RfkLQF
LdT41J7nhbIMcDHZ9i7hP7SACCyTFlvwRL/+hx1TIZqAUDUEpn3D0p+6fSzBx+UsVvyaaBtYoQj+
e6uLxv0mZv8BlqhreY5fivhIru7JdeeA9+ZMGUynpTqI9FzQdc71jOcrV80ySBGEHQpTNg+7FyWh
4QXIYQAbsRDDxWGzYGJ10Bkh5pkLMqeNHku2saTL+RPYNSiLaWK9UDVaARWeIYWnZDueoRdJGpsf
RtUiJP6R/lK3piNSkd6f2uA7SN6HX0iclJdOXMpS/k5yxxy7NIdiBiSSdsFw1UaUAVU3YRFEaFB5
h5/L+Oapqic61j0OEy0YEdTpt9vQrwv0KutMUZUT5pNxWqxyspKapJT/MwS1n4WF/g1gMU6IaBra
nmjWvBbS6OPqcOxmU5OJBd1jfkJ8JBzwmKw0JtPaA3dy5K5HpN5OgtULCRcfEOj/dB8anaRJEftH
4rBcyKH5Smrkzakyvg4+mCks780gJT66XPK9s6eHI5m6mKWWjMEubJGJFt9uFwHzc+AqMnF6R6P0
faMIMFaXqKJzEQmnclNDljJuMzOje5oBXezwXWYbuiA3JaARmzMb7vyKroUEjxGtwLbnmfznYTkR
xw9pc9ii5ayvnUNwbzececa4DLJGwYVJ2RZFRkXZMMIy7doeBBnFDi1wkNAUphBZu78cgdmY5dsA
+aDEQtA2INYR/IWiI38XTE4VnoHx4zDFj7rO3LGFmzTNuI9GByLfseS0xhjVCFgUjz6nMRd0iz3x
cd401rRfa8BwegLWJXlAKzk2qZTEjIX+lPrzdVYaJL/LpdvQkLtDGgXNFaL6n8r7OWSsX9/QUHWz
1f9iL0I5ZgxJgtQe5U8b2yGv1MUt/S62g2K/wOUc4yvkSg49/z4JKMOg2LPX2p5+1c3ZBmBH4mlk
bAPS8RipSROtE7jeeIzrqgGeTZ27vuBZx7IiQ44jaSo9Ql8bGkL8Qn7OslZklIXEs+ktuqNsQLpw
4P7vg+hZI0wL6oU+2r3y0AMnKemo0vkD1XDYTJ3t8SOFZvVLZ9g+7FPh5MgUOnKjvBzfDoTC6LdH
MNdJnArW6kyyiRrjsWutGq9WOQjoaIgcdgIcglxwjkAdEJBJS7P1WzMZybmu6msB1WD6iMwqgX82
T5OhMhrEWA1B4RT32mvF7n8rU3jr7BwrRFEy51OIlPPHbAR9z+xjrumk0afCzWKt5jEJqWcP7cIW
VOGxUGfqspf00bge3lU57WdRh7s3Dnon2410xUcgg1Vqu87RWMTpC4KQTGIF3aZK+j1QQZZ8lvz9
YVLvMR82oT0VnJAMnAJVjH3JPiC+nJyj3FOmGXw/rmnOnX2GDzcWCtZjIrg8IP++foA3eSyjmI3A
d2kSmv5tnM8VrG8mLPNVWaqJvBT2BsrY+4DhPBU52V+NAPZCxj6Tscod07Sr5NB88+NuQ+D7J9kA
vCPbT03ZsnD/RPPOFqg38ruoQ93UNS2TqP4tHrAbSsWqGbZqEJtaUwtR9x/BIDaktltaDpZWcufa
IGHlX9ij+/en6fhOOXIn0s0sN5erl3mQvJfVOBErLWKcuQCcIDWaXJpsKsk6mWGyMP75leLTOY8q
nfxmU3cVX5IG9fC2zJZ5PJuDOxq2uNOua/3pbZwV5lWQacpWvYBDFhevUGNnFOIG56qdl8sBzArF
WJ1lxuV6B3dSVMbCj3qZ3GzgWlzcGqyqq9u4z9Onbm2idho2PDwuolco0fpkxBSU7hZnKCyIeQJo
msylCHVSdMIDZ9xZBva/jbP0odqC26pYTXozQdOGBvjeRKLtzrwn01L7RoVrOTux3X6DLauF5G6L
9jd5gNi41MHHHt3o2DjJRzojR77tNv9GL1U0WmoHataroieHYzo56SAViznbKVYPOw8cC9jPqcSE
wjxTf8OWT7M5ussHpv1yYgdA/mVLJfZFbaHs9ujDuAxtjE1eB9rD7Wez/AJBfmgWjBREQM7T4UGz
tO+01dEvKHLFEyoKgrzbeZBW2erBED5zgcfgaxjnzgXf0+gEvDC0U5DiQo2WggXXkCvQOzJZmeEb
nRsc8K7XdGeRbTaj0K3PkHtVhr4ojtZhvCWBQnlTzgxfrgJXBAOLMFeYBbKSe7/Ojk7aiYufyypE
yJUZaLJ5U3+BC+GwvbImj5kga0VnyP49hWQiZ1OXtvBO+0d/5jjP7aAhfv3CUzB6nlMQQ1hQNKxi
B/3fYGApnyhHdqc6E6iuHr+wGS1lPyxg85XSLZDsj4Qsyh8Dh4Opv2miENkD9CO+rY2WzD+dRSbR
bi3aPY64mFHa4DeImtthwYS9rGEztMhekgMo+wy12zweYolqZzhkK3FRE4MoTnoJgAIr/WHaB2Np
oWuSH7UETrS+jcii8f+GuFtGBsVqIpae11ZrGJkCTJ95gaaHq0U2+HlS9/kEHtz29KllGl5IpBFl
PSX1piVXAgmO7jbtespY60QCHlOtq2OJvpWYORokL3Hzj4U9tR/jMAo14kSOfq3HM4FAgaC+ebk/
l+pFKWkPBXWlswGYKxHH1iJ0GpdIQuLJ6I0+EYKigd/+zSTOXMRKsWB9rUuj6LADyjaO0e05rg1i
r3zmlZNUm7aT/Q+oU7/fGvBRD/PX1kgSeml8hwhpw2YfY4wsDGi+ahG6x1OOox+EgvP4YoSTA+kV
+sIQy1d6sJ0otL4h1zIuGAn3G8TnjQWT/a+Onbji94+0/zbPzA3NhfrO5TrMtjwC0iR3uJogp00O
mks1Kr2G/j6QrWW2eSVaL2CzwX4hRVxhIzrozUTMhpUxABrFHOf3c4dHoTheVi4EUqOisiYjrn46
p0TmSIfvoXvGX8AYAyWuUa5Oy414P0RFWIy/AjyFpizbpDTigVFJfptzE+HEcG4HFG0XXFRRd7cp
c8BAzikkSoqMO56UbB0peOcZqXgFOn/EATdITYr5u/GQR9f+jIINBgAYPxQxeQCxhE/VWHhNMaaJ
vUgsoWi7xHabs4r/zTQ73O7f/8I17zRIIRFixqhp3U/nEHlWQegCKqK3Mr0TgnPccfgXLUqgak+Z
ZLnep0OoOk9yy7vgDA1t1I1+us7c6cDZoYUzvBwKkNa2W1nB0Guc5G477HJZHUY43CTCBAdtE8Tz
GF81tVxTtN9Y0KvYfA3vTFAg9hGmsDErrMxkY1LAl4fz4uPHWadhEDllF3+xoNEFjaibGF2xBtJ0
gI72tuzW9rk95Pnrg0e17//2M69dXG5UceJ7BiCqOpXYm8R8xE60PKGUmPgEqrtmZtnB4MpThojw
SVCaAgR7qSUIbLjzW8Iw8l2gykBfV2RXdFdnxcbwYsgEwSieBc6fv2qoUXztGqZwDhg8ELIl6SR+
/1p+GVoVsvsLiKwi1J+HMosq718M7XOYqKqbCDi7UX+84nky9J2sKQm9RmSmF0AKHPZXV8ja4gTq
pofy0deLlx80Ys7+4MrNNahXQwrSHhcXPjOpMsuJpE+lixFfFU7/v32hOp3z4o5XWeHAeht/MMZm
dkMlJJmFPd53Dvi/AASJ4XHw/+aryimSj7b63hAxwvnOQ0E+eb4VPVs0ItPHC4Wa5gZ67M0KxZA/
BICXVaiV8gxLEcJNUQ5x4h7lMqsMuL+3kZwFXZWfF5jdGRvQ5vXBArhKI/BfjGWcSWpw9tCjPTEg
34PtqAbNO0NwCgRoh4yDqweQn/2A2yFAGgolZoLl/UDnTds10mqbTb/8VZ2Rxaqe6z/8SbvOHD69
V4ABfDasBxScVwyFGLg7gVnOhFz6zgTvPnK8SnE4TqCvxQULvE/WlHMsKsqiuYWGAEtm40ooWXGz
9HcDISr3D9axAyzoGcYnjjfiimbB6DJoje3pT5ctoYdtKMlaoawV/oNklW01FFgt7ArT8QTcCj3L
I9KYnwY31Nz/3dAdgmsV/TZ4g8+YGYC03h4I7HF+Lkb661hT99MuGOJoAhLXb5/ewOqi4vXGTtc/
5sJziysS4ONtw8Wi3o2gWbhk330eBn1Fb4+BTSTRcpK+tL6YfWiFdJaIdDw9SU16OC+BVg+m+FSv
v/2a8mcBXZ+txyusDMJQWcmyj6e622lMInirqmxgPNM5BcTwL+ls/xm6CxzF5gVMZr5wzjT/p2HB
1x1btiMiCCJ5RQIuyie5wUrkpueVSATdw1DlVXfpYMdqEz48eYpXbeQkXKeoqb7Eq40k3F4QE0DM
dpyEkvwHRunZ6/W/PdYSxmIBLQQoZis7xU/7JNlx1QBvoufEwSULmercVPG8c2dc+cFMYvFO5cTr
xc12XZBEv0C2k+cbRNqvZzruVZxpsBfXoBlDISP5BPOA5VwmRctATWB7t9PA/U1D/X6HtoiKSI53
TFXGYjBAdhaWuHA+R8LN0H+c9IU0sa97nR6dmqHZX/YICHvbz5zA86DfC7m6xbzp/wD4EeTbeOhd
BxVVI/SlxBq4bK7kEHiE3hkXPNyDUfJ4rh1jqvnAfmAJ+qebNbZ+T4csV1Y/vMkIMPgiJFhwtJcl
YBtAkU9F3sYBx8wVXRbRMk/Q5VLye062jPYb+kGIJNY2ry59vp441xseSMlPWRrQOVUWNvUNjMnu
bfcYa371STcMvotfx9kJ2y6Sz2AsorwzhAw0aJ+dnTvoS5pMaGWBl+FxojT+9azWmkMD6WhibMGH
/4BWSyIU8sqa+yu9POK4enYnSdCWGUizC4kxOt4Fpzi5PFNlrh41g+u6pNa+yT6qUaavvofzC+xR
INw18DEA/+7LRIW+LtzIBBDNxRk4z4OfVzZUa0qmJyM02BgP/7n4Iy7RqkLZuv1WDJ6of85Dp1xs
ZmXZ0k02kqcKwA7NTu/LS9ziaR9zewd6g5cx+i4/lvMYPjCVQX6FC6JCuc1qy2Dl0/6vc3e9VUpl
jAz291NXXX8skLjOMveoiphA5CFMwEcyKqZghx/ImPoL27gQoa4A0fFRMWcdzyFUqtWYUCCn4XLT
mpUT0DzhXtMxjeguHGzkJ5TwGeC/+WtsJc85ppD1prGzXiBIEc0yC4M6yK7YMhAmGHJ9mFGbF/dy
I38CA153zMRsNiEw62ynZXNmhZCRPgtOp7tOZU8qWo9Des6B3S9VN6Ar4gyXkSkhkJZXBhwAUV/8
Z4HE/aRpTqr2giU2/XFnbPBJj0ERbQEDnfMTHqaFklXx7Go+tuNeavRnw58m2HJ2PXipUyVOCPBb
CEzig2Qyds7U3ROo91CigQ51GDdM5yivT5BkZ/w/0KfR6z8/w4eZn7/a3GTz+Oxm+x1iVIeiwHRK
exLNTtILgmIXkQfXQNpxVxd108p9/1pdMzWjNcztDSnyQuyLV6EislYTfEeyH2qx1IpnNbY1WIXi
mEtCIim2s/Gz2td+gFXYzOto9EA27GYaTWLr5uYF+uWbST8Ufqi3UAU0RNS5Vxr/drX+iMjuISab
N4pZT7Am0gZkF7cmbTceFyAagq8a3Ug42FNIjQx7ABZpLL/yHjz4fBZRhlHr2hY9HPN+P/LZc/E5
cQgmo0wKIGokVGKRCo/2ci7+8Uc+axvWEhTI/FeZV2q4QbcbPZIBPhqQkleOoNqOi6T6DQgbPtD9
fguTUemiL37KP+t7HHrqQwv7uL2KJjD2GO0h4GXTxpQLNu+ccs4b9Ki9ukzT4hVfqQN5ggHZ8J7p
XiyBXbH4oXPH1jXI3zG+/QmZiZaMziTMl/rnUpk7G+5dtM290jl62LFubaSTNXf6UZ0ZO5JKeABR
N0U5Fjn8PtfPIRtoxR1tyynyMxLss3NRWeu91GW6efkwhx0rrHM6wUlps042hBljKpR0DK97L1Xa
Wv/ooZJfCZtkgJy0pk/mTFYLaGN36qMJd8w64DN+KGg8He1QCZ0zwAH+0yGmVa0s/1AeCK/qsEsE
rTVR3cEmWPaGLmWhJM9viZSwNEmi4xfWOGmNhA+Kgwf/gfM1nV6OviCnbjh75i4ohbx54ki8OmIO
1CtvtPVuh6Be48jwdTy1WKgKKk4KTTZzC2TKeuL38ukGJVWFzZWU48+ycFSBeOQs9UROT2wDiYCR
lVIPR0t63bUEQdU7LNMhh2xvBFBLJ4iCDhjHAdS2u5Q8jWbjK/m9crBRnIspA2mWggKLRZbCD1YS
LaRngZc63DCtYrRcaMbJ9iIjK4Xk2twQD6JOD/n8usLYZ0GdwS8+dR6ZvwEedY4ISN7WulyHPg1U
aPMrEbbvhGCzqD9ZAFHeEHZ2HYGJ9a6v1KFUQsRsc5Qd9ubihTl5mt4hZryfAPh+wum7eviCZhwE
PiRuscdkwSIjwLeSlGtgd9L/p1VQ42cBzVhZvLk2gnXw6E/6s8pBHv72zETkTGrRhbPRGTFmEuQf
opE7zwog4BIx4arS7P6RBT6DZxVfW5v+rB8XXpG8iBg47q4AneGRPZeWPg860sorewW7VcvK/y5N
UUN/YnhEbbb4KkvUNesCuAQvpZvbD2hIIb12TybKues3MCBx2IyUxKCW08XsHcLyC/MQpyxIarK9
nMOas+WMlRLuDjeqv45Nzd31h0R4o5TuS6jiXFc8lxnH/ncERGB1LDC3w1cmkY6B8gYBM+OwhmUZ
m/mwY053miLmcotEsSYC3Kh7xXZhZyIr2bhGT6EdjUfYPlNVxHah92928VwKOF6y2Sp4NoZrZSSz
U/O0HcuEd+6EGWZ+geCt2tF4nKA6eKyu+Xf4fsITrBEzIAK3R/xJkpgVqoY//4IYeLnaRNkl66zM
KAPydQXpmoa10equRZ8pcvj4GbbIBF44cLxGYTfeFprt6Kpkb+R4a6STcTMc8szwmXliLmqB1DBN
a5YZ/c/D1UBb15UM9MMLZa6VaQHS7Ik64OEwQAm4THKcfxXwHIgWa6bTerv0jjZq5YUbj2tmiAoT
eQZrqsjOKQl+gQ6F8e58oUIdF2YNgXawGDKltueMu2hloYT7ScRoBo5MDYwy1oLA4gY/K0g9Qn82
pNT+Bqaxj1IRe5oYi9eleFo34HtZ3ovizqeH5PoiSPG3HQsRbDLit3r3YvfVhYC8JXbuACke9857
5CgWrzpBOyYZ1wIgT1BMJjtWhT8M25cUcfpmx0rhb+qxUDdyr5I6dHqMc40mFAMDUbdQETOcswpj
bTgXPMWW+7mCDik7II5GIdd61wlSenfcljama28BGu5VS6lHHcKKDA9C6zfAneuMdzTakCh4ySa1
iR5d/EeI7RxADXbXHqwsDOjmL7rTt1Z1UySBIoc3h2F5+UjirLd1YTt42Z7mw7F/aMj9DX5BMS7y
Dy75FORAwxTDP2/BqTMmbPWmmJCWTH79xc+aL1O41DLylzoJjU2bLBrOuNscyGHlMN+kaUNOVwZL
zT8dmufaUJIRvFSaoKWZG4UMTiE5cj1h7Tnxsghip5Q2thepFqGowK6/PRQCi84W8LIm43USZOHD
FDR3np5P9FTIecfyd5YnSajGNp9TYku1UKbmByWen+uq4hcYnJnNQgfSF20ePjQX6X/QsLpfpAqN
F0mscpQybLZuuxHLFj1Xnl02l5sirI35PIz5dFaOgEqgV1A3cu0Nw0ZNp7vWpQ0Ai7/2lkNpweuL
PYLd1EwLqVrwW913dlkwEn+Bua19/CX0u92sBOmOjWNKQdg4usVkzlr6/G/qXVw5UhstVJ6FZ4dO
D8ZGl3qfd+UzJGMXUZSIgxNI8PtlwQVnbkkctuCHVrZocFJvpSA7nUqPS5nNREUN1nobPLUCn/YC
RJ5Hh5lZmGFME1T+YJl2sJdPpxWKKx6tkVLSAdi8FKqmDPXZlIH++KDlK7ps4j6iBhBiHhn8yZnR
bjxjP5Q9yCZeVBj418z3IpohdRh+4iUgze161+CZUCDTvDJLTMkfcma21ASg6Ockg6XdWEg7JRnC
TZnybCT54u5tSOisEnzO0SvNyJdu4TvtpufcY0+6/+96ZMF475ylH/kY+/ghumSXRd1fc/dXr2XZ
Bctojtgrp8M3IZcNcnyocNiuO6GcrR+QwBkm7rMlY2He3gHTKus/5XsbegiW2cubNM2Y0NQFSRag
UDTnI6tw9nNlG5W/RFVsAd5l4CEvMBi1X7LszX4YO0ha7HxMd71ESND7v6arkEvXHFKByoS8HduA
l0a2+CgnESo7gf4hoiZqWq3Qgrr0qgFhaxnMgJke+VbvqyVCfVjh8rXFpfqcrAw5HPrqPoXBcEiw
D7S5tfaV50i0QBMXBvLOU0ADR25BBVW4Co04ThD/5naNS7Mfdx9N2JT6vRHzhpsXDI0gCOpJCXjr
zmckQbKc5v2cQi/IWp7Ac+LvCpSZwXYkfYScvfNqNcuLb++PrlmlKMy92ki6BDq9lVTg2VaLBqPe
5rCB/PbWvTWkiHuM2qC/ze7xFG7TbxgfW4iTR1DxjM0qdT0IDhJPrdICjZh/9jMe/ooaA613+e9q
F5VR+HCJLAcqA4rbumDtI6SNEpCsFwZ83ggqwCeTdB39U1boaiIoW7EcSEAFR636DtmcCVbj/UuN
IbVAsEtZhw7CmZsOy/XE8kcnTxokuuUEJKmRyuqboqZyGIVt8YXsqWnafl5k5LWcu9Yk3hJiw7ja
4v5GisTtz9tg9be3PbFvGRcVFdTOqrB/ejmuC+bxv6LyCnzYbZZRc+vTr0o0CojAnQgO3VplcZZK
2ZPlb3Ly7cpLLdHTBrLZRBe75MWEmdpGntMh8Zo3IFJTdW5c1MFuQnceSQmtsxt1vlyWZV5Y3xpf
znnAnRZI0AV1s9bSykqNBVZbEPp1a8a3H1N62+vM1thVIpv0MZiOFCYRwD35wibS+8EVeAOVTIuH
mwfXlsHEAg0NJzqP/+STx55jE2aY5RYS3n6ifCyhMu8jrjMRTvMWnmZZcpyU2TTRfiYuBlpgmGbX
F8Om1L2x//nMgdQHFKhSGTDjYttjiXRF2lIduQsGA2zNjh9d4V9xf1rVMvEuAyT+4Ftr3uby1V0/
jCxruewmOKUWbZ150t+Mnv60t2ilRYiTODBf0VnCONVG+Xq9EBsr6v99UNIuJHKSAR0c+WNISR7V
9koGYYecRUPVkHv88ifCChAb5mC8F78VkBy7Rfxxuhv75UN4zxHKs/BKA3mHvqEMSclPY1YsW1jQ
6ftKidWafzkqj+/BQWy3dNapPeKmNB1TtuYY4QkcTUUjg6C1rM1f5hCyW2TysVswxlC1ivHlIY+K
+I7aslOmLNIAL19oHDB+QsKAlYXYRZau64MQqvmsbInTSkFH51U/Ss+GrVnfYQh3kx++anFzn165
cZSUc9vYxFJGXGgsepa+PbQVt6AfLDbGxgwfwYfskzO369t7casHC/AN2ZApIcCnIhP8+PS6ewl4
WvLifPS4IuTzViGVgLHl4kC/rEcnVJ4SKEzF3g6/bf8L3AmsCb2t1u0OxJDDDU4yFZZoewHg5hjm
Juf2jzG2GyxKx9iVMtC3pHIDTvv/XWUEZTGT5VA6gn7qMQjKWaWiyHMosaR2S5P6KWPirwEb8GaD
v0GHdBhrdFCTvNpOelo5CG4N68fDsycbONIcuv5EEOkjWX3VwAfhZha2aIh4xzMBAtQ42Jz4CdbE
Vr+PuaJbZst7JJNh3YT4xoKYChFNXlymjOS/W3e3qMONjmjme9/U9iZniDx9hlNvPy4gvwwhSgXo
fL0RlxgylQAz8YJO8fbIhAp9UOv2TDr+Nu6hEvoeZs53UG1ZPrZUbl58v0p5/P+4FlQ7T4iq5dV0
uKgPeyW0trSevOKZ0+/nxAisFFdIcmTXj73iA2FOTTudSv6FeY1lFwHUb8xdGDzs0Vv7fnPkKYlI
o+pv/5Dvjf+jouO6w80boJT8eHlUtTxBDpYC5HH7iAnPT429kvfP/eQir2Us9wdDb/8kZx186B88
Ndk1l96XC/jRlvw9uis1oaa+FN1pj+BUy3LmNaDDBz+mvoBuCBowqdKBWdPX6RGS5vAz89NvN3vg
XAVtinvZKkqL/nuctLRywmXSsKNAC5ILDPIoRk2DHm44QSRIZbxrcdNHCg+TVRqnhQj7moRrv+ls
4d2LlCWrrI41muDP8tuO2gt/x3kBUE399eEc7mLlomzklfjbsuosd5BTuNodjf4wYT0wiCBDMh41
gbbn5AiNXEpUZDYEp3NGLA9W8IvnYuFm4+CBY+i5zW6g3MdGVjvhyTNsZEC9NEnKbU+BwxSUiilN
bR/zNf3PTeNcZB40oZPt6ZB5p3F6KmFbZ1gd5UHpWuSgGdmOa3Qd/ZTUcOeh/fVnD6OssznglMee
DCMuALYrNox6BfZTPbqGMj3QWdp4Ht7a8o3zSeffVxY+17Oy3QdCDb9EolkT46vnW/8oz4Cjm/Gx
CUElRXoXfdOTdyQT1v2vbUVGhiIYc3P54CPyp1je8HUPg8cBV7gK8bU+kEoxV4OUJ3xx+pVMyHot
amh6QwTeB/xoeGiOEq91zqdmaA0R8waKjWc2Vi5IfCwVFf88VKBm9ITSS0GzEEap4CWBNvWwtCq6
1mB+xsR9u7fIRLEFUy8QCQsbMwjYEui+MePPxa76rx07be81ZDyaHzPZXE4vr2FXTDm/CW0hzifR
e0PRJpMcMR1CdVM4ImSYcHK8gDzhIxJjN2uhbLWRTj4oG505HB2pY7WjPbqd8AywbSkgjbNsxooM
07K/zYvtSdsmcloEO5rFDyhsnx7MRPb+iz6SioMfh+kQBH7jjjr7nUNy9Wq0c3tWKTOUN2faGMiM
MLNuz/1CGyB/oVUrGZu27Mgdq0/ETqn/hBUX0GrYYtpZ67DKytJLqn7bgI21SAugL34xqbnJgz2R
NR497KfOz8Yml33LEl0SB0rSvkUPpna0ko6vB0or/lV/ejz8XPj3PydyuydGRi+ALSqzfE6GRfWw
AI0wdT+GY1L6Pa4SniwUhxwdX41A+xkmhHCrCX84e6ctWDnpuxNb8CnIY3k7AQGaV6fr4Dk9pGwQ
fWHXK3V5whJx++wbBOsTGX1A96AFyetOkrlDEwWP6OsgbJyziyUrXTjnI8SzjPVdcyJ24ySstCTX
9xwZoau49QmAbheeSbopDwzbY/t5Bhza7N1/GfCIxhqOYRt695vJrIlz/zItz7LtJYlw97yfhcGR
AhQeX+bDG1jddZTHI0cELQr2VWfRll5f7t1kuTT4LtYhBriEtUrGYRVLyWgwCjsxvLXVFf+3CptF
eKFB+uYIJGyn+bZe9JbpX9rd875zEda4crY0VfN2nS9t4cNpb3RSwD330bB6QH7MbDWkWUmr6xec
RAD25Y/S0qd4Rhkj/MfyYdmCEXC+d0r/6jS40hkupa3xuSszQ9aFE3mF+P+DZ1BlatXM+bcM+w/r
E0JSIfsLxkdWuiPVACTdR5t1LuibTFjY6u/+2LbQ2Vkx/SP6+4pqfHpZSlY5tu/2x/yn+D0wCBRr
RkfJvyEN4kAIykNsfzeds57eCwDj+Y9YejwTyKJ19qbsYxW7FeslLGxoJUVVa6rdn3/Jhce1ER8s
StCZpJnkeYYZ1yQa33p7UEdFvEs9Cj18jq4A8/3NjWCtdNqiGzWy+7aPQzeaeF5wUdKUKyj+rGIw
fO6eVuM+qIbOo0Yk4rKI/9nFgF2J+ZPdhzls37y1FPXUWXw7fl+GO125NyIP+G1sK6xV6kzvwtGJ
8XlQ3P1sxAgplJ28hBpVNrg5xndtumISqlFa9748XgfN4K9QgRbPBEJn6lInxodz3XYV1qaB3YGu
AVGWxYG061YkAl+RUMCtn74XNLff4x4KYnEi5Bj/QuzupdtjfqvomGmdImirvcwGbw99psp9zFs/
AGB3zgVfSWIFsYWNQfVObOijqwrLBfqPQbVr+ztHC4VsisJ6bs6/i9VbRKDF0HZdOJHsY2UqKiDR
jK2nuir9cz6J4L13PqhjZlarzHpngSEuWo+NzoGmTrDcfAg4Vr+mIVRfhhnBDbxzp5e39g2IJccD
MZl1jLQn7HGfhreePtKcUg+bPEZBsUa1KO0bc7tQCDRGQyHs0R9pxoys02gsgfxDDgsEHomUkVMy
zIThm3gwJP1ZFhgYrovXVGRwOYK3o7/Y/WoANP5X9qVaLXuoBZV4Dwtsjcx2LjUXJaXreQd5Wm3Y
rR7EHV+JS+pwoliTl42uNIdTFCI/dPC32DgTnk7NYlJu8+AZAxctxWEVBTsW5exvRAgKEYn9Zy6C
CQx1nblQ+g3hZTgjbUpBA6SD6bUIUqBXHpxMPl4vNiGMSSxgzvqyu63EvCivqRTW0TPuR/kD0dkw
87r+d+ZMRyTeyvDk/HuTZL3K9nawq6jJfGr2Hip6Ipg1XB4Qi/Vc+cYm23uVFPHNvIvT8f7iL7Eh
PqIzVqY77kNK2eYcZfCTxvm45CBYWhhBKu+ytszSLeSgJVJUCbeB1psSRitXA5TL++y8vVF5nSOD
2X+Q66cX222Tx9pDn8RMM4KtukdiOdb3goaj7SGqqRxK0jtfXX/EAYDMehw5QBKPv0JwiXnvaZ7g
M0zUck2SMUfcTqwqifP2CbSAMBAL41kAljr27lGvrw5GGIKx59g8tb4FqfZdMas+xBMx7kIkh06q
6GN6QWz+hc3T2S1xg9bdzFCw/6JxV1ESyDM7nRiXFqnWaSZ+OKBfOU7Prh76UQF3Po0Iyvbow69f
SobbedPxWQOr7GWF6nNjtXkfdTPNQmtFsM1hID1jC9et2+LHlLsxNLHSoJxl8H81zZyjnGW6efjI
px4zRAdAEnm8ZhMxYHWMyooUNyiroF4ZrrONh9gYTwml3hmLIkA8QBEYappxBIGLcSUxppHKdUm1
xNAur9Mvzvfv1N0C2X0oZBp8CQC580y+MYKDHIvW0EGAMqHMz5kaasW9eWz071WOmR1xjFxxbtJK
vGFuquDk8HjGMyyf9x6pthVsK/ihy/O9DMeCfZZkxuf9mG0BOG3FyRmdcArk7SmMReqMG7vo7xNp
uvbPRTaNmvnPGdzt5JMbiFffou2fBT/Ngr/WB3QtCEuc0mWQahgJSeYSi8hWnWMyHHmQoIYZOqEJ
xsNyX+KEoBd57UIbqEDACvrztwxNgFCoQ5+1la8OGwX5RPu9JYETpXthUERClDJSCgLh/MaWJU0z
u+q1QWCoEcs5rVjS+EwbRrzOwMz/E5KTIqb5jK0jg7Ij+0joBIRYyPNDa0MvpmrTYCV284n3m8gY
+O6X7tcVBaYti+PgRmGXHamG4U/spcqlyWEaAMNKSiXUq5b+7hLax6T0BxonrFYYfnJVan68mfRW
pzYPnMxni2IUsurBa5efuf36B3NkHUpNTgd/Mv1L0Eo6GhpiFG92AZSnM2LEAobO830yMr5zhRj1
zU0X9NR+LL2h9nJ2AapkpedES+IeZHZ4RbE4lURghDJ0/EtxKUOJtC47k8nIjJ48f2jnmN+Swuly
gy55x2G4azYEBsA/MXmuw/EiklbZf0Ow4n2p+nibRYkkb61W4sxVUccUQcKpHBeO5TW5lUc7DWc2
y8ShDIbXv9kjZYEh4kJIrm769oWTGu+zbbYH66aCCna9/zd+NhMJ9y2tMRe99zHkrrdElVbOFbmK
axoOXB7B8HiyuaMr7DJzm84lFv1JI0tOiz+p0YAt6eZYDsQ7F05++yTmVhi4XsDeFHH62aB9n8S2
JHkms6AmXEhGsECAoTiXWZHhe3nV3cNbxx2kuW7LGzKRrJj9NfxqjWYKwB/hZ70c3p3XDzRENHPY
T0bvXMgI0/kMwl9F2u/NJEWXTzm60z1Obb9J7TNLOMLMi7uixipaMAHJdf8S8TiihY9jPz64shoU
GvbTCn+BZdq4yL6MkKxX5azIFHtoVEnF+mcCItalQTaNv4l+dJZABf5uhSb3HbTrCFtAjUDQzzwV
ksUri57VkcTLhyBCdtgAXLC4Tqm5NPrO4DB9rhsLGzxsyz3xFZlkFWpWFwqhmak72TZ8ogAssZv3
0yG4BXj7ImkO1wHI3/kITq3afgmh8DiNfcpq1M6l4R3q4pj3EvM/gNNYROv/iBgBT2RfdGh6Fdnu
M3Y6ZKee72awfKdZGZxKZPc2LgkZc/4yZU+fmiNfaVd2TIoRSX7xv7nBv8UfeG02Cy2sJQu9juA/
7up+z4eJfc1Ek8J+TBLg1nbZezOinrTOqiPg7jDYhF73Lx5JlFlRRBxMIXcwLbr4oJ+DeQr9Sm12
OuM3EIZhXKrpyNX3QnpoHmjlb9S7t3XVt4pDVri0s4hnXovu2IDrrbpw9paiYEyozqISNJWX29lU
aEMIM7As1rKFeE4nRAeGlXMZ7TVXZMF1rq8S0FdAOpCYJ2FZt+NiglQGx/owA/9bmpNYUO7JdPBj
CIRgNLgVwNY2gjSBdOd6US5tWJfAUpI/EouqzxF+JjgUzy4KYyF/MmXH11Wjh1301BgPEufT2oF3
gcaNkNUNEax8wqHwjOBx3ueYGOCGOZb14+ZXMl+Bq7eEwSvC6C8ElNqERF/C/m80vq9ePjLRsEiL
I7HHXL528kIqBsl7v1Vt2vQveCfuFfKcXr9OlOY/SUfLXwAgUJBuiB5q8FeYGQVIgZY0a2zEEx+l
UvXOySCFIw37q0WMgEtJwH13+PTZ0PBgByrz/hgDqn49NoLAzxplPlCjYVAHz3JddckLnfzfMrOA
N8ZmyTKWoJkSZxtftbDreyVSUlzleak4QBfPeaud7TLbOvHfPXnEPuQrFu6n8d6OK+c9tbSVBwRI
4nDIfWHNMGKNm2l05TgGOhDAKqhEkXq8MEEKkYLXN2cgWwbH6KErUTcVoH4EMMdYZQboJE+5LCXQ
8/g7HxMpUnrgGXNcWjlV9A3BP56An8TBn5znBgGKDnAQ5lCUrfZhQDO1PPPPbHXcR7nAgcyO3i++
XiFUQbPCJO6jpjPJERBmiGbbvrCgOEOfA/mkCxH0Pwq90g8oUMFbTs677o813p6EeSlMKmccDk8H
+L25BY1VM0d4bbhBGECJONERNTvEi7l8ZkfZnddU2g5Phz28l0rsXQntgX+ftpzEobskzH/lRl4a
6v9Qwqzx8bnY7QOT3BUwUGTn9Guu7pVUh/xAyRO0NnlvyOqr78r6rz7jU9Kw6v+95rxHz/4UlkqC
OhHoETvFf8B2/YI6FDdMTNui4FHv8rqi8P4wybPVWh8rBl+szIh9WuL4sFb2qfOxbTT4tc49H9XK
j5Ar1NAgbMZmv2AeQzaF299rcITf1BipBflWvva9eq6G+GDcHEyHyX7G5ipg8G8QEOhd6CeIkvJi
6JtP1RpLg7j8aU59kcMHDeLCyJc0TCJxAeUT5zkCcNb4OgaLCsEjBSFvYBNAGaay9UXoLjvKdWDs
IzC4XU/KCoLRaHgqUUBaQ89BL0s/iu7FZcAt9uxdBSOtWsRKPmmgK+Y2tMoPGqTAv+hmQXZ/ZQnu
dHawTg9yqRad0YQUGsfpVwG3tJWdiHwXX/ZA8biG3f3cRBGFL+G+ZG9PZFH3dEX9H5F4a1THw1LO
d2Jtf6I0dbXlJKY5ESgOIiNnHk/YkCCwKRnIP+4q5hfXMwX/vX0STdjFvth8ao+h9X/ngv926v0L
bWWDhrpHlaeCuESH5VWFK+Azfcled3Hx+hYjm5RPPAuRixsB74EiMyam0ZTd5XDix+9M9z+uwcox
Goccs9T3V+Tjs67XergyGRxbAHKwp+JEtmul0IiIgXp/88SfAwLJ8CMj4xjumrfCOHMM8VvPpeu3
lxKgFdSzKns51YEE/ZYh2X+i7qWLYi2k8FQdf8N5w8Kyt/8k4mGdkXJeZBtAAM7XlMV3pxj8bgxL
QCgUWAdL1falRl6fla9aLGWiCUD4WgvotKEkWliNdnbhuHQmUW0t0Z0PxQBuAksle/keGjC/teNm
RqSY/wVFFZt/EdMs05bJJ0MGZjXHfIfBD3jVIkiLlC10tM6vQ8u+kbal9xBACO5hwXh4Bd9EtZ33
ylavmqQw0RnbizQ8B9hxniROYVHsjbspvgQaDXUh9QzQxJxhSFhMybU0U+I6jZ/I/LUhnhvzFbDC
9zeJ3bflxcC6C2ywOkFlWrVni2Odwguo23GUdkN9BInLzcYxa2tIY+Fa8SwSumeD7UkzrJsdrFfd
1HmEj4dyLQSf51HkK1CxhfH61mPnJWtBTgMnqH/+qX9oLEVXN1ZCLxMTYWWRbTZrldU7SEJkGBqb
c9iAynSGjPdMMoMLgiFa1mPjYOhrT4qB0UEr5q3Tu4Nek0d9ur+vs7u11kw3GSxl9YdHEfY0uDfw
X7655trYhxZXc1mEork4b55AaIW/TmYUVhkC5sVCpSy3kUTWddHs2uYeEx2f5Y1jlMqLDJbDiDJ3
PrwAXkVT+SF8qqDrGb4yR/JYp6c6oZvOkG+/NK7ZGnF0nxKS1TLCdDYs0y0YZOjd4BMSGUWQdQWz
0SYEmWLPZyBoSRWU5+jSTlMiMy5guK47xkYJVdOr9seOcKrfM8I1284S1mOm3TR5qINNQk8wlTON
a79+2RQRAfP8v+yZRYMkUtwcVUsgtV3GOEBN8B6SeUDfWUy7EWjWlZ1msZ7Mxs0qfO7saq68Kkn6
xkXMORl0ibPRRZQ/KP5SGvxH2FFVkai6x5QTru6oPvrng3sm53cz7N95bhNJZHbm36C6M5J2j79G
KszXGjKQ5FrilleI6oAIjNERQmS8qBAJv4zA/ngn01KWt2f+WL0oKanOVVDhDpAgl3K/fttHV7kM
QHEHvk8R1xibQD1B0fvRPZ/TTo8qiv63+qp+5orQLk32/ZKZ0fSWGxKrS7ZKMb1ArPrq9X8Z4FZt
RSQ+FqmyLZf2eggwPgATP6jNsnIgJB+ELDcRf83CwlfOxaY6fX47yw54QiDDOWAcpXaRO6fioTu5
6Z2+vlgKeEW9pXFzuISOQbpFcbOSvgGeR0VQLFXVxxAhGzjAbWEsDFNWGgdfP48n5rOS18KjMncI
8WP6MCH6ReGHiaxgBdAViA6gOSMSheH0iWIeqpNmkCq243ahCAhvUJJvt8B7SlKOWip250uh+Art
FDuTmrxJWEKNQBYUXw+YnXpJCYwrAcpjjsfSCHd+bQu7zMbicWW8rl+oNvyOZqZoYhKzM8Eb/CDJ
ZReiylQcmLh1mE3FoAD1HAQteRRfc3j9OL5qp9o3L4hUtNs0eQVs7OQFtDM8/vy+Pw0UZHieHEec
WaVhWAcNCWFdo4hyI4QJ1Jz8lS8xq+KjXZkAnnxdOP6MQ9jfcFGi58LETo9Pl2XFNTJpuQ7E5cDh
M/yTDcZkK6mgzFmLRzwxxOWl3ZO1iGFpT5CktVgVtFq3QpDIWKy2N8h99swBvcpTZLYxdscBeDJr
oi1ZPO89T8TEQ+WePKK3jnrODbfgPE7FMbhJkrf3YxB0s1kIC/qtkUJFsYkgy8rKdxk4MtmK8njx
+EKkp68R9rrq9NvFF0pdMl2CCPFmxS3Bg/ylibBC/m35k0tQfVSXW0kri5OQD76387c0ZZmfMhmy
B2ef/8C7i36lF4vDf/agSDpBud9SqDaWQWmzfbCRkP17QhGVkPa6xR3cuAT2pK5/maw/sX1zJiWV
orOVePzpgCGJpknFByqb12F6Mz1A7sSZpIcb1yDlJAY3m6beBlp1cL1uS8cXZuXMPo6K5Gqfws23
KcLvKUcufTjxqlVFkzdwIn/lmCh+9WeV/GhVyEtF/fj6nCguHe7aTgtUPuuXv4OeyoKC5Ow7Foag
XXaY2fXVPDqXT21jLfjambQEWkbClo04ygJl4fq1pH1QobwNdD+ncZht6FwHolasDs5dcZvcYXoN
exhJdUFOZDoQovM8s+QkTpFOz1vtT/+djaiWrIJg4RJ+DbDmO+KkSIKWJYsCap3XL4E0pjPNCU6P
y7ey906BfAtOTGAqr0Hrq/GvdTSEXEi3L5B4T+jQtB4ga244YfQWDbNXtJL9LmDhKiLV0gxfd/T0
Lg/OLjC/PX9j7jsY42mTjyPkIopmSVfIvxjYHRnTrUhwQogbzkHrzZYvm9ykNShfnUAYx2/rsNyT
NYOCcdTbGmKRY3fqrvV0Chx9YDDGdFF3K/SznR52OjVySBFThDV/fvKarvLZDs/G2mI6FyQzEI2z
BI4Y0kMfNELEzO3WlYWhY8z4/d5AQ7uBU1mCqTckK1x2Q+S5Xtzf6IDvDADM6RuEqkIXrxDLBK8Y
bnt70ndOElCn4dTkU2QsMw8Z/bujNxmbgFagIt4Mq7f4gn0b8apTOzfvbmTzBnCAekycEUz6jC4E
FndeYfPjyUQ1gzaIMpsks9WPL7cgJS0rdsCQVkL+JoBWRxMqdgcesRqiZedATE39+Sbr92YYbXp6
WkxCNgekaoaKHDwTlcsXevXAbSww6c3CDLZLB4TNF7wNLBGoWdhUlXKwqdsgpRVMgvt26u+MF66U
ieeicRMTbXhEPqHVcldxDUvWpjFDql4DMF6f6HBRpk20wgcDgZCg7sVibJwk/oAOrUvAtgx42UC9
0lXtxgIMkQAw2mIjoD4T7B+F7iQX6YIygfc9BlAyFz18XwuQOEbuB1QAvgpZ0RxJW8D7TQGJ65r4
MTHRBI9VhSAuhHtm3PfWwOC6ToW9oslS7u7TV4JlJqrI0bOTpW6WQylObTUky4E7Sm3RTXLhBtSo
uGE9W++l/Rrwgf/XGqBVkAQkWoYXP0QQkCFhJEmm8vfHJT6cC/MB+zWJeq+EfsJebDHC0C4oPT7u
DmHD3HWbByHdGqyYxvDGHfrdWoUBasJ9Kgrdg1bjDiYDmrnJqEecoIlUZBz7ZZWxVeGLC4xjrUsL
9gaANuighgozUBKbXBX2LSds9xWnjVUsiS8U5JsFCeZ8N9ibINoNtj9En8abskN0xCVWNHSF7ff1
pB6upQ40I3JYuPWTXHEqtIHiDbjKafnbR6q+3WJbFmzcHu++cHw4mgfQd3METfbSgZPJ56WgQhhD
8nGDE3Sa4k/Rn0ZKJmjENgGTOVEJvwbbBSlND8rjxVeW63DrL94u9aX9tOM8xRnqmaGx4S3+sQYg
+luQOUlIelFM8pVXSmvsTWisDNO+90B0gpAXNy3vZPIggXatQXC5Xmdjvm3tfIvo2Ovq+lWqAq16
7fWgr7MHsZXTbfHGdpvnPsbbnoP+j6FYQkHn0pqeJM/m6X1ht0OtoLtDaRzCT5vLX+vIsF7UXTeX
m2hD3WtNJB2NAFfE0jJK3c2+1hh08Dju/3JAx44IhCbwM3M41swr7emNU8/XOv/hZPkD/sXNhyhn
ulGENfp9Rl9Hc1ppZYP4KsMR/7Snv66IeWTNaa5D9XIp2VXwF9n0jIBeKGo/kMeJivoa+QswDn8N
5+C+OEl1iWOgPY7UfvBBmdwqgaVPix8GhHte9Vt0VaC/b7vc9/T5KTi6g6oXSbJ8jZ6IyO2KO3qE
jYAVgtOnTN9YN32RAp3UdMNIIGQT1Cvosn+X+6V0g4OyS14LFqdPvSZpSeGyScVb1cvXsLlSTMbV
nhSL1DZifdSa59iuwybYeivjVQMBKR82CowZBvBDi/UR07yNX2/J38pRZqZekHqEI3BeS4/Kpuy/
5XdX8g2HAKQTSOFG17UavQm5pKPyNIi/FzuWww1459k6qkNNZ1jIkxJZgGcm6wGJzET9ZZTA0Xf7
h0XyUvXyn/758Uv9OYgDcwPTwLqdSiNWf8jJv8fGfAqtfeZ79ucZAuULrM0QmfgDSuhPTCNTqYDF
ULf883eTqaBPE8yrLoIQgXE8dP4Gy5U4gmzmhRPGvb8AmEUkXXsfLVeovLksx23g28tcuwYwQUge
JNLSH3+Uu1jXkbFifNJzw1bkjsHQ1Y4iW+JekjK01LF+0wXpQ/RTE6xNIQNv1PB5Krd1ABfMGC7f
3X1t++fZDjZqH7K31LFRcuinm/0885Hbc6TgpI8iJAXeUtITSTPY7GECSrbe5NjOX5Idb3WqTjGM
Q/TwYhLe8YxdUzUtDmr9tJ3iuAxleXNTIkUY3WhRWBv3p1C7cpG/Q0loc5fQAhAUsEPs1/g9qIji
H15UcSlANCfHpEO+BrDdC0BnzHmABs8S1IVTB6CKzU2ZmoJ1JS34QBZxNmYCsXDqdtv/xn4f9rHh
ZfL2w980WOzuWN4KHufov2dL+P8J6LjAdSy43ASyiOKSvW/gUoFZqxS0bk4PkciCfMxnoQ1XOfbV
43+a1jqBRSvJlNMFsGG6dZoZwt6qlMDpeUXC6VVj8UMyMyhtusXCixTsInjAcOem8cC2Doqvhft9
PokeLKyD8mcO4N92FllbM2YkwUzywHSYQCNlVgXnQziubZSjRh4LRXcd1cJVw2SWsFsLVT0IQv55
FWfZ/Aj9T0Lh6jSTr5tzjT8fRaKlb6VyV9/wsdrhS1DTbRc3SqX742cZt1QoMwbeRU4ePh6lHdOO
tmvLJzp9iRjpyxvMhM8unpaseoDeVSIDRZf7W/uomrL2EFHgovTwySL0bWMspQsDKIM32hMJYIjJ
328DCI7LVlySSFdJuvNeMn8ytfDIySaglevCXp5zlZdTnq0v2B12jdLlOxGj4FBX705FJX7RHnnC
wgt/lKg8eEWV063EQW5TBLibRf/Wv/7CZDe/A8kA4H5mAXx/kPLSk6XO+IDkSz1D4FUCj36TEXVJ
Xl/OO3ngnjXoID6Cf82W1spu72PLRz/EVwzeh0Q+l8eTmqzK5EQl2mxwDTBxCraXb6PvTX5gd21m
wlsPbNB+YR0ZKPmtNv5GnGZejlVxSVWsD/mZGBtepSblLSlIoR/fB4OQPQ7eoSswC17eYJ1YlJb8
ATyxBO94M7yLo7P789xl/MZcOQeUesao9COe7vVjnCiORMnIVQsM8Fp/+MEQ4wqqG55BG1alX6Pt
mdom4V47MUBO6DszWbm8M8e9LJzGR1brOIrufrNLGPz1BoXK8wJnmQlQ1d6iRQ93EoPyJn+n7s4x
XaiBJ1GRqbjXwjIdmhOQPRrwjyT4yiNH3+a8VnIWDSXyX7mGPaDiRjKxFkiyfugt+nVkWngpjRgS
AgoNKUdxBbopmkay0SGAuvwCfcp7rE/VPkEnElsb3P+g751WmziGr7m1HUgQ+VTX+Qhjie/Y74bq
3iUJ5+6C3Rf028A477Z9ei3skvT66z0cA9hl8OjgMZoHTJBd1Z5a4QtrxCPrriBVHrGEsPQyf0dh
BXckRaplcvzaMc0zDkjuwxj7pa8/JmaToiMvp3G0/4wCWZTD2U0+nilmIlZgj7YcC3CnChFrIVQU
AZxVv7zQgcMQWScEtdHKHSb0es+e9Ee8byTQVCGRnQtMxNVFBG+BA9PwiwLTX8ZDHee3aA3vLHVS
3PwSVD3eNdTsohtEXyrSB6W1io+OpBWGfeSK6IPFyUnltzT8euQHY6GHbYk/J1Sok0opIHZsgzS9
6//i0fHYvrm/3wPwar9BaST4MaRz0irsBF5mBT9YdFAJWF/TB77migY+otp2G5xC2NwNmdQfEc6u
KuCiHDFL3RiwclbNeksSR1qDPrcdiI+zoDKFyBK0W95EeJQLA9Z+xq33QtIRQqUhvIqh5J+0wbOH
s8xcyBuVVokCUDjk+ds4sUzx6OekxqZsD+BRhqAONzmZsJkZd705Rm3SOiml8YCAxQShDIE6sgcN
n0URGJctCwz+z9UNsgHtU7ih0c//iVbM7WeUn91R4HSs1jsmwiigr1OdHnimMj76qxyYkKRi1wq4
FcO6B9VulJUhoYu/1j8jy31kMWsgMjrJ5wg5hVMkaaAoGCTvlqkOl2fon74Fqd/0WrF4G5+xBUcz
rGs88T3YipE+lbOMh4Y0spbEwHVaQZyFz0eMh1Chm3k8SRWmJGy8qRkqMqNPpjnq0BSSYFXeEwn/
Ih6Tu4ItifD4S9E8pagZpJ4yTQuvCUJzq5mDcREVgLBUtRETCKZX0up7I1rnXc/4Jk1JJWTXDoga
MW2+64ha5SBuWttaaf0uYqjRW48CKaNx/yiwi5yYdCuhWliHQGR8zoRDIXqUu+Mg1mQ/ShLHcTwx
0amRsU5oLMGIGM6wYqUVQGsoZxlskusnKCWRQEHloK+E0fnYbEV95+B443dAOPvAIcJyVKCQrsIr
t/2ZDlCuYPxCVP92R09vxnMQrjg0c3DIs5ZBEs5AvBD0wuB87z1Xym6XvQU9Oa2cWiqTsxT93M83
MW5cnVd8GW5qFXzkdW47diVZs7X5C97sYlZLKh0e8mZyHS0Vg3kmUuDALw6ShmuIuvIrI3yK3dVy
pcMSR8FdFKx4Zc8k7ISf0DH2xJWnH3aO28+kRn2D/oEAvy/STVPYAYOf6YcbQG8PML+VnsKhIbDV
2EjTyKig6P9udzZ0M9RYQ/tvC4Ojgsq2/TNj/1GR2RHo4Bpe7NbuUP6e1WNQhJTJ+CjonLRq4QOQ
C43wKsOsheyi4aU3XQdvZbkj0trrzqQLfe2J9UMxf0iGm3VsW7sgKouEUx/+MSlkjLG3KVpYq/sf
7u/sfnn9GVrTFLkOPy9p2BEPALQlp4M0laIHDbfgHKxCH6st/lOHN+sMLQ2yogCPR7MOqH0BUUcp
ET5xSdALe32i64FGfX8lMogZWRTnd8oGJ1Lr85zxG69A1UhEML7tipodEvG9BUFc0KRP1b7gk964
4aI6z/mdV0f3YafAsPeDZ42WzhpmKuQN0Q8B7ZUHpR+MJcA9CMs0sxzXhFv3hPcgSB1aZH+nMJnp
kNPE6ZV43eDmjG91M4kFs5OpUSLfYETi34DWjmbjoBLozm9thaEku65hVZ4HS30zH4f4iLI59Yjf
TFOih0pEKqG4fsspIZZKbD2Rbyh5nsmAxutSTq6ARmtGMmDFXA+863PkosRvtrMjlE2EaB/jlFdz
21RA+nixTvFwjcxrXdJcuil3n0hDz0a93/Ctt+euRPclszeELZsfO1KDBQSCH20rK5zkmjCnB9J5
esP0rDBMyqm6mm/we3E4h3NFns4vQfQfeKVO+dX5ERhsl/LGGcTRBJZtCnqk2RTpJU0oPfLMp9p4
6EHqC+4y4K+3NrHUtQdiysidL4eaKRJBWYpDldq+z9b6/B+mDKzm8890vpXCQZlt9iCLsbD8ja2C
H4dAolAEn9ZHxRz1twthth3syNZTBgZyFAE5KASjXJ+5NoBxBljHzb18N41kLQstIqKh0AMri7dO
yeCi9l3GVjd7gUs6+4VCGc8spB0v36N98kc9gpD+hz9Vg6gXefZAhWGSa5BgeApy64grgwn3xNE7
w4rAiFkvg4W0CJ5796sOk/VR539ISXxFVNeft/Dji3Ubt5T3emrk9BFL7OBbkuAYId9g1JARuBra
f4Ew97cBx2Tmz+r1My/2fEgF42NiyWUsVXLtMbo2L++Kb/9KyAbD3V5Axf8TiLqDCfpSeMiy375c
ytS1ruHV8pbEzhn/SOdMPcYSJENFCn6XYraBufL9JVwCvU64vFtCfi8+5vUIwcttwS6nLZfxzd1o
FPOxlXos2KmzgizHTizDyTOXQNEGL/QNxL2VPQ3+oZoaxYzIuIfMTCQ7jBjh2eU92ZZ3ebVE7nCM
Pduaae5iDxmHW0pjaul8imqKtKGVP9f/aHcOKOaQ/gaeSmLXU4p/5d50cM8N3nKItaVXtJy3tcwc
eGFC4JKZfADO5A41zmrzSk4REuff9l4kwYXuPFUFYuNYMAf/uJRbt04/mcMdofqEJusNT6+H/yY9
8ihr54KtmY8xYOPXUlM7KZoAIxrVtnRW1RbGx/24fsapTs9zJPBh4K+Brr2A0lVY+VD3iF53PMsF
4k//Iaq3DQHoPLZyaaKeykBOXwZn1eB0FLcWSiC8n2ksCR5A3XB31FN7BwOFqS9NSHrC5y3JfAHW
GkV1nuAGD10gPRDI0UDrXoVUMc7fiOdeC/eA7phwSb4AduQgB9rhmZplJSkmzlBsgbcWX1Xp2GFi
j8GUGQ0p1yRt+3JgGw/ZOXmC5+DHusqaoXGM+ON49O9zTLyi/O/sCtzIoNL/TTwSC1vTQkionE3H
xdc11gHaezSK4QwW0kVuEF9sEKdcjAiZPvSChOdN+gq6936XxtYSxgs1EqYSZ/qQdC2X9efwdVP1
RGG5cllXOEf0Adx8IhiLWj35L95WktHp8CU/UW2CCic6Jroup76sSzeRi9ATdEPGrarCFHX2401Y
QFHa0z7/lbYwcL+MOjYmPCyZthnVfd5iKk1eBMtg2NmDn5H/eZI/AkexzHJIBhluil3iRizXMIG/
qHX58bp/ijtxa1sXLXD9jS9CsprbUr23lbSmgfn3+xqusFxegjvAPaGCnwkb/5J+FoAkmTjjoxrS
TyORQ2rGXae/LfrTTPwu5lkbkyNc8wMAAlsAaEffW5YVTDNh0LGhKHiJvnwmMHM5JoYOt5wTjgyG
nT/o3f9xMhuND0ncefIEmpHXP7/rnNgPsfB6xM2oOrgsEX0MNj0KqmKuwY1ePmrjWe+OUiug+TZF
vlPj9PXgtyveIQ5NKn1dI6FUtbOBRYL0upH0If9elSIH6O2SGGdWbt9oMJV58Y0pdZVNL8/rsDQG
aYNlEOsUhNQKuO99onlP4nGEbvS45mkJhfXJJJ4oRVKsmJqdeiga9mUObCrY9XMks/yU6WB4SQuM
Zt4vAEmMOduW/Zs+BearsEkyfiI5g3hRbeY1CTzsE248NLnK07j4o/+0RBApTMuOvDQuz4RJSy/n
HCf4tTKhhA+gjXa547irxgcBE8DyDyNs1j56JPY0tQncv0ZhyNuYGTHT1z4cyk+9AE+uQ5/IpwEs
AjU0K7CdoL+LFpl0QTWojbboEZAvwGZb9i2jPZsOG/8I0fWcaSRlg5Hi5UdLd1aCvVMx4XYltRXt
iAB/tfEDGlxFCqZEs6E3P3MAW0XNjzIjuRhw2k/J/tetOrQNQ1JSveajfdaX9VjnGDXxadqoyPpj
GeAg/XoEKM56OmImGax5L8hINSzM7eRfNxHFpMpdDvNzqU+tmd5jrDbYAKHtPi1tAVc+ir1IP1Yv
r5285DZjEELIEsUtwoSI/Sf1ppCxKdKxSBTbXiNSlUQxgKHTDnmNXlEj6NEOsgnNv6q0E6hJP/UO
9LoUBy5YcXI3SFssc3rb7UXOvZ/CiCmbWcfkF0qAHEC/HUu633pX9wpoyIyMtJb4BiOVAjUbYnxM
f3P2KK58HMZKj9Ou2BTELNFk4pXA6XsnjptlhssXqKX4JU8ZDbjY4tiLB0fwwspsnoY8CacTibRR
8LGB+8MvOa2rRnWmZSqkAts8da9V5e3xXLQ2+JK6VW9cvzGdCFIeg4Gw9KOixH/wHKYnXiDH56z/
j0V4t/5p6lD3vBcbepHQikPgTSNuC/XZEFxCr2x32XOWICUSoejJCuZsab7WKDsi9y/ykxSd8lvK
bX/5auXNaF8pGe/BNeufjcmHG3Ivj+2KRAelvgfPheXn7p3VJ3r+OYxFDUd5QNdiqYbVG6mYbcY+
yArY3Ox/eQ5F4boE03vK+kEN925Ao66DxveyoFXoKVqPCEonlpRrXZj6EGcAivxJ7vh5uWtqcXpd
cuSKQcNxAS7cwHeq7hn8MZZ9rwnQpAyUn9MGZbh8F+Q6rGuuzpCuma5uNjujHff9MFPFlCYizZR6
D/B87/N+3iJ06V1UmxJRA04g0xisVuBYpYNLObQvkFhAzk8MtLlun2bWDt/tidqGSlpnR+0ndwrt
LdMwz/kweSOhpgg06sPT9hwsaPSZsU869SVJU1oDGG8+LjPcoQkb6jPNXMNfJDOobFkG9QJSW8yK
M43aMYQ06dZhvgv1H36j00Ni4Ee3tQjgwEAaCXHClw4P2zwP+JC4U2Z9cAHH6vjykih03GbJiUr6
4OPptMOhKUNsoIMiYZp/Wz/bCGRIUDjbMy/NifqJadsjvCOk4H1jLr/zcwhTGDvbsae42eQROmJ+
pw0i4pDWxONSc+yA0/VZrDpMGt1qk1ChWprHKBIz5gGzK8jaxxGwtUd80R+GqjlRVJCdZ1e+swxo
NSgMvBIlgVQsWSOPW52O+eWvl8isQKzyYEtFiqXypxtJtapgyMujlt62tdyAorWR+09ZOsyxcpnG
M6ot/bc0JCthpVTjn+zDn76PHZqf+M8Lg9YhGe4xbeKGjkhTTJ9Xt1Q0VDFrjOnzJEHd2q9XJsKu
yYtZUitrU2GV7TQSfqUa8AdBU+orxpdHXEBqeyw1Ooq3SUoabmfBGCQy2b6y6gCPc0sOwiQmVAwL
YIaaYfRFU1HtXASjpyMji/KswIUVAIDKAi9QwC7EveGnrt+q+E2LAfi/KrTN2dcIz4c7nysYTrW6
OyUMhHHT/L3i5y9AkrJoep5ouODoUHWDIiVKsWo04cI/CuLAmMi6g2D8mUs3mlIkK51w9qUqJzfY
NAhIWG95JqA+i+QgmaEscY1kc1opDQHiEn7JB40C5QWz6haO+XL9xGlXbZiESmDmgsJaXTs75Or3
GtUUb2HQAMMfwLNC9M8ElCzEJGxaL4jaSvj7VK/cM3IAgMSg+Sr/OkInNGOsbrpUcG6J0B+JsHG9
ksDoVpYUYIpU7xblZY30QxwuKx9w9vdaP7TUOhxAhF39vt2no6uYxYjQ8jVsmn7ijrynQUGavjjk
rRtdT/5FGy6lVg6QZI62OKH2dG+/FYeOtQJ0kQohj4PpOUM1rgzb6p2dbq2WVelcfDq3LiC9LJZK
LNWGTlsBsxdoqDKZkCfYXAnDulsuUBciIz33+W9RfK8s2X+BFKYR51IqLXj3nd0hTzm9VCDZfLrF
hPI8MuOEQNbUzVkZ/e9bxd6Zf9KQ+zHuYq7XE0NhgZyFrwWpz1do1wybSufmgSX13ywHpvvADAbN
riLRCb+Ow3jfaoX3l3IFA+SNT/XZ2U9yy/C00M71r0vBplZdKM5GU0RHGFv/eKb/KgKkNsRbfmtl
Ak5v1SA83w51sF3bpSyfmGT2816dVlvnfmoCYaM17kjJn9O9rHUBQZv24WLAqj+s62xDkvJKdMS4
L9yo7jnaFNi0JG6n9VbTiN3MEHoMbOFURqEvro/FNhFh3y0nKpCC81lOfOoqSyGeOF9k5ZymPh8z
JrdG211hUr5qH4srqPvluQC/f21b3So/I6N2d0qe6bj7vNQDZW7A98uUL50w8Ypzl6dlT3S451Dm
SY5rzT0rGsp/XI3TzOUlx2SuP8NyF0kUu0ylQlBJkwKvpa9oApYb2qwbse3XREzFjhtwSERPtMb2
eF4JmnmM1FnUhItacjZyoFbW2gru64ywburQStniKSYGdh8U+t8hwh/3NvbylNGKHd961jF3fmhO
scT9zJNhzYgs8wsxAuzXXjLxFrWIAOyHDGdiSPS4HnuMXcEZkmKN3V/j4Xedxt3rcXRpJfsDZfd6
2dh5hQpOlvViG0F9tUb7xBQuxWLZq9m0Sytcu7l1czYd/CRX9BenZw7tWvL3ldQSEOTuR81RlZFz
WDhpP7Z2W/GTvZenVgitjldt3fmV86QlzmDPWc8jNU0pZQ1Y6P3Hok08+e2BAczX0na+bxIN38EI
jD8yVxyZNUIDpdz2ZT/BiCxHCZF4Orym/Apaaq3H2PoEl3v/18pVCrn5SSEtrrDTAaLVuE20nMjg
QTwOkLLUWCIezvoqIMKuwACR2PUQR3JI5mlDk7tcOOeUo30zzM905+FtH6vi3LeFcCK2E+VlGKqF
FjkybBjabBO1q2QZyDu5x8Qd43HOrC3Cpa5mv5omMLwa2Z2LpO/loQxvcN+rysPxbMhMjclnEb5V
M3EVWD1eaR/gP43ATrztRCPb3/L/JgFmGji4/bD2uLNKy/kuLFmoSnI/HVy+Kf9S1V07+JWaJ2Hj
UsL4tkEDkMa5CY9/XElaMQ3UngJ64PO6T1oN6b23VaHMX/qHUwO4lh2n0tnEaTjYH/izKizBB64r
ump9sOqEP6bjOGxea31qOMDmu1XLDXYJgKrH/oKB2xsm7nxnQytcurZyUSPUg31zekGavtGdCQ0X
Iex7n15YLmfsiJXwVTIjDsLffCv4VWwTdL/lKoIPjgX/PE2sUzhBJcnLyRULK1SR+AZmPqF++miC
jueMIU2YMqDrcBYW5Efu8Qut5ogvPeJ+g+G3gV3F8toy+lgFzlUfONWy8qrlTmY5LGDA3QvAwRa3
IbmF7SidzGaEZ38wSfVCyMNvx1ItyKW6iVFXXEeTN0w5P6ht4bZrZRGthi8t+HHjdpyeyRyipj8B
ydGJfkej07oEHNJzgrtwHX0AlseiaiIw//Ek1ZhkAN/hY7dYMUsSngr0SgVWYDA6X6D+OkmK01K5
FJwW0oIPtISYsUd/7znAeRYx14j7P+5lQOgHnEr9+5Lqf8yEjxynj/qcz+gXL/smbkC+SCIlOcot
n40S/A/aLC5UwFxubsbrA3ohgxm7Fem62r3vFcunKvhcC162qQU8cW4aasDXNw2kq+EBCxx0PXYl
zS9ZzL2pmG9E5I9yBeyGnOjVdqIQP9coWMPB8m4INrFkwkzxM5zvYSNJtalor+lvveZ58T2670LE
g76Ar5s161vEaU3vt9tzl92gRfW5DjCQuV1GaR3YjbYfoIi4K+/s4FjswfDvG+/Tvat4qxKUKKy6
+cSn0OsawLNXjFEEi8mgVKjVzkw9fdnkPTr9mRRn/djwX/WXzQINMPUUNoOK92QbLYaLK+zf85pQ
PeCQ9VxnzsdOmL1waSNMk0bv3yWpBnPBvpZhcVO6DI/NcDqNLCSSO49LD2LGwbEhZMylyNnEgO+F
pVr2W1iaCrwTIOgilAlCekBxxkvH/g5s09taLvx4U/EW0WFMa9THILiulf0+JX5yL5DsN2dLWS48
ERCLqqY2Dh3GHzLijaNy6I93SAoL46oXeied3pFcnyJgMcMZVX/SkS9//bzYswi6UL7MI03cLz8z
H3WjsWn2SHFi8Z4O6KN88LBEE8AKH4lPt3axGL0uUS4Bwpt6FfslCDj8uttPkzeBSpicVRnO7ALX
5N0h+rVThpI9imEjI0atnFxlIAvrb3g48+FE0kYrlkA/10NIWNpdH+K/mUin3AXPzmBpXx9CE358
D4F9+np9C4TGRCQWr0KbdBHgYX3KKZAq6R4NUXrc6qWN5wc6xyXV0Ba0fgtvrx4gXk7yljv61iCk
H/UNzGdhIF5MVFRKX5CsVg5liWeiY3etUtdLX+K4qp5nit8hTZCbxW82ZHXFJlTlkeUsTtRsdTsi
0KEVa7PoJjqZkD6XrcR5udyAVvZE5i9xziU6/gZ2xTyrnqKj9ulshYLfQJGoHSzONd89dEAN6SDy
yqwNJIFQh4MBc+g7Iu1EATMRe8PxPCgyrrUFitSmgd1eoVKkyVevpWaGHV98Le7NbJ+C5zsIMXEL
nrfA+wkCWgq5KJbvuPzu0uDK5eTXd5Vz7Nkb5EP54rW7ZOyz4zThCbt2tWzQI/RIYJHClz7Qd68X
Ro8Et6lPqIQ9EgTwF5YzUHYuhhRFGh/GkJsiY2YS2Ump1tuAWuPN7vqFV8xeFWuZsgcgsPef3ly/
hd239Mxs3xb7KjXAAQXhLpE0pK7rRqs6RrEvQUP2AfpLq65hN+X5/wCkUyLgmzhXFJ20jWtfBxpd
1c8s0Ff1BUJz1H4Eg/JDCfg0MK02z7aasGzxrUzMH3G6+yQp6HyszPKYtsGEXOvcCHkbDPkhjp9l
qsG0RfRem+gHfKPYXnnvQGGJ+PXLT6WER3QExzo9SaM7d7PYqpugxPdKfbAJtE+X4IQr6q8vPwn9
GU4eUJCkswp5JIpUYTxLyGmGyME25BfzvnnyBcuInUZT5iWNOXu7rTImk74T7a4U53sTBDZSAH//
2+LSY9Qpani/Zvh4hXNi8SNYSLiSwpfSqXB1v190LT6/Ja8K94sWL3Zy/9+ueo9rlF1fXUGB2ACY
Gwfde0ZNqYlHRtT9QRDxg88Yd+VVhZgRRsPtkiaTj5htrYENiVnv4Ch+SNp8MKH+oHFmG3riX8rF
laPM6KXL5Yax6ZAcuiDs+iddVJWyd6Ds6QpAqomz26nB9p2o3TaN+Y6LvCF+VrTdN2TNrTmHg9c9
UotqkQTIj0/nhvoFI0r3duKfyjDJw0HKmuqxdp8losiWtddlbRZ/NfuxENIg6mx3k8JwuavFsMbP
ioE3mzXdR5yK7aSmxWaocjX9ubHxbq8gyJ5TN5cvRax5CRYn4xmvsv90q6MsOmH2Y5S1FNhywTzc
VflRlFNvdc+9lXlInQvg5sVXkvpVIf11TpvNLqUjCZr5fgM5e2fL4Tz5R+uuQXWDkRJAnDN9PO+/
P9IHxK8ATT0ztDW20cm8hBNdid+rKjwdwXJ7agLSGFcMVd84+oR/YiU6ew2riJiFC3hMi9kRyFSA
r4t0rVauUk+Jug7hkCyEwHeXnA8dlj/GUiNFcM0PfpVk4iRV/IyaEvsRhVch3ERq1GKRCYe9yTX2
qH8yDvA0OCbzS9FU6wFaQNlM47Cnz+CA+UaYaaabZ8u572ZwD6e2iEvx6hNSixuQcdFN8v3Ng4ID
JaA3mGg3CgbRRM/10JoibcHE1d77DaV7qvB8XaPdNGKckSYHZeADMtxeLJtHh/aiP/GwRrK44+Do
fI014Efnisu4xBgyLZj4W5vwh9/6gqLrwNGgPNiwGjd5U4BNp+RfvUN8fFt8BmINEiXBmsTP06Wg
lmwu/IAMdv2jyoFHifBtix9XUUm7oByTKg9LxX+5+EC94wPIoE1URfEeh675psHPO9sjKZFZlu9U
a8oOk5CHM4MqnCEZBylvvtzvQfh9Wyk0dpoXsiOLU760cIIZzRFt9O0/MZQahMhoQ9hmN3usNUtm
9HmsPJI7Uzft/3yyQruPIJWWf4Ho6tviNxjQmfKafFuX86vcgZxIk4IXElIkd/+MNN4d9pnZJYFt
dDE1OmErOgeMRQrRA+zVXHgbrc4shDtkgi5e8QUAqPU44Ooe42MHRJ2UEEN2QoZsuP1ghaD9/OS3
6nDrWLP6kjOLXucwj6WLqAhIi7ZWWmDVAYvS6r55+OgM8Wk2GNtRYFlZCexNraH3b6n2jNBi86h9
WbBsXCcs6D2OEVUoZPRj3ML2W+GsspyY4XnSs85UQPI/pMktiNwbw0xF8L8NQ6Gi1FAz7un3ukUI
SOC7zc+hmIjAQosk0eJZqM1Kmq7bryuNCeIoHyiWD8oqcfzNmN2lhJueMYnVdXgZCDP16+8WjNNC
1jpP4TBB5w+K7zGgddjHyR8Wz52hGgO0dAtbaUhTxRo1f/yp5miK97z248ZRKnYtCwCzDMvpPl1c
NsKAPtLaoBxKMYxBgm6Tvr7QwUbD5o9vWvZZb2Yr6PD2nQg8H4f/S3cfeXXfjAvzsVEv3QxpVLr7
VFrV5xGl0KsVMZ6DaD4JQuJG+dkB4nvyTUWDchyRLqdfGAcOg0ia0lpSHmPUNw6xPl5Lcl7wUKUu
5XgKFuKsL1DLiTRn5gcJeioKsG92l9nG7tqLTh3pOcrbOuNMhCV3fFuqiM23QZ8idNfLZI+JGsXF
2/DdRzoe78WI25GTBth8wSuR/uv0XYNz1miYiU75mTuTPlzX00ud1CNht9AspZYwUcl9HzY0YzPj
26B+8bCUgp+dgPqJiRZgscKPgmwTpuiTmG2nEc2495BqorZjcXqIkfP8axdno366sKyxBAsPB0t/
R83mFVyTpYn5/mcFdI3STuZPIfewpc4EHfTqo1hJzPLz/V9HCgQwFBSmhLUYEJ1dQH/yILPkB9KW
klIs66HelF2mrNuEIvKwOjfN5QM6qnHhSVkyH6R04NTrf/C1Zz7LkPT9oO7R7w8Ke7vmdLunf8dN
GsOwuY+vlN1aSxkFCD9cIAApWm0mwl6DYIA3I/7DVCIqOLXhGGCvU0pkjAqEYsyarUo2S7AtLM4y
m9JTeeoWb2qjN5ZIzgmFid0BKNjmN8HcpZuwp0Q765AA1HwM5Mbge2WR4dD7hhFPrsUCaqihsNlI
i2pmbuY1ZwxuFp6DidVZlU4iNw3f/XhYZmaaJ4i5TrxYLAlBSd650xHNif7opUR9x7OV8EwEDqPr
IfTlK3ziiaKvOnoc9hb0zq+6zCdFHeOyvL/RPRfJZKCCnl5aZi116EBvhi2kKxDxIIs56sUpwwJI
QywxcRWZnjDksSD9ecewYIlq+2K2cWFxAkLXhBkKRd1wQ56PCmiTsz6i4ekAy4UFg364vHr/szlU
SZhcHJUIelmcmV3q2dAYwl+kZQ1gUSXzGZVm7jFgmFTQIGUr6aoaz8nZVFYrM1NMjEcdYACnosAQ
YTvum85I0q+Iw/hlCjJbJXkvSIyw3XX2T4Kul8mSVq1GQQi3Gk3Y7mEzrqHjtzTloKLzDie2KtSw
A6gLAWUTymHn4VPxzFl7TwBAmqFofc519OU639PrcxspuxNfRR9PK5m9p0YljRAn+762q/6TQ6Qs
vPDj23/rJbX7HWfzmBlF0ha9hl72vaOqesfN+ituXN6wF4rnz1Y9tTyV5/8NZYkllfxvkBmtZ5H5
iDyJsKBggDRcP5NqMv4Hg6sHSaat72QJS1HM3kL4aDPFEasvjrNpsPpKPySNaby7L2BJv8C6IsCK
y1mQUpW83lmXaxfs8Cd0lUpEJ1mUbEPv06KNKPC+Aol6TtUl0qwLQkTEI3Ui0AqRu7UzTguX8wiu
Hr0NSgUoNsAoBcJ9OL8EVEw3HiZFnNpU7p3Jjw8t28DmrqpJuvO09f+dTlgMKt5uXtzuKMD+4dU7
VV/gnTAJHRKk4oMMTQM32GMI/iMOjuiMtyAw7CY3sz8JamfJOeJtqoQ654E10q/Wpsfpfidlz6Bu
TfJ2rojFqlco8ytogDdSEx15MozD6r36m1Y4ksklCSv78AwDd8yW/K6f4mpkecNHbbZc+bWOg9GU
D1bT+TCt8orKBTboo/G2WyCTQBxZf+fT7l1FyzGziH+YlwZUYjA9S/BV3juVFR/ckUmCkHVj/gY2
508T0c308SM6mDGOsICbcTReVXpTcUcg2lN7wg/HaKdGPVZCjJmZFfr9hd8sewBnnJoyEKBc4YmT
Qz2oSXwsiD+v82xa1SMmVE7p/2m6byOu7NQe7ihDNibSH7Mu0ccumZZ7ZC8tSsNJwIO7T/O9R3u2
CLp6IhSYatcnkksXuWnppTBIRApk2n7GNwoRJ/Ku2ov+/Jep5njCwrnB9ZVVBfo/T5hlyP89qk2+
8cCIGbeKL4XNt12HDizdSMeEE3YbkwLhEc7Tp0FtS+S3v6rF7QmmeDqgJQWDaxC1X3S7dFOuTNqE
7diP/ztqfdpdtWx4bfO5RG1bsX5Ec8zG7YTTiY5FDQoSeYDgX6a9KKPKO67VGDHGphoDoNM6TC6B
oO569bYp6Bisg1QsCg/U9LWrtb1D8pLRVLnG7YN8wKeLPfAUeOUndBmx0oCIL9QGMMRkAQnKPqZ9
AcxuX8Dq8uBf2xbuUH28wbV9NwaLs+gEOg29KNyEa/5LzFHDNxU70QPnkcyFRfHv8TiLDjwvrCtL
dcvydgIUOFz6HHI8gnrslLs6Q5o/7A59aEPLBaslF9Lk+GKkZ2eaGz4hBV6vbTYA6aWbppfuBo4m
rQNLEao+x9Z9Qu+3ZwECEjo40IBH3v8gJq3D15BxglJeP7Kzto73/o15MkALyDIllsw9gsYKXnF5
OOxi95bVTk5Hq8kl55I2If3Qpd26nTHzqkDoA2Eiw2bKhAee995Hmh7DxhxDplr+EM/Wza4ip+iT
bwVsDKnB0sE91PsAKOHYqiYohSWj50CvQaHCfk7M/SQlXi+jwmMEe7pMUNOzVQ9Y8ubU9JyL7Uzs
QXQXRvL+0MN2pqnhRdhWsoO0ifKm5qPNm4+3ZUAmRnsOjagA7ksUnK0odSIVwdiH4lZJxS2FHyN+
dQCQKjVnCSc/OVuP8sU7DXZKBJUsijgFnBocu/iDPKliFpIsbVoJfS8MZAj9x2VmxSUVAqaElQr2
MD7xu2MCq0vTahAR8YPnbDjZ3dMzcjzlh28tPPENguAsJIjJbDiTAWlfgqNsMIR5A70w+/ac0Uvl
/gsAZ3EAAM6rxl1xH3p4amvkA3e3nupmZjzCXidwnz4dMqlxX73049UyMxIwvzhzE9gkFuBcxOUJ
2JsHpZQF4W23aRyFUiZZLcuhvXAfpXnJo/l3REQmjSFHpy7KxU3aBiamP6OkusL8MPRNVo2c13og
mr2f0O+/NYQ73D6yito523oV72VaXMiTjjzP4AxqzbjT4eswzbf/ycA4v1VIH1vFrd8yS7aeljX0
/tmVx3MU3aN0fkGLeMQstpT3X7m57CXuVbyHSqRCbLE3LeyrdRARZFJI06uom+fMGtXI2HDabzxs
E/uRqW76cqaQo/LA3xul/vXY+D/CIanjCNu26Q1hAchFkbew9rj1sWuJTACaXcDyg/LfLx2K5yFa
LtTgQbDXnuSqw11l2bLB1j0ZfYMCZ0Njcm4IPkRs412V0Q6jPPgKQXn2Vr2Qhv4Wz6MXGDfDmAWR
MvLtXixe0spSX8uxZlbSTws4UU9M/Gjcp/5flE8s34WorQGlQ2ahwFJ7s4MwXLtYzNaypX3IdDP0
Pe+rRdJxWHSPCmFwYPw/IlZ7C29dZ6T5EGxiLtj0TpBUEnXJJsYtYc9j/pGHOVwfvhqBlSA8zCDj
f2fzC8x6+9rdEZ9iGOarFxASn6Ml+NxaZ2swA+SLfaXVmf4awmFG0BBkTNrJL5cX5q3HKKOYFnpL
+UZiJm3of1zeZRxu6LtK6QPegkIOQ5zdvYwMggmBpTCRIAj8OgTHY8THcvu1pEWN+tdZkXB0s3Bn
GcKCTVKh/EfEt7cidB5cBVNZVleGAFQDNsIXekSQV78h+0GwWuo98HB/9WFxeWfImwBQoembFaw9
oawFFDVlQYvopnz2f24vcnCiCjWp455CHpucoTYw3mlbBDtlQ4Kabj12p9B3zKKDfPOIIYu9fwOm
p1u0/CZAa4GMDAo/++t2exQIhAbcTNZR60PmsE4R1zyrvNVKwAy+f6vq0hvHJsst2pxI+voh+/E6
T/tdD3+W2hijuADlSIhz/dz9Ck1Wynzb3ILTGTdiHeDWoORd51YxyRGWOHCe7koo6vWmk5rXHcP/
jm9w3b6Dzk5UzZ5KSP0Hyd7aVqJULlUghUCaqQZfyq8vc1me3Fz65BWCgv6mPtrOjeB1dmP/qQYj
QAAZR9Zs0CSuXTBcvBCEjZpdxEwln4K9fOSlE3R1F1YjW7pmxN6el3CKnI+ajw9ZNer4uefCozdD
AE1QBnt4HZ3ef76x7L3VWeoqosLbXKW6oQ2uh3YE/Rum28wmkG+7SZHcjrNWvSX8Ark052YP2EW8
MM+FUlq2Jy234SbT7IkXseXE0BgO7a/qq8oW2lKmY0ymfXmvLTKyOJbEBrQ1i3W+jcqmvGYLxxkO
+tPNA4LlZv52fvk8cSuIM1pwJzLXNSdQ8nxaOKyalhDdSJWSmdYpW9kfpMMSYdtavV4M8g/5SV7E
YOPux85Q+8wBLuPWkl0Y142cBNR7QKGDJMY7nhrakW0wvXlGurliIYNf+M0QbfISKB5f9t7g9JAU
96w0MGuPjE+ANA9ZGtgYo0Eajnl+vO/mPsMWtEtNifSKxCV6t9/AkH1HwN7WFltJLmw8x4AYwtZ4
ZjYnkfG/4XOb+uMkrPiFUmDe5XiEIFbLujv8mP8l0TI1mAow2USt69++Yot7fw/ZF5EMlhj8e+YU
RFTRap8GSamzIuIx/pFox3MHByBJ989gopQ85j4/RjXBIjjdZxYkpGaOTOL7FwO1pYCkqLjI0smN
XFsmvRITwJU76NZTdiUQJUPFhV95lNq5eOY4c3ts3AJ/W73oDUymeLSREWUPtorz+UmV/BF0ZmXh
Fn82u7KZYsz1rOLMlrAGH3bPHeQzb4Vkfa4ZkPg1JK9L0LqVNJBsqubDIOvKuePnRLgKl+I9d2TB
bZlkI7vRduFOynMelvO9stdsEguZ71tQ6SHHSyLkyeoD62mkOZfvU6ROf2Nxq8DQgJuyvjr6NpuX
oCHXhrS+JTDoI46NgqoaBj/+uv1O1T8l2rE+l8gFd9rD0Qd6T2hjizS/JsPO5g+og7TLvVltkWVc
WBTkCgJc59ofBxW143aPDRDegrBeMB9V6ho9NeMprviQteApq+o31sboBl19S8cITFchIJHuq+l8
p9mWYyqQ+mAh2iFCmEU8Hc3TkFexE0fKmTHofASOX+2MESi7E8CxBNCgLmMmB276rkXS3KvdsxPo
uFS6Qz3dRl+ER0WDFXCflrBlv27+OBoQt6Ia+FbCHumy8wsoR0tdnVNYzuulJiR9+S+ayIiB09eE
+EO6bi4FD9Mlca7bGm5jcugVRSUD+NlH4wOKIeyqySuxh/puO7RsDoqilnt1F379Ne3r8j0ZwZJI
AKmfl6kEEGjOISPxASgWXKBw0KOnEy+/nU8R7ZEaUjPwW4C9WqprEiB+5uGn74RmfDx0uK/Z9a6p
N3+TEKR01LvXkbOVejYXWduwbffALETiNve4Io+aw0g6dWOe+jydzWjJ36xn3Bp6DtCsAnqS3yaP
KiRNhAG1lJ3887/p9Fi76lZcIsoj22+nzBhRGmsPFWEAOUvC6RMJuYNXva3zLlTXUYLHWJ30rbl9
5JYbfwPzf4MFCPVcVYC6m4p8RYEwh8QfZbQ7hD0K4ESHWoTJ6iFmtdK45pELJIoY4eskL6+t+cES
sGG/2IGoVY7CTCRR9626KiDrvx4oTEPdr4u3slH4Mdrabc5l0KRIn9Mi7dNi/r6qNFbQqMFPjgUC
0wcrObUsjiXJA1e/ht8HSGa0WBplP3sQzAXovI6Vqh2iIbhOSJ3xL+gWM6ngfDhJ07WJ+Fdaz05a
h8zbwO/6iGT3+9m/UsndusywEOzPoR43Pn1mnh+B92vNwccq1fWbVMp/admpZ4SlEw7NiihyF5zS
lbwFJSvM0e+3OmVvCB61eXn/Q9UbG3L4wA1UDRfSUo3uMDHFY11bMhbokDvhXwFqjH4WjOgs1j3I
Gc1QrvMr7U9p3h6ppDwXVqX3+JOs4ntqUvJLI8VM8q5xCQJ5KGbHjsotNcpVGM1plKohYaJ//smQ
E/6Y+CFB+zaRCxFRXNmKz5Hdmn0cXPsVk6HaTJ8qgfwQssOKcWxwYb3d0oAR5/hJHUx6t3FXWNiB
vLTA6TmN3xbcK1C7d8bXxPhUEi8A4IP/klFUYh41loW1gj0CkWSfRnI6kXEc9QlInhjEZCyLC+bM
y+qsT7FTVDl38NtfRnoKFblByY0CQknYa92r5BiVhavMAgItsRDYM8ARt0MoBzR+sEdHsL3rr0WU
EzoM9FmT+l/3S9XNdwexhAdLratwvPSh1h//9kVu84vvy2pm7sghkz5HbI187pZoCLIZhXa8MnOd
QBtV48QtBMNZ+elGB5vwqpsqy4dl15Om7kMan3n2+4Odf9GbLrEpMXHghzY2PSQkzxoIL0UbvJVT
bESc1u9AMF7X1pXd7oxwa5PQvb82VgM1zeMBi2FB5XsFqGNbt//rB/djNvfrSrYQLFcMkogbFxDc
P0KshUqSVG9RiRQDMj84q74er4MiEy3cZyJwdtDLupO+7oO3Fu4R9HMtDgelGQ7zhNmm0W5P/3gx
hZlKZfE/Pvvu50xpIdrujQL74iCD+C7QN7D0JcFVp7ctHGvfwtY+jv6U9dn448i+VI6fSHOziotX
weBG/UfPOl1SzVhE+cxxv2l/BupY9v+LVI7KRcb9T43d5F/Q0lVjAGrB8HxCk5IQZICQpvUyY+S1
L1tsas1fdbe+24fruTeBm2B3/bUFqarWU4WMt1rYJrEDJGkDq0NbitRyb4mSBHksCnprL+On3yp+
4gWgU6vOPu4yWEavNys5bSrcZNKFizm4BLdZzJHTEymD1O/0BYSdRUAd7z96lKVPDgoNIyNbMsEU
RKks3g0NEXjnyBd/PuoQECO74Xo9vjg6blUFQliseW/ugET2Gf1LgJ7+3avSgOaorgzbRPyHPWg2
7YuiKbckJB91W34TPN6tZnCHrG3eE+muc5xaKLnRG6oW+oSrcqOZBwfeHaAFRV2cQ5T7HFtnetfz
HL29eEPVWml0Qw/pq8UpTXibKyG6Aj/00NtD7R2AbYcDEh/+w3dikRZ6bHe77uw4ljDPxAB7QM6a
QBtDx9Tg5mbY8dfgC06hsVoZxkv4nfeHtakK2Yeivm5wm6bJFN+zikOwLqQHGt1uU9UFPqadpVu5
sjJuwJmGQoLM1h+02njATlIrcWHsPiuW/880brSodFpRcdVphkzH16/hjZhaWuJembEmN3HQTMcx
j7YVnm6sNMuKrw7NK2Mfo3m4IaQCtEe5uRrDUw/RLZbbkMvKbpeSqcpTSw1ZcyoTpNmvoa4epg/V
EtneQa7VrAfHRtJfJZ65pZspmx7j8LZI/ehmdK3vhjrEM9M/AhssyozB1vjtwMc7VZ/bUiNR8IEa
Kc7oKhHcFxZm4uT3QfiUJSC7H8pSAD4ztGr/IdCvmkuJoUQpdNwJPaVJtxiD3d2NUwYDOdlkUZz0
ZJGhMChYpy+YuOymkK8KX5M8t6eD1siJt6aasD3Z+vLJTWY3IfeE21iey4P0ZeKp3U4FSvy/RmDR
50oEeYcuYaUpUhI1q+RP0fGhmyWYYbjCpD+K8KJRLiiQRLj1SxXXAJcLCaJZOffEaqMDM33euZCh
pN6kma574/q3cS7dKWprf+AQwBxAwCNil+IEbO9eQ8G2ZbS10LOYDYtWYcJ4YJz3Z7ZAfGmUStGZ
jgr58xGZR7gBQBAfmrUZQBpxVDzFkmbUqbNEcVY8j5Us6ap+otTyyjSaiC4PaUjabcBQQV74tgSa
rvq/zxycpqaj2z40Hn754i/iIhbCN38/p+ZJzdqYPNQxDaSlN/ilCLtMgXw0/P6AKnI/IUXxFH7x
Usoq/kFWYcb5DtWK3mnPlsiGoCFMMyH07HzQySOZmtE0VCzu51xRj7e1lgLpEdMmKb4gQH9AySpC
PGJDNNU0WMZuDXaFKBmLZ34FZVMgLUPYg2WGp0L3H6XuNrCw2lExT43O6cdx+Tj0d2nM9dHNN58J
fZab9kZouzGN1iHBuy8E8VZeydPj/JiD2v7AAemuW7LcdNHgZy3O7dPCb6wV51/Ny8Qm40+q3f7u
FTTEXTMdhXGCc5O84zpK3svaamUpOx1eAFqekw+2IzE6JhQPvyCV1Og3Wqz8d88wQSAV8106qZvC
DemqS6Zkr87pkvzU57h4ZFrYW7zlK3z+KodOj1bTlrU0k/9tsX0rhJnyjMyd6JJJ06KfJAMIvc+3
PWdUSULJeGjtoaOFdsM5a2FrpPkqDdxelhAqGfXQl8nMQzbKPtNvhhsU6VXtcUlqMud3mnbXMsTW
mikIAuJX2k6IRGOQUBjXCdy2UjJQ9XctwG+BdRYTRwz4+4qRU+jsWZp331HG26w1EknDhdbCPE+A
dGK6NOev8qyp+FCaZvh0tnOFdJDH/uZ7VKxzChm4FlbbOvWEAsS0ABrE4HKHFC5OG9vc5CFJbHyT
t3daDZILsGo0N4JQh6hH0IS2U2rcpAq4N5D+lRymGvEm3o6QeJQ8dTE1CF+IRrhqeRvX4BCvugnS
fZ2Kq22K/n/q2o6qJvYU7GuH6gHSultET2Cg6EYx5OOq7EICORSws3B7rkKVImYbr4StINp8rp4d
mbG21V9QmUrIJC2JnGC6Bfr8tzIorECUCxSXsyy7q3wE68h52EsmSXN5w/wfu9TKLlZvkm6ESFmh
nQjaSiW7W0cZ7BbgIJ+mWdsDzvufqxp5JQh0dnUCnLl/gnEJ81utCyQNImkmxb5yVmz/rGU8kt/3
TZnwJcx+1m1W/Kp4chxN0OpA8rGfOaUGkHsFMGNuKfsay+u3+6JFOKuUKU6PHr7GB1+mRHT7/j8s
5ccwJrGH/eMv8XhNlNr3IQazTVXlqtCx4E4rYRBBXYoSpUjmOb+wkqUiAjCFj8sG41O/gnVJ07JQ
vM19xnRvYVLKhd+AqKk1xAq0w9lxTVDkCBM71xmuxXU0dCUIa64qy7YlikMF+Sphc6Jiotce30Ie
rK179+e3W9iWf51h6Xf3UxpsVPmZ1oZ3qDnEhBTdyNNkbM7OZa6phhcxim1OMFaHRW1YzNRfSBEq
0Y4DER5V8IgYrCYCsoupbVUG2iHVnlUKL7IN+SqwqmS3CFYBZQwCYokViji5YFQge1XoORyLTvFa
Z1tSIM5sX4GahVTEQ9djUQ0xIC1Be08u4070oNL85wbeTEwXz2dQ5q/Sculi+nz1p9ScOKHAHEDE
ZKsEloAYcF36SLEFLZNEMfGzrQJReZ/DCRaSZNNgj8HRTTZ2CImfKz0tpUuvoQteM6lscEzFzrOO
mljWR+k0byFndgkojLcRsCHNknfeeYBEk38T671u6Jmsfq1m7Flc766vPdaCUBjm3HEXVwbsCV2E
Emvjp8nvjAooRgvHKaAiXTkPbZFQ/W9u8Pc4Y3HUdPLkWnrbq+hUV8L01gAop6XsP0RCHwcjGOrs
fTyI+kJk3gm2NVbonPo0cjZPwjsi4R5Zo8ZbYjuKQpcSi3LjlCzpQfmGQItbZ2tVlkfk05TTEbWJ
hHM5JF/qLcsX99KQPxSTJVRm8+dyKSfbbqtJL8HAGo7naom1cQthdvcSwribZXzyOnCoBa8NH2hu
Nlr9+LJHdthgUSrZls0FlDvZ9AeZjIVtmP0WrjlMl5hY0rqYwfsIn+g2rlsQhERWXwc0VAV3oxN3
Z0e9vCxG7hTCYKDv+3+3q5bpHyepmZI8NjTiN6wWwYIpUWtA8dh4WfrWscsATg5jPTqUhlEhZ30Q
mbJHDmp/8r38NAFkY4Bj2lX2u9L5GXJgmsv79li1nv4jZ0kQN4FgFRBVtM7Q4B3AfPDZeRzsy+Gv
1NDL332neqx9Nu552gK9V/cDSwYGyYt8Z9gksm0sEtpXZXdpZt7PzxNoo3jymxcLmuHZeLeMQ1P2
+nQj4n5IZDYvWyg3PkFKFbnhc3R20eDFy1poszLtS0hKgnCW7odBIXcg0TeiTyPbl+ZfQPbPGhJX
fW+zsXfiYeVDszmapQzchm/V9AQb+MMJPYuf5/KZ3ur067pcgwmvx1i7R0B0UnmqpnrNWPCsJBRI
JIvWqVO7Emh+TPhVujLHMZI8oM7LLIPKZcSQR9/pwJgm7Dieoa1UX9po751C94EOxpB7rYtJJFfj
gSSRcN6tExhIo5FvGapzB8eqYhl/qE7mQcATsVBOGb9GFS9nnDxnppEMn93Z3y8RY+oKlrMST+yy
qym0MiuWOw65R1xF4bFPloDJQQp//4f9sZ8dOPu1WQsIPlH7U6TltVpt+RH5tz6KiSxl+3MQaSI1
aBaPe1yST9iRxJDQ+g9RUbgDVXPmcI+qgbnOOAS3e6onPvEp7hJn5b7ET2NqBWJ3HvXmC9zx+qle
cgvKv0CcIUL1QLmgpTbJ99ph2C4Why1RXEA8pXItr9aW3UBmU1GG2Idk4dvcLa7aHl9Kez4+vR8G
dITo0FTF7qqU+mEIXpZHC/nGPt5w0lS2K+/B24C00K6dQUH1fulNhW56U9ooDMD5yjhCGljt+xEE
CwGKd+MNjHx8u7cs456986DK9xFpdpu68g2MOnj2cGau16x6I8NP/TpmUI03dcz6tM5dv4Bg+CPr
X5fD5yy5t+P4lCSBgb1xccnWD6Wzgh7pd907l08lB3Nd4XMcqL1xlSkdmdl95msxcTv0YVnmmZ4u
VkP8pyb0p9blgWdU5/V9Ygbd12YT0HY/peRTRtt1OjtDNM5w6VGG6gTpuhdVcGXv8PdbazLWTSIF
ZdxTGQnAXu0ozsJOPmzQ+QeRzfTUYkqu7Ow2Q5nP++74RP/prsyy8qEb/DiS3CM1EgMCe3y2AeXo
WHuE5eUPhfr3FMVOW8/+8+/GE++ePC2CIgcklGxDc77yCFYvYAt8+oEB6cOSTcvotk1qMrOjQTXO
iyxj5RXuBC6oG7D9POxSYfS6NfSJTKYCdbLshmSyK/gOSCULP4G2H9nh+VhYElsui4hsnpOKBFQn
V/F0ddmVGDNvw0nqHbilcMzRhyD4yp1JXicyhe6Vi2CxOMwhub9C81F/ScamCMAZJ5qtgMGRr69y
TTWlj+FoaCJaz9/hgj9gh6Ym9B9jevjLOCq5fZFRsg5ITiyIFddIX8/Ksbs5DkN7bygKzp7UT1Ky
GDOUsqSZ/HhjJiX1zu98KYAxOo74AihNm1Z311teRwI6yYz7mnnF56YRqCfZ+jnG2oe9g9yUZXVa
3Oy7C14Y2C2UOArhizVUXqqGZpyamhKpNnFUL3jqol4tbUgAX9P7HkHE3KaYCKoFLnAQcYS3UUq5
Ojitai4m8qQC4wQGsMQHasVRn8kwh8ruPz2FInz2qXFoTePIXk55xezu6sbZTpZJXq69xMzO+cI7
jvXV+xM9Rg7vfXQ/O0btrm69oTrzMEcL+dH+0cDBwamaK7qqdID3E9xrNGLs7W5sZ/LOkR3Wj66V
H+mMAaezbe9XucFjPGdedLsEWAzxOpT86rDXpokALkNZ3IszIK7trGcVnU6GAFsspldcLrb7OyKZ
gSSatwRQJzSxXP9XPFflQw/BHMqsHEVSid6iVrQ+BzcgUIZ2R0QIYYygnyMVy8RCXqMeYvf7HgWP
1dgkS97qRg6E9XHqSY0A9GYuJwuXBEky8JT5AhiYu4rzAep124sgZsechYc1LPfC5VwFGAynFwTU
GJaweow70hmpEtuY106MYQ4G+6fwD3fXUIF29p/wUXr4y8p83AqO55BESHrbLmqMgUwwk+cBpceg
aA+byGrP8mvNT6ilD41ENFewQiM9wFL1O+U0s+9G7auqoi55qDlGLjJnXg1LHLaLhzfudAROEFq6
4gg2a7mRgbwD7ldoAM01D/XGwoJHASr5hmx2+4LU7eN/2qqDqBXCnmx9DFqh+pm00Fj3seMWshlp
L3a9bD3qIKZxZENp1klmYNVULWh7wpL52qZJTR03RD6Gx+Y7S3KpqTlgD8YvU5ozBrfdGXJhuoQ0
hFJeSCxxGR5VhC1rxNhLvyEw1Fe9Y1Se9P58UuZzq5Dp/LP3Kw/OnNgr2ORt0oiP7dpeuY1NXHDa
VNRaT6r2OVP9idnJJ3xjc+sDDssEILHN1y12XjZrgvi01I9qMKXCP7lDCyK1DBTydljv0A8hUxY5
xtjzrj/rEO4SLI/IPT5/bcqiHuCUnU+6I2eZK+Cd/Er3fGd2DxFfSvpcDDBfIl7FluNSQtRiugPi
0uFWweR+wEE+KI0mBqkGNuEqJtSIEEdEZjnChic1ElQt/Kyf2DDYfgTIHvTGPvm7wF4bhV8YmPCt
7+1jPVSRovIoBg2SAsxUjFjmf8nFA1ZdA5BG6BB4VzdhV6SVoQRpTC6jQkPV9/lr9zzmHqZObk8L
zSHutyOVI1bIACq9WqAIr38LfYLH0BoaVtCclptUifLA35cjoDag6pPaTc3MXOjyVCC6yzDzuaUh
DupMCvZtW7a+D9qNh4Sltgjz/O61rvP625yZkrsDQHXYx+O7Nu+MnRZTuOPxKSisNArN9+5TtGhW
kG8WRc9KkJGFPJzS9hKXMSWIE16b6NNcQWxvy7+G/GFx2jD/67G7oBKFo4zdCMk2UU09ruARbJJ8
q1eMCg7psEXNcHt+l6WyT0rtmRBgp4wJfL0+CgYqb1HsRXjQAj0ELDSA94r35rQ3AgvCUBKvwcVz
2AZ/8TpgwymXMyZTfTBc6wcJ1uMawH1uNhzA2KTj0LYBiyV5lb0RualJeym2uJTaqW5KBTrojocJ
8rfC/K5pkGFrw/bvLEr8gM5mP8loYz7847nD+M5ZnS62K3s9HSwlRcm4c64yHIrCjMOyGKX5dUz4
qoc/375bVfHeUnIpWJqZ59S7Ci1qT8Mbm/D9fHIZRWelXVHfrOSaiQfrkogXr+UIraEc2wa94CqP
aZDSBbKLnsAhhfZ8bV/8fg4uaw1uExH6mPb0NV1jiGqIuS2RLoKi2CMEqPNJa5nmxAlhGHnZ2sqz
6Seln/dMQc5OYbEs0w0vHIA6LtHXgj4X2doYjxJarV4IPBs8DhpP8JFqF2F6iWW83Y8UpJqtucgT
tbiCnV/gauqaFUuDMz36nK2rpBBm/aEluglzD2i+wOfewfHwvljgtiRSTvwR4a22ls28P6ZrR7KZ
QMeQcmwAhIKbKaA4Rq1/kZgxGRb0BwFs66+E7QpP2EGnmafghzlBu7igiZja3MJyZ113yeNSOMgm
xcgnK6miX7UAbWmc86qZOvLEGH1vL3kRaZZaPVeitW5jTi0BZ27Vn3pfB4F4QAu+JK5rNikLdYHo
qNhskbPmn8Sww2MHmGHs1FVvpi+KZyzpYVfhcUmCnmRr9OmqlSgOC5NaNmXTVl/1SQjbHHR77wN2
MLn4OcQcIV9oeHGZ7uuoo1c+xxb267hmOI17WmIqoM7N8xCZUi1H8fn3kD+pOhjOqlKG5IqVD8MT
+ufzpEUlTCEtGDMIr5G5cLm88789l2pzFfBV2HoDMV+bN8GkgZJpP0zTbblHrtkqzJ8V+qZFCbBj
oavSOzqlXVyUBW8O0C/sp6JOzSYvVvEoPUpRBa7icBvBhVyyQT+BqbgseQOgAIJD0f7yN4wy3lLE
uhRn0KrpEzy3LOAV7gAFUy0RKwup6MOm4xNo/j1PxyS7BbjJfYijouyAi3uO1DHZf6CpqK1EEn/g
ix6aHz04V0W+myFFhLeC3MXe/JoePZQfljJ4QWxHaXCPlbJy8/rVIzP3BvPitA7rLvD++YsVHhXJ
8+yRxKhBN92Km80cDOZADeBdQqOFTCNuzbrP/smnr5zTxWxj/uJHfPcjfzr8n9EJQVBfPKuG7sLi
roWCsDlWQm7hKr7VwZS7b1w13M9rlBAaUB/arZZJ38mwrJB74VQ5GO6ikRtxT1en0EAdVUv5Ene9
unECP4Q/cYmivTAmv6i9coVPgHXtwjnBzPvIq3Sr0dr/IN/RiqF2AqVpOaKnA+btPw6ufUw0g29u
ZQuYzjWk2IAJpRs70nVfrJO0s4o8G8wcHyU2NIJkDbg14T+UasJ1Iyrt+J/gPsTq89qj7ximFGdy
XKz/7oLjPAgewmLwgTyA0dKy0zrrT3TebOXgf+mcQOvoyB4AUg1r3N/vl6cMbfYppEM8Qrcslhip
M/Fr/lDvtePCF6j7F+BcflSisSRClDVNRvkbC6RKsPoc6gyxSZ8CpndpFFoZ1aZAzYTR/79fhT4u
kGZ6C0VcBKSa8DLbbxT1tpiX2OgGu+BweJMd448ha43lr8pCytMetMf/KdI2SzVp1hN0z+Lar659
RGfllB9x28sdAjsa72TXw6XDbipwUpvBY0ysYNxlGEKP8qrXWgW6Tpi0UjGlMQWFFQP5IzD8N7DR
vGmxvKk4/VRX9Ck+ihMrDnYMOZFFetj9AmyXoy5wT94ArXWsnMkSmSVOSMoubuJHBiCMr5BNz3YE
ErpBZ3cpv9DM668dDbJjNAsZ4zVdA31hi0l4C42rnp5qwbfyix+3tWMVlFFS8oDAHhZnAEv9PX/q
fIqJ9OpwkyNYrHK8lbIVyiDz5I8zU+R0jprBNqtHFhVKQlbD08O5W/LqKF+m3uTqmvmS5o5HPYXZ
P2YnMuTTeHas1NulKC78I3tBaGajmc7L1NiKzIdEpFcLZojstLmomFHBohRT0K1wcG4mkR3C5bfg
RMzyhTRNbZhQS9myGhKPpbhXlUn0JBu+ncjmATiDxxpu1SS/IR1F8a5/yuOsaydg01RyG+jDrAB9
JL7XxWzZHgkxytyOz1vPxaNTuKL1Oz+9+7fZ8L5gwhrKSAfLqNlvmTKuyja7lwUcrXtgzMBGI6qI
Bye0wMwsoXUmHf45d5OTEC4Zh3v8ka8I6/62RLpjkGcRNKHQRo9cLW5+xGPXiB7fUAYcgeaJVj3c
on5xSmm6ufdVHZXOn2/ulcFAl/SvNn/3hMF2Gdiy7mYPzs1ETO7IcDEkaM5Znbn6bwexnzbSIu1E
4hYZmWvLhieE0G9jON3rbX07P9zFxDbKgRhvKzqhadBTeanbMcfUlgZdnGRYCx2VFXisunhfVDut
s+dRiGwtDvtvNMvKr1s6E1MajyYAdIn7ZJa2Cz1EaBGygSRUpSNsJC5SX3BdqfZ60VjfZxkzg7TH
d0e/xRuLKSyjfI4ydKpbh992GoBSoMWAXrndmWxxtrzMZP0LsiySLFnaEPkfcO8Uw8oEfMrBEkxw
wJ+or2UETBqHt6ueokEikqMWaBvD45gh9cmJ2hX24Yy0yhg6Tj45wKiW+JalgRO0u37kVYVy1fJx
aFSAb6Bt+/I8wu+E3+s2Fd3TEwzNJGSeKEawn0eD1qN+clMVacb4HLfayTHdSqEAOvPPZwhJ1Unm
A7rEjY2V7yGYlkZHQT4l+NB1IpjAb1WHK9Sdu3ybWmiSfboL4eGbxH+eTnaQd7I5RVtf2KW+Dkfc
fQYf0KI1wphAyfKOnzDVkx89kSPa7GBajNGO5F9wXBSY5LS7e2gy/TvWn9Ie1U9lSzh7ZZMlAxfb
OT8FAs4lONZPdfZW3QgJc466jfUDSg9wDL7zbcqv0RgP8FjJiimMQdJP+dBU2KwV0m9hk65b5lRn
BhlDWNJtKRv8aQARCw+BFgblNL8jBsI1A92oeiaXg+O9D5JnC7JEYBHnbs5tn8jmvR47zMVpvlzI
P6GyjBuxVrp2IR+mT2TS8z+czuaHPXfO63POfprGil6L6BkpdJ9x4ixqSvur3Ui3VoXnmKy8Y8YG
rczjO1qg1H6+uy8JAbbYuMsnnfHFky1bkNMmYy7avsix3CT1PFGCvKJZ4hKPo94frKgon7Ul+U5x
HPcn5eePeAoqQ30VIHwj3HabDGpjQbC1TmUlZZ0FeKwYPA3IIqxmkcZiuKsRiknzlOXtW/O1WbO+
LwoTfuMINiDeqUYrSJmHiyBMtu6aNE5cXZJJ6PkRFclrKxSKksEn2pOKfXL6Cuan9XCt6Ua9Mat5
GxMyTavGOMQqcVvqqiMrtcOJLN82mg/Fj8oj+o3p/x1l4n6KnHoa459hSyi02+SW5dHc9KplaX13
ynpulWq8iufZbBGm+S/JTq9RORcaQOvxO/Q2XX+OIzwoh51elHlzym+r6iNmvoXSPCMKnpaO/uxS
EI8yhAUi1DJ2dz6O4zmY3jOX3mcffo4MbciVWowv77qU8a8tXixFVK/NtLtK3Al/bLCw2BuGsb8X
iR4DSWRxJDct4TjRbBbyKilvEXutUh1c2WdFAJaU1AWG5tYWJ9Zow0cvl4bzPw+kQ0M6C+xvloH0
x959pZd+u8KtxX5vjz9QkhLitVyohA0HTwZsiZBGEnr2RETJBg4/XEXcEAf2H3no1LyNa5cHUepW
WvAGVcwH9JGtXFWS0eV1jCZ712W6O+Irzf8dpCa6HhuqXJtFOsU3IpLOm5GFkoIGnIhvVxU9BBde
vetOfqpgh3W1ugCnZK/rCx46Au2hJ68mVIus2qZaoW82AZnJrq+aDeHGBg1zsBQ4A2S5m2PH3x8I
zC1J/1AKWeuT903Lnf9TxtwAbRd1FMDbYhrKcZKP5+vd8bvG95MwAoTnFjTfDDbqv4t3IVSV4am5
teLYud+FAk6ejHfIHBmb2vi3xofhMRSufwhff7PcGaOnlROFvpnsBqdXxHnmdQZYMbvCV7E8R9ya
qAi1TfZ5i8pe9qUKbyfAHe9WTU9vQvGCWyL8c9Rra7xWFfvk1P+3ZQfXBmbjae4hwZK5q75RISt6
JWScvxXP6KUE3fFVs67s+gCwn2E+5HFgY6t2vcnxogEyIz+txfyA0qcp8yLVF0EKE8ijZX0zXKWp
vxsOypcRtPsh/PD99JqRwlJJi6IJaD/ppUXLK0g7wIfqzY2DpPKfnUj8NJwC7VZTnDX9WgMB3fLz
FnaQ29HqV/iGnaTFn/OohAEujvcHYkc8XslS1o7oCQyb59XBrPP0d6FhfYrYv4p6LHI43ULKZLmB
VAP4xZkhVeYDEV0IJgAnY3zUQ6M5dyEEb0nODT2z+2fgD8gEUB+L4y+8o/8/bSmn0wd7e40T8GRD
NQ2rFk8p6ukmXG8bc5++O7dq3hgkE8gVG4uCJb2C0iw+UCBriBNXL4nXWqohRd85vXe0MA2I0zbO
Puzq/5Kiwpa4X95uyRFSJ8UhRgoB4V3OAJALt6HS+Xw82VkqzHW6ZyTPL05Tumqw9Hj7lyfOEhXJ
LUtEv0hUeukVucjA5HTkUZe56z4YEvYExtLdxv5nJgCwtqNrjCOm9Ho3DmQe0lwTCvjlKQkitVDp
XIde4k91ECQVa2JV6fVhmM272AsdCAjcRYVAkOOezJBAeCEqgZZe0HkGdOHL64i2Z9qcAbibbsKj
yToXFHaheCaXUykr0sCZm2upRedMTE7nng+mo377U9YgnlKx2D04/AlgPRzB6GWWJ9ZICZ7lqoXd
nAyphopwNk5TN9xKy4S70llILRBUqcBwXzl5WZ0vCErgZDa4yqmHBXIPls2sRmqT5xvHoCizsQ2L
+KCKodk6UCDNYtv8ZXsVeQuom3chRX+GGTBXMIh8c+GEnTHEB/tH1UWJkABlj3udqO2lg6/lJfzD
0nINjWgLtcAzP9x0/s2UBUQcESLEukuTKKWIux3whRq4et/2aLl2s6DP7Mdg9cCIro4wg9gOM9Ve
KYNkqXq+Heb6sXVZffMOIvSmo7G3m4CniMaUImdTPHh1u5ZnFTpzVn90f4wMLH8mF67JqyNBf85X
tu59OL1CU3KvAT6L0QVo2s2hvYTHZWV9H2yvEr8e8zCW5XwIKpFuVM1Pn4ERGtm9nedM7PF7KVSS
Cu7/2gRvLvAejQabJ1vyyQ7sO3wGZ3g4Av0WlVutx/EEdnq0L+AJO03FVsbSPphRr8hAHbrrx+hs
AfOptwy4fpnJEfquCO+CXhd1eMatfKtY50BJ35JxLnvcWh5NsySrwf1aQ5WFdY/UpWLJdxsn300J
XULUj7OKhu1pm4k5e2Y50SgVMfSbXrJOhpJW22GLFWnBHFVS/rMsdUCtiR+YNPkmjhQY38rDDfA5
mzOLycvBGcEGIsfzUbVkqm8TMVnay2BlMoH/UdaT+Fa8XRMAmjA6y8rQ+Khx4ndxGOWCrV7RXbV0
JiBNuChlin8hBxH8lWgtXEPSjzGNJ35/UZ70SgKBVXv3SPAjPwFuNpoQu7XplL7mAIWNAJ+MYtM2
HfudPrj3LmBlT/LyuL5OuP4E4Da2O3lDr0mJSaOehKB2ODwPk2nRGEt+51NguJ0ne9U6NB2W55N8
xVY3W99nsGd5nZ5P3gUI4I6oRB1V3a78p9Dny2nMkdTepM7TOrjft49uSCEh+1OAJOwZ8o6VMqNG
Amvu6sn/BZYZn37Oz4FAx4MD81Awmm+VtS5+s9xNUZq9OMR4Ctm8ryphx3ZF+BxYuGaobhp4TEZo
r3jmjEBzWIrCpUa2e5KMNz1PkWYxKyDWUbLjJuv+8/4475vwgOtiAnSq7w89Ev+KL8itadb3AU7Z
QuWBQkc1KFHSGcHRt9BxEDkYgxK5Ro3Vb0TuUt8s2WrxvDWs0DITW5ur+Gm+ObEXIFMRCgeQSLj5
Y26k5n+MvRDH+VySNs3YS4vVKkB3VDAl/40bnoJFQC/h45rcFz40g/6EoSEnGRpjBuZGOm/BKylA
2zBBtJhaGFT2Y7RQOBT5jwl4IhqRqZ/etPG+0Z6yF4julhsX4EfKlbtngx4NDwGp7bpYI4IFnag0
kQfb9bbJuFOjjIuPYonrdp4Z10mtFa0XH8xU+0xJlALSesDb+cKz/7aH2AuO/Jf49K8FkfCDIQkb
jOHNXtORHamwxN/KMggNwkMquC1XQITgr7JhsSKBKMF4UMnKc81tpb9SAwLt4icJEPlZOe74gdIG
d+6MoHtG9VWTyhFc2A6M0lCsGSQWQCtXOch44/DmV1M4zkzeICPiKlOJOJ2yMCbww5ugAy57beTY
9UX9JAHaIk7Fm/BUYNcJnKm2KSRta5rJWtmkA3i5r9F5b1+xsD9ucD+auxOHh76N/6FJL8dig1Vr
w7GcccRzc6mXSUgggWNli2OUhoWvVndycmR5XPIkIwgyHEzKD90zlG2uSxug6HcxI6dNfezHjVgM
v0qtpVlMgu05Ar1UDMuRFGkpL85RJwFG2fBp0EoiqPTLswfKWTc4bIUXVGNbAnnfVcdpdfT/RZUl
yK5xj3sG5gGU3lhE5l5OaUQ3vj+WeH657mW5U36+zCSZt8PDh/OkoZfVse1udHfYZjEDO/mQs1K+
FPVhYgrnwV9BYfom1HcpCbURt/IIXwAPb3/gQIuamQeHJg0N+DZOD+Z7YujV7b0hmOmCS/W2wOGI
AF4EqAE2BsXJ1RKxiiHYaOEV9kT1hMSMonml+8vk4S5T1pZmOHrLr0nLXTgXkRkGfb6Q5+WV3001
mcs0dZ2+nSETs7jobHIS3ojw0WERVze1qEiYlfG01m9edgbARREm8+aQ/gCE75M6a1VtM05JGI++
dVoTFqBu14gg/hLHiRRb/vawxEVULFyPKAc4CxTi8UGcvatVpQpJ4nwDV8aKZ5FQ5SKMDsF5oLC6
oKty5kBm2Vns38EkwdA2g4dv6eMOlDyeIlj//npD0F+j8+Ex5jB3lkpucUazNFebvJwBDxcyAbcK
TlME1JO3LfQBQ97ulUIL+7V2wPrrM46xZXsdS0wDaPqZUhfgjvq6DQwr+/TYZs1xQ/uEtc1Ce8Hg
54wk+oLis/IeLXcDvXrahYOcO0enY2NKEV19gGMsf51DnxwrrU5UK8AYXkOI1vPX3A2p8hYUN22j
xytOGOzTHeVnw9Fwr3IQrh3fZLn6U1SuC283PkDtbm6FI0vCq6w9XLHtGgIK2VKl2mtK/qKH7f3i
cvGD9vsrm+GFsNNHzPnxFOrGAvq9cU/SZZj0diES/Ohpil4T8S7/DihJfx0xHMi2DHR8HkhjnUKf
nQhA8Haew+8g/PyTs0C0KkT/WqhGe1a1tyNAyyb2qsmd88HqUk+Tx45Bx7N8Xcdo/yeP1vd3/kbB
nAI3VfRC9KlL4SgdMVWPWqQR/KSm3Y/pt4qLuA69N22L8U9/sggff6MImGPyspatJZ/AOelfjpN+
krfXq2ikNqqido1ONj4bPukmvmFbo020Et/wyU4qS5ies1wEDh2+FLsuBgDymACZ3FNtb9ZRv7rk
Ic4XaKkLieH7hupPb7X5HgzSdYpwSpmDU8CqMb8lOwyxqHdwI0IuG6C06gVQFe5QJMRImBnmWE01
5NtyAEY0Nne7y09W+5ynGaRyckwW+RJy/clMQOOn4CxO6H5492u3DFSAyP+N4DN3O8ABku6+IVwQ
IPIOP09vSgMuO6Q24ezKCemdd47aOZ9EtZlhHIrBU5WjPhh8sQAEDR9OWkvBZCBAoI4HA19qtYO+
ccskjtPRlCK5iAty6M6slzudTtIMETxza/hPikiKweimF5AMLRHQwpyxivP1BZ4NJ8Cg3IUwvhjf
sYh9m/0pul+Idc+C/Pp4AmkS23lKQRASBjzBg5EXfvMaNcDH6t/fX/0ekYHVxqp7nC3wL80S788n
q/UHvMErMv4VO3Y4CBlAAZtperEq+OKlqY4Qx/ODi6u44GAdqbr1Hrqlk1F8NdzXP8ZuXqWJPesU
p1hS88WHqilli0x1/nLXy1j/xIGKBjEW3025x7piBeVBFSquG5dmqMs1raTaq4JZj/PVOgAXeUVG
6j+81RB80EYp36ZCXY0VFAC3PFZpFWWSu7w1+EdBXiQftiBrGceJH5Yp0Or3SObHf8RZC+B2WAht
W3Z1MN83jqC2uBuBWOJ+OBTBLolvTbYLQja5lLy6jJ0ZMjVEt7dYzXjpK3vfzjWiGrKkv7FWcBcb
4R3FVTNN9Y/5Xj744k95zhdcA46qxSuELqahKUVVG3QJHnOsrSajhJKLElolcDBeGh4X7NFJvNZv
Anafcc0jw5KQFaoa6Vw+E3YseeHbbYQF0vgLEhzbDKXo6EZMSKMfkwAOXaE+OSUGccpVJ28alq40
OhcrwObMrilJuqv3hBxHTTIS3Xv/rtB3zQjvS9fFpEs8SNDKtio/Cc/pDndCZGurk2HK0HeK2SUH
IOoJQu+UNXGRy+xAMytH/ckb47bHk4G4WLGLgsRCKC8xEAf3V8mixPOJDBAmxP88MRa7uJ7NdJS/
WIavtQyCuFfPrfK+iyM4muJFOSszpRrl5KNksGHhBqk3UpzlNCCYQY77FM2Idiwu9PKcEvhbN+oE
+lXeom1cd2YYybH/hoBHxFsccb90Mjox961uQf5ugebcZ0jHJXlD0dPJ4g8xic+zYYW1+V8x5hDD
EJM8dJ+EcGtpnM66smIB7Wrg6pPsjr0x7yeEcqU0ZbFC5L1Ei4DibACs59hQ3+Va9uypMBclUBMc
1bWWw0eypfOWJs8VgEX6/6a5MAvXDPmLiUPRcRSTY+YerxO7Z7yhaFGDKfkIAyLs8ojXK8lMU3wD
xOIUw3dzng0ch7xU+p9wREz28itNHnFaZFik3Ew7guON5+y9DoFUWingBQlBv05tiLgW72k+A1Eg
fg7Vfm5uC0Bi7+MqMhoj/Rv9kAKYpWFvaie4DE9gS83CNrv4ML2iBAJFyTL/x7GSsXY20DVMN26L
kgcyJJkFVff5+RqPns4/d6DsAHKwAeTTtLxgCM1axoC/qQzvqkjp2YrgyH4avgnr6vG4Uz458ygs
qAyQPNslBHyLCG/b0hFoTJ0U+KYdX09tWkjjygPCGaro3QBXogKMLWtvkwS7twYH2VwEj7d/8Ve3
k6+cOeINrgTM94x9XHh8xnqzLs1fsQS0pI5NQx9y+AeuOuKksvhZDm3/gHPFa9BTsin9sYgN3EEa
j/gWJfv23xviH0SqKjVmR2rjFWcbAXDtt8io7XEw6yDrdajXdrqf460Cew9h0pmbnO+H4sgIG64q
KVcCqPX4K49G7GSry/CD5zBAfhQ11ZUjglXmtdrTWCbfsAPgw+3kkIL9tW0QwcNfVhkoi+nlNR0W
h10TbsmEC72EArRLnV9DsTlHeneEu060p2BwA0NjeYvOhW3w7id1rVr8PBJwUjdshoE91MEYbwSg
owxTSMpQTp11m6R9zL3xy5O+s3tf9dm+e0sUzQzA1UdP7ASTYpL9YLMFmIUd/D+NzGQztHTjnmFl
6vwP94JXgGz+BVU3kM0WzM5Ge2+i8nu50mICmSMFcU/2jZUwWRmfzR90o9RFBfDG8wFTp63VjttS
WwqngqCPeRbAtlI8ugagYeRckSfrtN45Oa2nejVCBPwIsF6K9LJsptVKbMNNc8v7r+yHWSixYsz8
AnhAL39U5k3oAiAt3EsrJqBLSepLNbb/pLmoLsIRNjGm1GMZDR9fkHw2bYKF8r6WAoXh+o8rv/+n
ORKoGHEHxV/yCRYj1+pEImXdZE67b8Re0mU9DVxsmpLuHXTwgPanTvr9pyOdoZ2+SYoQSxRvUh/K
7G+giEoeZKsYn4FvDNLplCEJGtAOdYxU1wDhDzYI/n8Mq58v6vNWnmSMbDVI9uVzQsibhGVljFXL
+vPEuwpl96NeecvOi0Espqh+3fI5bkIPUy2qkbahHU9AB3EOK2AMYqxt4HNeuSBb0s25bBvqp1SO
pouYHBSu+/kh3a0jjIelbcqth1+g7wmeBltsOeSAApDkYKbRphgAXlqHUZLHSIGyKzJvgCdsiqLm
mTl5+cON/UvbWP27at+Nbqz/cmVtorP/EgtivrX8FriozhY6GLhw24j/7UEugXL2ishwvhzk3nXt
8DZH1CCQzHilOHGGaeTj57nSwIPvWjVJKiiYWJuafawuCNz572E29JBmG1SoC6sbPtd9JLR+XE3q
jbc6HoASXyB9VPwymzXjiNUfukknqkZ9CxV8CfRVRh+I/C4oBAQiyRQRTAILYmbTK7FWq9zsohkG
hE4fzkAwFfBtM8HgzQxy+Ar1VlLOrrePg8RAqOYU4fQ32rJyMHp/03ANLa+A9B2+2KxDHsIWYBVy
hnTVQ0x0QDTNMsS5bVb/gMxZs9PCESI959kq9ux7NtWNfWBhfae1okTjdjB6YbPr1lfyY87xoM8E
PnfEMT3YbJoXSY3mCyr4K11BMBzTLshIf+/MSrJCSbo7YTYR5eIn0DihKno3nV4rRist3sCm3wcz
R+JxFs7FlLrtQ6d5+JuVY14xlFJMV1VEy5DBOlIT7GURzB1xPV/uCG0QcoKJEZUMC0O43tRdjFsP
0ne2OuFRDUiB0d0Zeqx9bQzNANJlOpbL7j6O4K91cXvMxovT4exaHDVqbLlugkrLVONTwKYmoOW1
wSn+J5eVZY/5vKtPKrhlqfnJUYf8p9Bc8sC0vgF6JlcfiUmTMjtlu2KdoWbyInHo02OBLlN8F6GA
n3zWIAsgpqM8E0b/DlbHYhQzukVy/lDidCsCuHQX2nszcdqxQZ6tKMLjJVFz5wGOKTqG9Db8vUpY
aVyXc8ROeFYawGDypqFfpbMj2M3a6rjA05WSGryW9P+UEsfF+59MjNZUfXo9vsMeybP7WD2Jv1P6
SQBSpbKVu5dVG1xq4ocB40wS7amSHPSBx5t/f/EHulKnwiPqwr4dJV7mN1CgQTE2tBDydIBGxCV2
UsGxDqzuLJqEHRomXnma1SAdhdWytcMEKgRtCWB0cD6WwXT+9to4TQ0sWfw2Unc8IaySOE0KZQ+m
fbV36ceJxiQzwbGcnPl0gGNjnMvm4SgbEzA5AtJz6iA+Y/A+I7l5ogxoE9P6TAudo3UHEfAuVu2H
tb57iI/NguWxJU1v2Pr5q5FZeuu7WNhH1cYgosCv87m19AETIylKkIfwoYaoMd5RhqcXcSC9jQRc
qJn1wg2IWqH0y+9XO6tJIXNZc2iYthMzjnF9hM1fjLLtTmyNKogh7Wu3J/8XXo6SGtneMMjKnB61
C2zxBQzZpK22W3SNOkQtn6vhNQrZzdS2bPnSc6jE36u33eIs1OL0gZ+M9aHsvlNY4JJ+4SI4EfLZ
zQ5g5VOrWsJ2Df/YhqyR3RJf6YqTCYRrMAEOr+erN1g6oam5QaiWp73zknEFpDp0L+YCJqXNEQf4
d1fk5mpOJy2Qaz6RvHsDkiyTChTH601oQBzb7fVI/vrkXG7SWlfPiCP3Dd3B5iCgAxgeKlTy/p6h
6RN/IGX/NCI2PHnEP5WHz7SrvOSEd6UYuZEWOBWAmF0Jbj+13g4yKZ1a9L42IfEd4RHJt58JDE+D
MXorHBkFyBjd0YOlbrqO7a7nym6LGoMRkth1STv1fIjf2bKS4iAuXsuM8oWoHeqcSnlzOF3j3AUY
quWvkWYWpfMbIak/9frAaS7u8IJ/48uPCIgn9lOAX5W9qCD1ytqipJbBsZrsdTxs9MO2TbTSKsUl
ymA+25QqiAv217oEFQPXbeUa/fFrRQ3ZAz0POn42+D8TVvc4dR6nJ7nh8rRKY3saO3EGRQRcgoHh
RqI65Bd7LZI07wqjPLcWYrjV1nmiP2lHc7bCaPjksiavLzLi/xnZo1Q2Eli7iDttAxN/cYfduMYl
on+wLb8Osm6GyyWr1bFGHFKX2BQZbVxVO45VPo47/xFkTvidEkWYFQBHG6ORM1THFWjm3JtqEssI
R1MVKfkhCNTb/uVbZwURjft3TDjnRK56N/tYAeCxihYZsEmlGBcPDkKQRlV/DCv2nDvOKLoE20MV
BhaFthZ32/B7FMasbpTzze8x+TdVOVzcW3lMbsYFMla0eYajrvREtdMinGJMD7Ye/C/Iu6XI2ebW
Qew3WdaBw3+QkcEPLLNB1eZ8u8cN9EXu7jbbharFosVbY/IWvRXNiRDW+qxsRXjSPVCB9F/FGt3I
uTov4I4hW2D7FUtO8KWJCRmFWa7CV+NJLuLBIJQw4vRXxFL4J3/wEjKpVEMwAc8dpxGUblimGrck
q7krF+UHL8s9m/CQM5SiQNPWlz23IdSxHSCcx+BKUh0SSHuyMAt4LRcvP9XAKPL224vPDlvqudZu
c8JtXzj9fKUwn54hvJXpc3jK7lVEiIVAyXPIeOCKHCX4vXVbfFrx50ml5vxEH9dRtu2FFRNM6QHB
ceRPbYo42DR4vZX04h0azxGYWaXc8ZPG93RqOS7W7CVPTDoY7rYDu9lAH8tbn//ZmmW+g68D7Gjw
iOlus9eGYFiEIAN9tLAQhliaNP9iyQfdMA5Flnj3iNBTHn09aEyhB+us0KWddD5ScavQ4moIS/t8
PHh/jW3p6rbuk0dpzAfwlHVakUPlPxmwPrqvG/dgrihMQCfQO/sbYPQ6GniZ2cOZEBkK72jfTcDd
YbKMw+7E9qDD4R3gm75vZNRxXvnDWbV+5OrbvqOzMtM2tagx7GUCTpcAiqH5BqKWKuQfUprkHUi6
URQXaf+tDqyNN38xk5IbRH1o/O3Y/obzSrHfLnfkgaOLB0WxPFQX9rpZi+GyZUCbejLvCCi4gvND
KQ6KRddnYzYQs2b5E1V7jkvVnmmWhVAA4lO5uSSGTiKW2NAaEd607VlN+uYQyOutQQxWHPMC+1ZG
VtU4/6SsMGqLNMndJ5VTuug1JWVm2o2PVoDGKAroYz7kzZJ6pAhQVG8JDejetDb8eo/047VLlv1L
2Nmv20p89wFB+13aCgGWa1km+xCPmIOKB+pIbjiFIC81g0Ws4CatEKcyYXxmolEpowQuQJ02sNSH
0tu/nrrj+KrTUSM1g6P5VxGSjAC3WtlLMSvaoENnFcPZ6syCWbU8dmaFjHkgOP1/cq9/Qmy9e5O3
EQpGNBU1WWg6zTJhBAxUu56qijRCyMV0S0K/NVAYRRMYL81POOtHFraloqYC2BNYZ/TZEvQm5UuN
9N6V6hApNc4xPpD937LjQEd6gzz/0cszmspkNNxIMjgTddrCmwSRckGFlLdjwltOfczqNKgizlnP
WN247Q58ZBxIa2OKJvq4dj7vcmvYcQi4c6w1IaAyzGiHb/pvqJFq7QsYNeDrTnb8lWkDDbWBNGeG
XIdG3xXoHrThQ7UMWNKe47MXZWjahcBbSMoI6AneR7p8/dMt/Qm7HFENaLCz1s3FWNWYz9ihPz6d
oyNL03qBW8p3ofWBGkJSoWqTbJB3TODIKStJpYA838UsDDuiKC+nQDgZtJpNusJY6J+6UPFa14du
bmf/qeCS+ER01VdvKKjyZV1WwPzZ/d7OSVPWeq1SCxOC3oLMs3z4Eo/eZ/e5r3kedB3uRpj6eI1H
xt4jcZ/ZDLpEAayJTRq2V8MVmVH9Ot3LVrAhqhRr9TAm9BvqKbqitq5Na4OIB7dXo90QZSnIJsRn
t6K0aaz7ss4cqB4XyyVn5AI/T8CTyqXhQrW0KBY+KoCie0ouPQVnIQLg7kQFlBuuXnjvPWmGzMcb
EUqkGYQx/mviT3HBRMhJN5hyGGVIsiPjlhXsKbJ3qPv90wyA/o+Obq6hNMk510jZUt9UR6KcpcSB
Znx3cCk8D8cW3XBa8z7G2hBEWp14OP8KvREEuzXdTRNdYXSdD+BQx1fu8WsbFLqDYYQii8IIR0wR
OZLdqT1lvTqvsOE3hIDIed6KDsxrw/zCCNhxa3Sbibdv7+lYIlRW1ljWUHoKTlMMVxRsPG7lnKZG
SYSKbP2xu+JO2Um/AVTZS5Ej/CTOKWkhbUl0C6woEIEzddp/HqV6+e6JgLOefDQu2nTZcwyg8+aH
DTREVQIeVS0eeCsRQOHYik/BV6mBvhwscodjJaF7vfBC2EchseHX9b1Ms7kYNNOndBFqxB+0LSt0
f6wrUwovRF2CzS6MbZxLampFIZdAB260CeZhpL4NnpelQrcmrZeKxpXfdNQofWZkQduI02TcwK0z
eyxNry+8xYU3JWVW9sHZj06CvN+nkn7Ugsln2acMkdzSaB8+zuAuj0VHskxKAmdm0hmBInsLAI6L
TtXWZtyFZhCT7xPgCoQ0tWz0eGwBrJY1A5JdsNsi5ej7QZfzWqW5lXUx9CHKtSPJfV28vA7KGHid
hzyxkgQHNRGfiWoJCmXRrDl+k5YPTBOsMVTskDuvGyUzM2De8OQqUAy+dANWux4ovsx4gkNOUNmr
Oy+2szHYweQVrmh9yjQ0ojECIAJ9vRNkZS/fcqC5xDYlGrAdXBBxeRKL74EisOYKc3RSY4SPZES0
BiDpwEFgYK1sxFqQI6R+94vRF52W9VAGej/qrY5m9EB/tdJ1nE9afC8dMmItscLEB7hXPFvdMw0I
ILJ40EX2w4kGDiotahml8+bsvIbf40hKwa8dFKQzbyPSoGcAK4j0t5mfgEzB6XdxuZPTFVtE/fDy
DchvYN+NDkbwrJ0Ka3nfkdI2ETpMfy3OTYhnGV1nhkNFG42YV3/P0ewXQ++1Rhwp/y6sl5BdOprm
qSgWOIAxfZfPrBHuL0jTwCZK5YcZ3sGScA68idnZJ9WSDWVlDhQ00ilstlQlnLsBLs10fTCC6WVh
zliEb1fx2jMTLH89mMh0cZT9tccCy1lIsTVHbJ6G0I78xs8NnqsC8EzjfQkJp7NMezqar3K6amQa
px9GE50+Voy7Oxqf5KOG4kfdVjtnUjb8WB8TWVnn1yjDIUvtjPZsXXXT/hJ99cwCWomQwqqlbDW2
gZ/ujql9NZ+fT/zrrPNeydfNrRiDXIjAUdFvKNHeJ7gCrV2mmWBtyEPdMMuBvSCQQ7g92ougbgdW
3MS6dlNXDuuGzyIQbmpRfVHFt1Et8PUHgtxdGE9o7czp9By2Pctm8mjuP7qq30REhm+MHGZtEp7y
7n8VJ65PS3z/B/xZIEZjn1Ew//MSUhDR4X9W2H/FPZ09fV62QfTECnDwz4+3D1Hu2a5EvAmN101b
T5/5HgovumVTTL2YBkiWxW3UuUTI4InZZzHzt+XI2yrHcNkSDmbUMxFk96mYzsW88GkA5s3xyYke
+s3RBg3RgUA2usUq4jg2vJSG8PTF5KoyUJP2JokQjMyFSGAkRqgw2V78se0Kkep0pYD4g2T0vWbO
KQM/lehL6KkE7D0ANf31ICqbybJ/X6MzDMpczCyFOg2P8JsggJ8s0OH0s9M6MnAZsLrTIEppEvTZ
wH21X2tf7eIORUezfsh9/PbhKX6omVtfkCN2Kg8mm5N1J8ThuqzRY522vybl/CuW+f8EE1PkgwVJ
ysTnhVBk19c1yIozycucJ2EpYISZ1OkCFyW5UO3EI33v4bxRSGqiERVYALWCr0j6YAqxber+1xYr
iY2R7XUYlvklThd94Nmeii+gyip6Wkx2YCSYBpxsJc2xYNLkdc5FtaQ1tFis1r6y8Qmj631Z1blL
dhJzm8yeCxLB7Vnhm98cu9Zhjvzt1QleTn9pbNFtyUf9+eGztFWhecAM8vre40EoAcg+R8i0yIm3
pBXbzdlZjxDdUlmGDo9OBGF6bhhavE2e8T7cyqvGqEF/ldZXlqcchq62j6uItxSDG3ATyTZLjOjt
pTGM9nkJSOq5zrqXlJJkT+uemgPTBr1F0VjvI4aCLizJ70oCeJVhF7AisyJowWV68kjL81Yw5OzN
/QDvJSVeKapAF9EHjiFf+dKx1Hv5caCW7SrGv9Q/DNFS1JNr+FMeedZM04TZiXXXYd2s+IYMWL5X
8oGtvzRiTwp1RPja1TUYc9+zBWlHUSUsHpc0hx17P7xRVM6xSdMgBOX15y3ixkgxDyMWJdVJk4NF
OpaBBsO8bhmEcdPlfPR5oS4JVnCKDqTSC4hrMei1supZEvj8JxeGgxA5zZAdNuWhAIoQm3Hf8eKb
OVS6cZsi98SkrcBDEyiyiYBpxZCo21OFknJ+qyKH167QQ91j/mqq3LypKDBH+5rZLL6Dd1H7I+Qu
P2HG+c3+OpuaJUOvhv5ueid1/h7GnN5rCalelsDs7Vjy/DK9n81yxNuNfEP8Kf1VOGH+b6RGllU7
KWcPd6Mrub+3pgt9fgplBZPCbwOXTBzdudtuy2B+eHM2jrZPFuPj0BEtL1qT1YPqkiiKuGbnpWc5
XeVP3rSGT8MT0/bJBp85vBqqVGCtlNoMugC3BZU5sA8Sj7f3btwFrdYUYzdCFlqZFy/CRIJXGQwh
mRm2vuJ8sD9erPOJB2RkRd1PFsM93Hb0O9cWT6JOfWGA7unYcu27sSdBLMja2UpbPQpPxDYGXAlu
KL5a2Y4LgvXKFy5UKjwkXuidFl7Oe3UkI12dVjyrW/u605LD7e93dPfgyEqhU0mRC17X2KXvOFMi
t0+P8bdiACSrcnLdh/c84Qwm8IWp2TAN6ZVF+Mko/BVOewM//l6LlAXP6r7k2YaM2YQ4DzXbajBD
A69oYvPqmPyeP1ExPM56nwqdcd0e2Hz2AtfJzZq+QTP131oQn+lq0dzLHup+PepEadfulQChK6eY
xg1772kp1cng1+npusnpNRoy6k5Ja07tLVMYlCbsgRekcBE/O8ZvkmpCPxHzS0ZgNHGys8jkn6zX
W3F4j4QLTsVjsmT1cE1z1X5bsdls2sOqSbemdwPDx90L+OPrK0ogxN4/qerktAHlpx/Hh4UkfezT
Bo1xpza+ElJJLRcGbb/fBtn1noY34hNVhqD2k9hFIfSi8xSQG7pKWYRHFgx6CQ7KXFT2MK2bB5IS
fvSZ7PEa236lSQIXFUYmzXR2jIK7nyBv9kskYt4+IXTlPaVJPrHQzQxgH4lB/Svh++AYiV2peFLv
pRiX/3kzVW6c4WOG820VP/DVmBbNbY42AA3jE61HVrdwdnKUDyzBKejATBLhg+zWWHwIwlmzGZyP
nkRcZPH3TvZO0NigB564MtIuMeUJVvRawnErfBqYagkLpMe66Zh4TfbuZ+agZfehrknqAWq1Gp+c
JEYqokM4quko+lrE6U5jGN1urySziPOnMXC9cH2tXwBduqJKd5rc3q1aZUsV/vaekb46u3v9laML
WL6NDZd1i86O95PQaYATjCdpTo917r2qtZvN7Ddm3XPUHEyfx6z8weoRRUrfCQv3Q9O586iZ3gyM
Fm33yzjeG92/gZX0B9M/pqL+GvzHuUoX9G3OW/6X5k3yqqXJ+OpXXvGhZm+xEHb2EJOwBs/X98rg
LrPqKTUpm0hyWpP9hs1X7B9VCMYQC7IbunARZYSlASASyhcU7YdBszhCdn/FcXAUtVprJaPnNF9l
FRkPWk3IJ04kuE//yi9KJqKYAOXHyDrlZWExziXbD2+RUBCdkTkjHxj/qMb4aNg3kjI4CrTfvXMg
fh6uU2gg9B//T8JgcO6Rk1o6TL53N0isk5TjBNvuMO1zNcZTP7SNpy+Pbyfb4i3fGHc7G/Z0Hc2S
sN2/uLam82O+eQYrN7CAWrV9vucaJo3Ngnzl3V+fYmgmVHj9K8g+N78xsE1hxT6qy0FjiB+Djmag
+lPaWzVnLrlzxDqKYiimXyHql17zWRg0A/lOsLxrUmi4h8gEsOZwBRdSEvEh9DMUPFPmhjjOvPGf
HMmiPt2RhLTZqL+bJjGWhVln7ji/qiHunwG9ovYccHRS1jO62uCKMbj4UgqUKroL/P8u1qrw5G9l
uG2sQ9nHySdytSCuhAUArmRyZtWYTVn1jZteTr4A5VJbULlpMh6a80VgWxN7GcM+E/eAJtmI4L64
Sfd7Gu/ji68z6EjuoL0JlPgGynmPv562pnwzAQV/82smyKzSHooccqEiGpzA0oKCZu32N0d2W3UY
WLvLAYPndoE4b+en5wf9dkUTvMd/+InqCZqo0ACNAr4b7g+IKHK8kwKgzWrpZ9L/YV4qx/qlptVT
opkLR43+cMWyQnIytOWodDYsPAfV54qPXHEPRWAAkuKAtm2AFVARpngTCOOBEwzl+dsI8zM6R89b
z1z4kWmC9fryUmEFhZvDtlTh7Dr8lpPVoCPrkAjm1aG1R3RcLCtJsvnjsMEjvNRrZNAEKu28qUz/
MoMSFuYhOCyiRHJSYkmRMuPbh7Z/Drd3aavrfZpQZjrRBklIYYwTFSQVC/5muN4O8uQbqAAnLMoy
gIbRHxQ/8YniK2c9kG5vXP939TH8qO4dXP4SU8bCnMfFVXWSqXtktBFrfwjRsm+20P8kjxPOTTeV
9AZ430e+cQirWATTvlGfeIpJBlr6n3BZQLYi3TwN2s3tjFfUSOZEkuUB7DG0T3V0sGnXptBlzuG1
avOeyk6GedJGJtNmFrIwylJdNL31aN8i+GtNEsg/Phz4eXidV1JSHUJdhtK58xgFZrvlDZHFHOM7
zNGdjkPvlnLvb+EIN1XxIIbvIWXVgjD7MJHmLVC21GeLDBu/xes+ciqo4F+oC4UJ1DQdZwQnugzI
tOS25z7ASt76Sfx+7JwLx3g+3363+vZO0QLCZd2/yjhYv+2F3SzDmdhNMfz1+K/12CMGZdM2kzvi
gE3vyM4yD2O+dNmSBWjSaSWzESTbh5/BgLGwXvX03dEwjG6wdNoaxtmgEYF7wDNM7+ibKW0HLh9s
UezFDbmnNJ8AeLB18X+iuyyXNni+aZolqkG+z2QRw7nbIAS/2Q9IVkz3aGFbYMtymkujDPYDUAnO
gLLuN0kX1niPgL6XgnHPCOqOtEQGX9rWDHI9+slVZNPcRs1mCdqiRTfo3Ud7NMzLqelqdkHyWuG1
7ACml6rVUa0/DbvnyI4AwVVkAolHoetLhE4FSqZ1l6XlCFODvIWIppkqwWwFCw9QqeYzif9M4pdq
7rS4v/id3K0epC9ORF5OiYNSt1WJI6OdTDxjKPzJWTM36g4m0bVfluzzFcE/5APYm/TlsYHOd6MI
3JE4xP++t1UgYabWXTXCizRIXCju3viin7cNeWF7PDmDMDVucwPCQ9MUPOt0kvw1fGIgmtSFNUfu
dMhnVO4bKSq7rQLzi5d/jJDbGUmI7qkwiSPiRXQ6ZfjzAsEEcr/VWVZ0ExmAqJZwgDG43iDXinsK
N3U6xzY1oM7I8dEpO5Cw9abYr2rgTW8YVbNoq4OmIboi6vBwgF0qfGr0BfG/aU8LR9fmrcNu25ZQ
+RN/5DEWYJ1h0DWc1wmoUTAnGH0jDgJ0K827fBWsZ7qiPohDQmk6op+yXkMuWTGaRei4HN0caHhe
tdZjX7rjkenG4cV43a7DSaQ29zvRnD9CvJpSn2KCDLKtfvhXZGG9YDtFAbbE4vCv5/2o28Ialt6Y
hisnmGeX2kYCda+GIS6E6yIi7ocy9bijHLXtdkxmXyBSbG6sBoqhDEGVeZmQWoD643VaLA6HUh06
FY9jLD5+HGAo4wbk0yairBSK90FuhtwEsiAa17SpgQFljUfpvMmA0c7hqFFcbgTG4lsvj2MZmZPO
9pAM9j9o+bm7sfu7fmviY2YNe6ChqjU/cFsstQYTQg3uAunYXFNX+tVtnEpCCCmQljXoeYnrhM6+
BYQiz+sS0msRt+eEz1mC7QRSM64/DjA6QP8fwUh8ilB5vUUeIfuqON3jrciErOS/ekRh3bEZIKkA
HbcglKaO2z0GcvkSVxJ7lt8kV+XgvdT5Ch0qcrBEvjorkistyvdmCMJG2Y4zzeec5hp+zjdrutRV
BHRLls+oQc31hhh60N+aDqxFnbsJ7F1LtAQqRnMF5jEOg7BHzMayLDJ1Dr/TrtdKs/GDZG1oRzjE
70791hZB0/fHho+SvBTsP+E7Cvo6RrWoqcuHf+wNcEf8jyPer3j5xXVNAbamDWeXJatj4GkyXJNO
gVsDvlX+Qn+IgBV18b0OGL4S7TU980NykHnUwPUkfiQvgmbzUpFHsZrRapwMIOZORqGeP3qq4pU8
1tWm8OGjarCZQkzGwWOZ3ZXKrEPYDd09xQndOqaHhXa6YQ2UaNI5CfKmYb6YHPhYjWIwmOyskJt5
nfLJK/iCTk70yQG1gH1Jap/boCgPbbPNbhGOR5hXcgmd6ngYwzsBH69XsgFcAimrU784N9GlZ+oX
I/e20ay4uszYJbe1LHwvQZbdFb914Q6KpTNyVcdsW0ZTpja/0mixQs4B9KnIqpGSJPZEwt8/KXij
XNEr3kQtvnJHwzAGXRVoB59eMeb3hUdu3FmdDphg7Q1YOZKZpLY7ZO/JnC4TlBA+pUBUyngUd/xG
biVan3X7bSIIDvU5BQ8e/wMqdpQV8+pmkNk0TQNE2w8XhbIyNi711Xb6U+4R6JNSRP+O4mXqAXC6
UuvTJ6DTedwJsF1rZQj9PDnKeCjlIT9CLQKT1194/rVXRCXVEgpgNCoDEjryVUZWbhGIKNa17WNA
VnfT2PIRbkC5ry6I4U3jKy4GYsdWhnx+HlqgDAej7lVTJXZN4e588WAanxAFlRUhYgKlWB0dL1DV
XLXmczwbqWYxpE+RoTe7EG5qvVztnZf+OLbvh0Hbz62WeLv/zz4aoRjpFGam6Ciyzf8t0N8z29dn
Jz5dZ5YQ67pQxUgmb9ggfHMdgJ+MNKufE5mHcZm1qXjGNgJPnlJ3zbmspF623fCoXdO/CaFl3xNY
ARFiDAxkBIy9nJ6pjEHD8n1sWsEFbx463g24+mnj7GhxU2SKg8OWrmcF9MrIGSNxA7BcWS6tLSYf
sGkh73Kj2fKY2YW4uAtttJNhK1z6Utt4rm6sbuvxroZf39PwkBT/M94m73qZz5R5YZCYjghMKPN6
Fk+exudXEcovurm1ebn1FnmfKDIQIOv0J6sdp+dnHK7veAnJCAbTLk15ZRkJFJv0cUZiglnhN9bo
qU6ORTbaU6vfWWXtSJsLNoo6Hwpq689xU0iE3f8+KC80fHZM7vst08V441RDTRsVO8t7tdi5JRcb
TkDwVqs0iaTkIQzqijnuY2tgjaYTxFpUBUahaB6L6Vg0BzZy1knKQ64LzCOvsICxmhgT+bISJNUV
vvXRvNTYv6Zoi7CL5lo2v19WBBwcKaTbeKGDbuqqeNC4bYJwdFRt7W1F6CevnIKTh5KVhzwsnY1o
fnHTTzmlPQ5fblywKIQqPBdD1A340r3OdYygoMPEhc3lY/uCXJpT3MSHaxuPTtEcEn2Ae2ieUeUQ
Dj5dGi16p/gzMWoVg9lQNCp62traOhqrsIiePIKX2b5i+DhN0igAzWHEOxz67KIEJm3rMHTZ/5Nh
p1eHrtlDgjChYjU+GSoT8eH7l8EYaBExagGmd+G9ocyx1Dkvvz8wwfMfp5kbd0NVSoGQkWoipY4I
ERgraxGYzFpzyaYYv/or5tmXyAGjrTthv+eECJLEEiHQ7H9djv6oEvgn4bwLH6sD/6aGKzIkeoIZ
TU8wqPZJhSaRVmh3kHPlIcLcqiKOMx8S+jm0tVUf5G4q0dnvzLaj/nJHn46LoaeNAJ81S6XW/oLn
rAj3El/qdYMNtzHkgGn75WHdhDXuwnX+/sdDuwJt4gK5gpF7Wiiu7m9pTj/dTCQYRqTc3M5yau/F
06hWaY0ZgSO0jNfTxuS5Y/v9GcR3nmWRuzIRjuPtP4YHIE6EzAfYvwqUuG871zm+qpSE9C9//yhL
7MC+DT6l3aBpxJYEWSDfgueA5Hjb3zbNHuda2IqAmhLsqIGEPj5GXj+g93cdPFo+1xLABfDj/baU
pQOCELf3xwPGhREMKqkXWdVZAbkQ/Z0LUX5uNLve7wO4gkIg4YcdQ2vMg4eoTrcUP0mPcUQvYnH8
MxszA1iN6Orr1R0O1jP8M8eXR/8FhFSZP09ntNHAcTfTQSksvyDRmlUg1YgU0T8QPPN2mJ1dVWBh
kahP0jcp+vY8JVei4D69nGmWzSYJH7DV91DzRyk7ft0iZt0jD3vi3/JX75WnFb1IwC1BP7ZdcN1k
YzLVxNxjY2gLW5qPoDRlehuEMu0dJd9Pwiz9GqYaALyBcSfP4vZvn7sY4wSNzfBHTVJ7cx+c2gqh
s+iPa6pGjbR2alAZRmdfygauxt0J4Edl9JPWcwrPSZtn6HUbUQ6rs4HsdbZgPR4qOY6QL9aCm86/
J5DGYqNQYk/vFSK3k9sFUp533TgD5zdB+LwFNYMNw8ydfOIdzaLLQjYNRSxdS/TFMV+tnXFxHcPc
DSDTZ9wImPTHZ7vdIjdgPVYyqbx5QcB78EY+kW+c81iEOJXNzjcATflpfRzYlV+fUUN1YBgKzcAL
1TPqxLJUgSofgoF2f4HA7k8A+h17R0g7AvQBqq/wXrUYAl12hP98J10MOIrZF0atKBO14dSbf8Ew
l+pP9BbJRkX955gCw+QgzHPx0Ow2h5sxfozdOCFLDt23XFK842GfgJS9YaBmwN9yjxofZ8nHYnYp
EBAgaJLwU3Q4XohgkvbQFwudalxWkhSUoA0dL0fs1WC7Wp50QW0ePNSWp+xnZT6EPladxrkPrx0A
PXZieQWK5dScHSoqTXUFJKL3e8Czj7Jr2bk0a8Kj3Eu+b9lIso5E/wArBBpBfn/S7DD6ncxUbi/o
OEAGuJPsgg6sda2HPD3fKU8AIhrZH9CpmlkQYCV6d0zgYeYYaORAyAMMeY6xYSnnRuiaAljKhUbk
NtJPdeeTVApIqD9ZuyeWAClc+/BjJDDPO9EJpeAL0/T0tgrN4LU6DeSJc3XcHFVj3LZKt8twXiSn
t0kQEftGXm31g4S8gfKlEu8vxCR1gN2z4VLI4W2xHabMBtjiN5C063V1vZ9v2hoATs2sv/zZnwJN
aQINETEhnNhI/F48PDvvtG8EDAyx86sNSyolxNeqx1wW3+Fa9aQumZZtwa8hT3qX65jhCfWHWOYM
UKp+KqeCNHAnu3HjxnVAtUv9FwigHInafzg7pwyxTCWh9+c1R6FOi4lvZD4KdnfQliNuyng7ZusG
SzmsHo1Yp0TCxqSGJcfW0fovNGjZXGg64rMOAWmCrpdkhy8otjew63Z7yLAmQDYLhr7rfLR/nhs1
i1FG9RQb76dxxvnr2pzwevNyoT3M2s9QBcQPqffQ/k4/BRBD4fFNEgFOHRO+OqJY40MDLb7zm0aQ
GGmO6VXeTtNxSN/hhZtpvaZYjI4LTOXcz/yW07ftYmQeGI12DlLVoOxJO97OY3gmin1C5XCzi3aG
Q3ZMplGTCVWPKjahnfSWBxeoQHRNbKRXdHhG/w+biMEMWANlC25YShcMS2RLHwN8p58UrFctESgn
TnoU5KMF1hgh2OcvfcUPwMQJ3mqBpbg6RONKRXExud4d/Br/WVgvrC/vmIsP1gCaZeuDWZYkFeY3
SkPJri5a6VdeytBlUaK6Z4Ht56fu8yzOlUweRzeUxgQ+UUjTxsBjozpK7IYyFkjC9dRQK9dtUle/
y3pddY5o8Mlr/Q62Y8Kd/NaNYdNj11LAK7wur1MaygTN3RIu7nW6NXSvfMX+0r34nfwL5+V/uAWi
zfhlgu8gdQN+ZrNB26kVvjhaq/uJyGnsiJ7Qzco2q4XLJi/oMANLTi0i0B4wXPryvZzkWN6HGnxC
KwoC9Lwg3zBT6O5czV+aIbhL4DNP2JUwsq0DHScJTNaK/XDZSnDhEw3YvK63tCcFV2OjO3EZ0dsO
GaTip/BROiJaMFOAX0kqtDHQgy2t6TlY/cDH03bqq3iQw0H0aVklnoBNECt5/PcRExMqj9TuOiPT
Q1DZDFdJz0cc+2pMrE75b6sq5nkJ2V9ZCpksv8COerGiJWlWdZ524lBoxGe3FvaD65aUfwTHn8J0
91a7dXKgj6+348vRmP54MN85zH0WQA7eFYrHOmA14Wmse5kh0x2AnzCvNPNAP1BTcNLg+YW+yWOC
LesJoIZb9AFc4nLsHPBUqW8muQZR0cT4l/oVJlyblB7jhZmCOAByKgubWPalZeYph8TEpKkmnszV
m/GOo3KeW9Ply3c67vfFTlvlBeAEJEmH0Te5WbJmFp5P3ubUjT/v/Nx0JbTHkNTuovXsGyt9UTyz
Ns0bJKfYtQSnm2P5niIThyu3/QLNJSUJD2k/grZOtqjm2kcDvUZUVA7aBys4fgbafTmryZIO/acf
2KZ9H/9b9V8WDA0Tqh+pP5L3dj5kIiUb8See2faawEHv5w+Se7cDzAcczqW6sT97vH/PJeRNhmne
cdjBD4zh+SH1bbHkEt2T96EAV/OvMWT5GX9ujZtSVn1aPTNmUaa/AhnhJ+JAt3wchNjeP7hq/TFZ
IfQFIHJ6qyW/icjGdY2nnmnuthwVi2hBCfc2Fca6eQm2pjwqs5/eiAFWKITPsmLBTdAK1BxbCVWx
Uh1rLBdNZYLaeICJ0SFFkHbjQfWWX5LH4jM8g88cMKpDeq+MvyMtzKCPrtLycdiM9ZzFh4/jJMYb
3Ig7h5DJILs4woZNlsryGkVtTdDbsgC32FjpK1Y/qzyBpuv3D+x1s/WpzMEEzUVPKEcDZmM2BBIa
Qmq9f36wu5JPcudOE52CFtDBBhgrXrGp3RuSoSJTkFqzF/ydJV1uXX/yQbRVhVrVjeVLx/j7ByBh
COQ175hjt09v+ETNt+XvCqk2vTstBbX8FFO2skSPwqx88FYZBZxZtv6iC77wf6SKw+17cRrx0TYi
3W7BX/YP+84b4nnX3wsNqUODMNTpdkP/8UThBmV8bZvjHiPjWV7qemc5Od481ynzIrDcW2az2W3q
DECnVcv/aTnOds8DWvdAVp0Trkp03r3L9VSeLxgnljz77J5vi4+YwREWzPq8M/TTn/xJ4JLQpQyi
brd9EDBd6OPD+CHMEAvQlap2NNEn3Mf6FPiDJR/kjB3Di+QrAvsL6+u5KFKtwrG6eF2DBS1Kczbn
OUlAkL/kcdchtGwZQfyIO2TlWMCN/3hgWzE5wfBPmfLKMkJunJrLl2dZhwasQTS60/Jf+5d3dSiF
GllBCIY0Atiy32n2ZzhkAnhUVugFuhu1F+bd6NOEpG/SsVOkXptS0rDrkxINEsVEKPiAQGri0Yv/
NXxUXRbdY77LcMeZmPeRAVNNul4CDZqRtSIzQCPLHXUHbmMTD4wJNUkqkA25qJE/z3EaVVxJkHYt
pJKr4klQ63Smfu8pIHxUMQpZscF//CMfr5XO4/K1Ld0e9aTCndB515MxaBU0S7mxPQlwIj+eGX8w
ps7z4vnCdwVCQjniL27fl+z/65oiQBW1HQaRqP4cS0Ig+xz1FntZsYpAIWIQB+Hif6nfd3Rn50pd
zkWvPjkBWZ16TcUjZVWYbz4RQIpKZN3ezTtX96nzPGAaBmmPbrGLMa98eBZCSNlYfaTozbvBtXw5
KCLl8s8SZND8v9p2UroK7x3bmkCI/RecGBjJlJ89kBZO2szVplwTTXqOqyjEvtSejgdQUdAy18Dg
UZj5zHomMkKemJ8vVjkCXe69aWabHVoyfQVuchJ0CfMaDWb6ZHvBrFRtEvQDgbW8OreME7lszgRQ
PTJXWcuInvdJF+i9LdHtbEmyWilTID7A4fQgs3NJgpKw2IYovVCe5b3b1ZKUhshyhNW62zNXvHBI
F6Us7dU0FIYzM73ElkVoePpttpKSfnPJdPjQYdaoTQctw/hBMdzs/B3Q95TFqzTup7QTKJ6Umx0d
45MuYPKutPqjsJV9mRPzUzyspwc0tRK7AajouI3wCUIbW8lgtjCbfY2bjVfxu0RcosPQdLn0tau5
UoXFDge6PZ8syp9xbCUVHc41GJywpwnDO9giqQY259q0k6wilP8wO2y4+Y5DbxKV7uYs6NxKPOTb
8v4RvdlXGhXFWNVgF+fpXxrJ/Bl/UvlyUMQxa7m21Ad1+tkII9Rk8OGTafq1a+SmYS/DdsRgKKNL
hIORH9JWwKU+aMxBrK3bW5wYY/2rjFkrI5dX3nlNUJKbRqwmLy5KLQswxSWCFttAmxkSRTTWg9An
JePjVXY9ulqG/7SSeyQQr623vcZdPT1SnMfOmVEnK94v4ZH+u9RoKupJGOVsJBQgDg04UDzxdWQx
9P0QnyXvMkA9dBapoeWm1oPNWzzwLwzeY5Ow2Oa3A7+j8lpqQ0CPWor5SRf+M6vUIN6LpG4Txl+o
qRPRqaBjVBqd9DwxOeNII1rsScE1FNyDfPBQEaej9cgoF4vgvtuuNLpGfZj9LwYwWLJ3VbNyCjMs
1ElOiw8OsukoYfGAmAi2seIf8IA0f5OsLQRZKNSx8H+UJDGZDEgXAoaGC7wPSHlpeLd5yk2nN4lc
tdY34fPiwCBMmYDyaPxO8xbpqGAWQk8HU4BnrtI4/U476yUCPrETi32Qb86Aqqmn+o2Q/XhZoUvw
mkpdbBLcDOiWDlTlWQ7sghl1BPiBqx0tXY8ZV5jCCgvsvgxvUzpRXuPCDCSdPWeNB5OPLLbpOiRB
aaNCDwc6lj2peqAAnFWkxQ/Y82AAL8K9l39zXhLvzDTjsnDfkzyR64I56se9oFu1K593STcjxacE
atvwttdP2zibmo5cB9Nm9kDXiQdGMpzp5Yt9acXHP+EDYtKvh7MnjikZJx24E0Sxh3VaL/dq8g5O
YODr+gZccpvJv8+46z2pEyw5uWqn3guZ5NV5nQJuqmFRjCvIWBzEncpWBUcr2CxVtV7wITfkSzqU
nhcyUnKdimmT5wf1M2s1SWXfiaLzQoyPhAMoWHk/Eqaw9kDajR5nGnoC887omoVCVvxdfpZn9WDm
NyDCnBqE7MnuFDvIMKym3pZ5BGlAd4Xwcl4PfN39rcFzuR/4qiP0LH64zB3VGTb9Ky25YJRsV38A
Gc0TBPrKwKgFERaeERn2fB2FKQpwaKrWTTK+Noo35432kNVsmEJ5Ph9a1KHb46aKWDBMTfF8hYLz
y7As64KBwZMN3UOCdUFNEblzTr1rJpDMPmUHLjBF+2Xikp7xaL5DA2qpJyu+LaguO/h0345ieyJ8
z3OvTPvUpq+wdzLmUqmnHdOoNTlKgPhuitepSS98ISd5OHxctajNWjBoKQ1CoDDPZEqhVGQnI0GE
k4721SXVasynwPnzLZZXRTJxyD9dsUneK13df2Sj3ocwxkRTtRSNvq+HZ1VytbHKtsalMr5f4u29
WhY5n8RdImZp6agdqVO2As/LqdBa8K3p31yhSNGxqaRIpyPKniu24S3FRRXdtN4kFBlgbl5HTvS1
PmxhmzLzXpHHxQ4O7UUgfPUDRXTed85A3CaiWvdef/FdfCgCbAMMIcXkec46+P8ZgXDxyJb5X9vO
U0MChLdIihQ6p721xY+pCW41iUnJlhDQ1BflItW/erPD1MBebSfsLG2+vh1ain9pcKGd9UBJ5GKS
/2k5j+BVGGwuiq31IW8/o+bMGwyVY90tq/r7RYPXqFSlvWF3Atm573D423ldn2C4rB+eU14yDTDZ
2J/QmuieLswfCeL/kzMYvBlCg6vkvSPpjocO4+kflK+AOAtX1czSaPyzxu2apCiHJ+yA1ni7x47a
nPfyQo0g+/pf4TALqedOa7kLva0kkBAxQbqAUaW3bGUxs/HMUUkGFLqaI0aUk/ai1ztpk2Vy9F8D
h9O8r1xFN8heDDNzr+u7BtOUGNaVRD2iUmLJYf6c4To1qH972hkfwuNhYmL8J5QoS6GAsWWyHfD5
yheIcDLUC6O1Ul/2SQVkZNgC/DxAXV3odvs9qgEJHpHwtMB2kzvVf9/DLoh92rYnruBY+GL5z+TL
mXIQyHi9SbVrW66Y/ky68YA8hO6FggTaqw7PoGVpCPXq9iZmHJLtimEVrFYP3X2Ia0XIdqoTaj/z
VzsVQwuB0FZIdFGB9fV8KckDUEyb9EGPq37GrSnwybXLHi+be6UTuRclMpIVWHCH7i0G7gYm01In
gapadvI8SyTgcEsTO0BxLL25TLZP+Pudrw8R6fBoUI/LkE8ZM6n9+jNzW1bDUmD9urPHqhAdW9sY
o1mrO9C5Wo/w4lqlZ67l7uzHS1/Uy/NzApXubWjAVmNzc1Bfu53JFXJaAgKhIpFV/LE/pnYgezYd
vE7zyMlpJUEr2BhAssrFgQT96IDLoQHiaN0VyMYQm7e0F53Wrmp36vQvdGOTcDcJtuNZSVR/tUNu
UC5kkF08ILOv3vLzioca9xIeZZ9aAmqiWveYHTtd6hP495fsRHC3Fcglkm45MaOF25dmltNcmYxJ
sUNdThmfroLHolLHMpaSbGKJg45xTHDrdxcYZgSOELDPR/lP9GazcA88d33xzynnxJKCrRY8LHnF
mJtTeONClwqgqco65/N4DXe8t8sJTzNT3m0wVt+OIBFV8nMK+v9MRrfuLM0tUrGQx4bD9zFMSqOd
B42Y6eJoWJD+P4XQH94P58+nZ9pEoabdmH+MW3YPyghstLmpaF2VYV1NjO445OVA0LHly2tMR6GY
7+46h6CsAEWUmOEyPPwH650RhiesyOnDY9oirNkMV6ejWV7GUdi9cdJaitcNpd4m4LgtR2xJJS25
RSwIUSvKNCuzTfuHol1ucE5c6P8l0c4ji7AAvwvVDfsBFEss0G5mQ9Q5c3g+JWF9gu0QugQRpk0z
VrOfgjU+32d2/DEGsCSJEt/89jXXUH5CnAHNhyFnMHzQJitjtaD3ZOzs6N7X9fNOysMCaBKQPGlH
dw34aP9VmHFTP/lV3YOSl0FXobfntt3Fe0nyHV+DX1czfBHvnQiQRO0dDrrcvS6rl9PSwjF5qju8
dJ9ZeprBDE2c8ZQudl8SJAK9WRtTaOtT65hF3F5aeYM3MJkZAS/FGab2PEHsrtxedtXwYBtavtWT
6hSagsT82AqW6YI1X9VdRoBTm0185LNKHoUyJQTjNW5fwpsZlypqTmSg7RHBVMKzPvqbcnla4EXA
WzdxagqhJQqpFgHo9tSSjOp4dyslwOrwZnKnVTfBPsSAtRf4aKXv+WC/vK5thG4GlZ75uyNCl19B
seTR7n05kxzMO5jEgYJuV/7rbw0cfaju1JVVIUL9qgrNwbNvLRRvNEowIZuGBrefOKz6vNJhMOAr
fT/Abo1WIAJ9rPW12Hf90pFRglFHQoznlvpJWhmereMlHC48f9ky28VTqJdrP/xoZtsDa0huyV6J
bRbDs8d5iyCFSgS6IYM6+JL0ty8TwqsNEj740Ts1LcS8rrPogotIPLroVz+rVRc8L7f8voTD01Tv
rwkRbHvzv6fMj4kHP5Cx2G/F+iiMmxg3Sk5xRCcDhuQZleJ4jv+Hwec4rNfSSbxIR/W3WJ5t3H2d
4dGcprjRaCnBpyLXB5/d26ksyTD1g6cnEgM6s3Oil12Yk9sNIP2VAPNeMRG8/jZCUInuxjIS1uUN
cvcpUVKtqZLh/Su74g7uPc+uF0taE093GBLpZwiIrE3l4MSCBoajgMhhb16EyoYGEdbFMuTanP5z
i/+Xc2n09F6rWx9g8ELKOX4MOJhrADu98QK5yGlpq60OmKb0IwrXXuF6bELKz/UB6cSm2Iffp5a6
I56962nXnh9mvlA4fSE2Ha2Jjueub0Z8AZPgLkhUrUN//xcQAuhSbbs/RceJ9BssA9aMCP9t9mF6
1B31bKBeB4YiJF53dv7FRY9DJvXwzq3s9opeERr3t1bWZt4pJWhV30wdog/+OCZdBs1nZGizYixr
dAl6281IWreQ1TwIvJd7xRMlJPTnVC9p0QbaixumjYgxPqWlAz6jx53KtAKIl/40y+B6YXbCFoY7
9/lOio3n+UoQSr37JZsErShTTNk8Sbzm59v5Rim5BkR1YVyDnVE/OurxsVatPZsh0PTSi+bez5pZ
Va4RWNPffsqUkDu9roS9Qc28aFS/mBSlJSTH3ZWIa1uyx9OfWflBqRuIJ2DN7Rf2EGqeNoaQ+27V
auTj2SL21yM+3xakqTNxQ87V5umhuwJIY6SIhbvk9IWoVKRrQz4thpgZurVKrNNRYQYz3zs+XjaX
IkYBn/B7uhuaDrNEjNdFKF1nX6jRQgR1tpAwrXG9Y7/ShnpNvayy33DmmhIQhzdcc3HFxhsJjIBX
snVf3Zj2BfK+Yh40SmraDFry5x8jFV0ISTl7R9sHDq47QGRGU/PP+JjkzBY1KY7jCcJmSf5+n1FS
gxq+SRr0XnP0/HC1i6jttV1p65CQ78k6pvxH5bPvtYIEGKuG901IFFA0JQ3kQL35fc9fMZ1qKP6T
hQvLKRbZA6Za+BdXHyv7LADeodf03mqNQdRgirwWQUL+ObsUWTYFyETp3rn8B1u1AjR5zWarCven
DsoS/yTTf1sbxyjIEMv1gJ55mqR0/UGs4umtdhLIvT499QPe3Jm6BNH15ymiHDncq4O5L7vAjk7E
d2HJgFnlYU4gzAEXkmcuIjFGn3IFRq4XJMHn96j9pyGElie8+pD8Ea8+RG4r+sxjipab45TAD3Wq
MIN2lzV148SC6Pub2C7XIf1bmTAGhjNw6lzgc8KFjbZXu+elIYzB+goFdBS12/PTPiKLndLt01AK
MHLdfTUWgahIsscSCUn9639VSBRkXYY5FO4FWZpH6ChjS1RaqxTMct9QiP+0jmSiOKKaLIGHft06
66GtwIuhm4IcQfDHGexbJlnnrqBQ9AEnCiz9K9ZuZI/Y3qDHqfHSunqqvmBUjgIp21HPIyYojIm5
mmDf53Oiq/37bx0AI+ItaggfTlBNU2VlXXeToQcVSm6OKnPBD3gXzBDJi6QywcS7MtAapkl8IJ8C
k7WJnBAoWuhdEHZ3lT8nprR9FrBxP5CGPEwRZxMu/BTtsqfG7/0Kgp33DMO9yY7+SjrYk+uioeNQ
acRlOq8JQs8Fx0QGWseuhDsrT7t2sZrlbOJgiPjGCGRFUrDltvwM0BgvSo9EO5m+fmNSNE897mhS
oVzQaycFf0Li6sGlfrMBvf+JLrXzCMENIoPLjoUMGj1l/SCT9a7oelniMAInvZtyXbatZAFvavrf
dHcZLbqhYp3Xi0ESCJKclpbjjFv+U75KCoxjN8k7O9wC6ymQ0fzQQEa/jxDnxFwKrLhkRreYpo3V
Y98swcLdhcPCKNIHyvxNE+eC2UtMRm+P2rU4VFou81WOy1NXZiRKDjY2UFTQhNnqapsdSsCiUang
CPdM6EHz7bc8r7sht33ZRnD7ePFep+1g9g1sPuRziweqTimZmptqAW/LQHW+C8zEiE3mrFMD3MIH
bCth3n4xDYyaMol/ilhi9a+ZuWHGZznvNKYdCq6DmEIXnRsE1nd+rxmWDEGQL8svk/A9lJnnowtP
MCotvPsfwtaIag4oewlKaBCCAaaWjDetuXifBsVFKcwPhdR531DNR4WwNBewmOPVYdKLVHhmlNYv
GS35hFVj4DCwMLzLQxFBapGx/8tJfjPlsw1Uf/AFS3sjE/Y3LEPj7kmXZWYC+9qkjSJ3arKLiwaZ
mN5wZ7Ui87Jx5JagGxTWkGEb0RfW2tgoeDBoc+pNdaiuHttc8CBsd6B+nfkBGMw5I6cLaDn1gZxE
mej3/fLa/MreFl6Au/vKddVwQUfM0ySTHhsJ+MwrwtszuHfgUmyYhX55ByiPXjml4Fu/aoShwzWp
skc9sNv4GG7r7BXcZe4h+kiGBthrpxEUJaOs9kXR9L/fANAv52/hViDPIalSPl76NuJN3XQ/i/Yl
GmODIIvYr/NWtHE764yn5elT0HI3xQGv88uQN0Sa5NjeBL6Gs58otejNYlkjEjLnaCZ4rMUT2UCL
j6nVeHSsPfci5olio9ZLG+G5mQNETaOrQyo7uPAwsqGC2FFlom7uWaBYlFaJK6wivA/waR/Y/tqr
b6RcK8KL/JGdcxRNtb/P08f0jyirk2FcC42NwJWFmSdCQdlK7j6D6WPzgU2e814BmMP24/GZpFek
3Kxp0zsX0+tyO+CC7TdClnIeuFA6vm6Wk4vbkUNeBR5X6Z/6XCSohh2ETbn5NgApj0EOtNigV9GV
nwkR+N5XPV+JR9FKSS1KLyQuxG1mQI6QHfv4ySuloh1iuc1rygWEeDgFvNxKHiaZ4F/wji05jBnj
uQCjVOGhF1pRRsIcTr3xzJ0rI2Um/vDzCMXu76HQWNPedQQjH4/aRGgmBBVqqiAHAuHiYnupxTgF
rVRsRcR1ySIvxQrArFmJk53fjN5JhQbHYf93XEV0v8LD8hyomlMw4rKbSxU0g//GQxEJaXdgHprt
EaFKPcej2CYsgKePSzRFkiQ4Bwk81HAKsM1StgkJRHbZUPPcome9aCqD1hqmRGSQh8QcdbBXLlVU
SG0acH6O2MGNzp2OwFL9Ufdce8JAcQaSA/R2ob44HgmgTH1H1ojNgXct0diFp/SsOWo6x47eXzuO
tWTA7JQivzqzaNESHSu/N0OBgIFKHj4ukdb0NgzkOP4KY+0eVURqiX4yen12E1/MQgGwcEJmzP1Y
7UYViKbM8XW1Q5XyjoncC62q5BMcaOS3/fVM08+HGTPQ1ICYBEQTcFQRd5d9vdGLoqG3VeGDYA21
Scez3UCLHAWMwcf5Cr7pBSyjAiyoHyRWzSFUPyhn8xjUCqwukzsPCsGRP6io8rCkjowUgV1Gc3in
thoW65VQRDD5eriRM0ClneNUrFzBvoWNSPiY8D7iXAQwzWDCzoUG+CVKgvxlbY+wCh2woFFKnorD
14WtSFW2n0BMuNjLeGKJeAGLNaib/AVUuwuDhTnkNZgzRqUoNn/hq1hoajJ0A+5J/cUV2W034EMt
ticaNw5j96VYCNWEW35oLQdl5/YWtkoP9vdhw2GFzev96cYPcsIeQiGIqWIoF8WBhOhI9bbt1yTS
SMc4+JdKLyXDyPjSP1fYF7VBJ8K/6uMfHcSAVJraCzp42Z//Jq6UfeTXeVCaI7GcT8QcK/Pdttls
SIcJ1aTADbpSOM/ovKqAHFZT8i6TovM3rSYMgVMP4d5s1APTZ4Z2zfoC8gim315D4X+EYPAsyYbF
1nbE5ShCMdIGf+Y+KXQ3I8HztroyNwKDmTJij9zUllnhEe5EpByk7Dppei73TPWejUFwIJUCDbti
AZHmc1rRIgrBBph03XujEp5nUEu5zAHSFV1DjNK14fMi4Q7qTuQF3bx6OLWoje+k5d5fAoiBiAVV
Tsuq8XqY5Dgt2PjzWzW5t/zwJ2uwm9TMq/oJdLe6UY/wPfuuQel0DYF1oHZ6ugjQ2saf9nBcq8jf
LDhPCW94UZ/6Bb60fHd62kBq3dFzmle4JRRQY7hyN4XWDG7N9YvVB5frpbjaTznDpo1r1LYUENYI
Uf0L03Hy76ygIz6hgJaVk8sOAAzdz8tfUuofy9nHhap2Zywk3AVBrUlWeDsTIg06LmvymfugqqNd
G+mHKSERvqRLfwbt+EWBnI+YhVave5fIg0HRF3G0gmtm/JgoFPaB2o1HHcPZMs5UUyvvLZNbo4sU
72hBatUFdj2+XvavAMb4TLFeHpBKTrSpxjUA7Ek/gNw99nAFTCLdltAjcAFAP3bG30STFGIVbDba
SY9OXMOqIlE0IdWvNysKhcUEdEwt8BiRRvXjtYKI3ag9YwK38gmHzYIvD38a945ECK8fz8ENCPUN
f9RIwkWrFqiiaYM8roCk/I+l6lJqcHGXi8uNzjaIymtHHJi2+2xu71R918RgVQdPjaMEbOWcXIgA
DHVoC0PYJQBcfKmiEGsXZ+gsmK01ywwnvopx32z51Zo6wAXtLQtDgwAv1t1gU5szlHpwgUyGqPYl
nXEgRUxltEJnDwqn62nJLprwCGUN9VVYQjOJHou1+q6dua2AzR5i424f7iBNrAp9iOgmD9Lb7UG6
QHJB5r+3GK+K7ztfqk/eIozc2eRcOf8FYOVWl3ed39+EW1SdrsKxojPeOsPxxSDnRfHn0Rf9XZDF
eJ5LwRIU3s3+w/cWrWYJK5wYxhgwc3NL8BSaRldTBYxyAIJLdZInmRO+VvluQRkxKujNSFunXv5Z
r7XyWjc9gz/apK9hQK6CoLCOnW5VsiwdQXqhyx9C5pH4FOa8eb4lTdRRlltBiTLnh2EhBn4mR/Du
lvMApZuSovyLpYsx12wOwcvLRK89gOQgGxrZeKVh/KV+egUeOLer/mkiNC350fxPKCPLUIkM5eDf
cR9CPP0v/MdWHp4dXMt+0nEDW5suRqDxmSbFIXq+Dzofg2kWM7lB5Ikhufz3VgizjGwedZDVUOS4
qhtfHarpGFxV1phtuu6Ibgunw0n0FyffCQuwms1GweOb9UjeMXTyMhoxNhYzRhixGVYJW3J/4SMV
448ig6oZJZ04J5U33j7ngNnfs8HtH1t6fTOqboL+/oooqX0GIyc+NlKeiqnaZ3HFh1vvErVbjP3i
6Q/f5wADeHTYpJjvCqwZH7Ub8sZmmer7WzpP6Tk5Z4vPks78eatJY7GH6imaHMiQ3JauvhBO5tvS
UMBKfIFLjkM8t2wCL9BEbHQyPk5lTSjlxO+QmLwz0f/cFS95ywjDvz/h99dDjFSMVTDzEIu/is/6
HIzO6EAMvw1DiUi2apdQqStD7v8jLgLcy/A+uuH+g9TfsrFM9EIgtewffLP0RZxEbmzXsU/6bXcL
udnryMhgEgKvI/ee5gYGbgEGfi7ZoTPhk6q+qCI49/I6nO5iFo+pgpc7wu4UYUUIpAIBgqdKXODE
O3nMZWOwMKoriEMjZetUGXI/pYyTiLbI/hMPYnWcqZkIvnP5AU+tI6XuQ1XmUII0GgbqZDXfo2q4
oIO+JaHt/heahbis8QlAmsAhIo34lAxnA3ZzSIlKgfVIEm9coU+LqwclHx42qC0A1xaTst71p1NP
QPAMJPItVde6HyV989mYaVgNXKBiLgFAYYDLwzPIFtBezMP3Ynld1KNA3WnRhzdUqTas92o7xKCu
rXwuXpBvfiANiX+SmHUVExk2mOx6lSPWMKOAYa/1PBC7vlm1hKClGAP0pQICzuAc1AjrTCZJ3aB3
H69bw18olnwiBhG+2hG7/sitBOBOFb7SgoA+PiLSRdD+ic7lQ41Wg9ud4jGzttP5VdIRqEeW2uHk
ZnAGdVbLmtVpFCvkAdyotR5CO11bCUKhvvNlKFI1bIWYviz1LOwxExTiUHmnJCQanpWqlvGWb7vZ
yQsQ8ZEuS3XHLBgLBgZxuOsZwRTciZlZy3lTZzObwkIHzj7xG9PFAGj1JQu6cucyvR87L2FUQUSm
AbqgOVT3XF6c/0vx4OhKdoeU50ayFhaVXnFSnGe2F/koWY9CGXmf9JvqSBEvZ8WAYr9/KJ8gEftZ
6uHXGnlBGR1HEjzcok+4grZ+Gar7ib5TuxeuAYwMjpukso30j91yMViw4lpdXm0pcKWNVCm6a9zp
c6vcdIbD1dZ5a7QHVEV7Jk/AQ+9tL3kebSKnvRqOJe9JHNO8y4SrU+o3LYEnrfd/ScUGlfDFQFai
MKTD/NynD5z41eHXynJH6kt8pKp3ZxjTmId3mTm0zritZ93f5RIfatQxQIRlPp6+EB8Gpqi950W4
6WUnYyhSkYndnhH7kE83chCxakGMFczs8qTQoa8+t/ozLaSQOvzLw3gmDeISzESQ1zoMNbueS2xM
kiTH8YGIoo2B+drNlEpZnCESGI7lQFOt5YYY21oBGKtspJ6YqC6sGX3/GXPbCcgWO4OQBfdK3EN+
VtPwqRFtN5ajNH1jv7MAA9amhTNlI/5cQs/rXMuP/Lg6Q/9X8ho50sP3HY4KluhiRFCoiwI0E4GU
tofkdYuElOoV6kmAUw4N11FnpVSB716OJqqBIf8MlSblfEfM35puXTqySaGrnRmb+ez3sbZTzrnY
PlpkNVqVxt6hyFm/FvU2nX2Q5RhVE6iHCDNO8UEwHBsvteiyJxIHXqSQshlMkFpvsCTbLc5BD8zr
IVX5n2w5eGsi7J6soSZvnD45tsNq1DgVLYwOIqGc4XqbNJbQXgGZCaFdtlUP4oxuHT+INXWRGqAI
lB4xc3QKvgb32vKApFCxmTYejixv8Rsdl1hPfjQ/NL68jj6y+FPu2uphv6xa8uxTJlUaAibj6GB0
amf+2EkJ93BelxRG3sOsakPUteMErCiy2+wh/w/r8/LnEjI5VUd90f3KvGEldS/FDiriL8aPmInW
6mLfStTnk8hv+0g2AOu9l2ziuye6BMd+axPS/vl8LVcuRbqkdoERjhrY1XapuVJT7rgPISzDhTWe
7QOy9elykdjxD7u3Q/rGY1G1CtPbrPmBcnrZzq4cl4siQFn4ekaLK+4seHeJJXccrFJRMw+aZOp7
Hdel1TaxUwYRiNuSGKsKqITmDaAawvi8xL9J3NM21b0lmWB4iTrFmqHCvPCuPEl/wSZOtPwSnEYo
+UxU3R23py2mpF5IWHq+lFapOrdQItnLlur9lTsmKG5sECkQ+fcb1jGepb/eijzOLS91K5e/HYWp
ysgfNHAM91/4xtEOGqs5Cs/bWeYK3i05Hcb5vmc2QOYeNTu0z3r+g6zqJM49Xx5jTfY07zV8ccgh
rl8b2oWR7Y8+QVjGl0svc1JkpXwt1c/QzTQ048L3+hRHVUrV1bLVeyAyHReUzCyZSftBlEPjXnRE
aA3jdusYJzJrjNzyIR7Hc6HMneSJxs7f06+0PTqE/En/x0XE0G4BnDEF3oxVV4rPCMsf6gYZXSpt
2epg+GCjcWVD+L/Sob3e5iKsjhm+NpchmqzuK57uXtqljHzoPGXqeIiBiVWXBXsSHclBdTZLAFQe
+fv2oLZMxNpESEjaEsy63rn53kLRGua0r5IyDRcDdjORli7R6ZX6/51wI+sT7p2740wUd9cIgx5l
Qt2gICEt3vPt9Uag/F5+3Az6e9LbEXiqA7TbUCLscAX1ZMTXIZs7HBDKsoRktdtGBkOY+RaHuIr3
m1lFmxCZoM5/rslSINhQfNbPUYJF7FAMgiDnirvy6pENF2FtiMfufERVrFawwm5VE/v6n3Ob+O2q
y/O5CRY7TaE9MPmk3fBA6r6iSt1EMrOHX5RpkCeW5eDUWU96sOmoQkS5X/3nFZTERtC6G3qLM/9r
IXmhfZOA84niDBij+Ca2ZeuDnNMxrAEMUQ3J4AUygJ+Y9o5GZEO5ezX73klBFgs/7zqlvDzyV41y
CZCpcGcPruY87nx0dieYqLfp6Y9Gp/wCX2QvOmQrO/eE/nHSQDnhkERZHQCGddCggQ777lgtpat7
UjYx8ZxhhmRczdWduqry9lbUnoMi4qy1qywTF8V7sdbej/2NTQUGEL0r2+kkH8frnf7kHuXl3eYr
VbUncsHg5TGJcicCImnoKpYUj0qE7fY5D1A/yHtGvkLC90k2xsUt7MsxVGkxhZPpHqnRrVm9iZAF
B+Wp+0ki/ttj2+zzJkRzqvRaQlw0wfpv5zqTvvZsi6/eGoLrcn5CsoufE8AuNqr5qiuOncl+aJdq
6eAGSXNQ7t/bu//nE2aDO5sIefdorbmd7h5bzB5WVA+QopTbL4GNS8suK7G+nR3CDKBy4ZBx3nO6
+oNf4o1xzwkvZQ31WX+oiTwfx2e3TRO9FPo8kdwBFQwG94Wc5sexQuxeTtrMTtDofa2z1EyevRX/
/8xnEYWXP9JKt6Oaard1PFV43gmFj4qhqLD6CKkzddjLv1Ee7G5lj7/nihyz+lFs6Ri9J5C9f9Yo
5Cx3AGdJ97Sa+HXCRNGSUGqiZxmFYsfByDTR7bMG1dsfiCW7Www3FLkHGh6+f0YHlyI8rJXrmOv0
ou6N4Qtv+15D0EfXYbWpNtRmmidb63rRWmJu6jM2oOhncJ18JvWgYgcUGlQasM+lWUM6vh5SnPvw
+wxSAsddsBotPye37988AfBggmiQv0t5iDJeXbNFyt4KDXzBjzEylvk9qLYJsNEs4L/rn69YA8bO
fTWKsqpv8X8DVZR1E3IRZszcST3XQqk8DW1eTBaYozYOgxgEPRmzKraMPewHwRgwSF8oa5phQazu
UJfNfi3sO2C2/acFugmaCPVKaU1bvHqvHRZeek5HB4uTcaElo9Xg+XiyNfEMLxUhbdolLNbxIS4W
J4JH70pLl7Q0TNJo45RYjNBI5cv3Zr8hpg3hGZRul9LIjWD46xlc7f2XwzbA6uObx213OCeF6QLX
+b1EXa6D0d2EfgsdHhKbPh2WVMyl7va4yW1l1Bl8wDddkdIMBZndaobqPLsIXUwoXY5EgPi8DArB
oV4RE0ETyhO/zrTMP9TOtMnhumdGA7IxvmOjgSeNoKJrXqQqhwyMNy2+LXxI97m3OOFbGd1cvSZD
xxSpLSw0xBZOuGzG/8rD8DPw0y9pUMpbgPCYoN3IcNm2Y9yLWIlWLTkpQ66Ewmt7PYprXGKPWrrH
3hyxJYnmc3c1fqK/fz0vNUm1NVmgIAL67dc3Kk0cqcGnLvA26vr3yTpRKJghWeMvtPIhjUTMGmL2
/JnRtdNKRW0VHfLiD/irh0PSnq26o2qNwCzaXqE6JMOm/87u+JvcKS5cGwBPMr5E4xBAtPgQi4WB
X9mGijHB4OY2v9tcHGG3U3K61XSjdhJbKstKXhkfAzo/WxHB6B3OOM0o5MgO6y5qqmsajpTVaCPD
MFMN7byYvVCAdd5u5JhfKdeRud4v+C7uhQUu1gncfSkw1EkMeJHYHyFQZ8MGJYiwHxy/Fpx+AL5a
ZMC36G4njhRl/IrsZCYwxHnzt7+j2As7L/aun7Ib/A6kzHGO7bS9QtT8mp5bxjePCIQTlYxilsFn
NFbAdC/KqwOFxKX/ObzwWvSsgK3pfOUo0YqRNsIbkb8EY1G4WkOdaLgfEW/1cDGD+7P93cRj8nqm
NaVEyDsm4guDhlSkKweoSq4KVdA8hB3HxzoHN6NojDv8o6dJOHMuhH/oqgm+AyiCcItltum5Sph6
vLIq1FKz9iQIl71NWIj4cxjIcWlZTC1X5eZ3dKpAXb5JJ8BF1FM8fe7aE201/0k87Q/fcHWvSm7C
mipQcOBwcAucAybtGvDNVNgaqZQEXfnmBilLMcpvXpNznrlOjKfPBMI2XffZPxGrlPcUj3DB/U94
masdYv84KXsCprx3DzJHADsCu1Y10A1vbfmS+nKl0ooAMpEE0dVH6FV1EfW75Fn+xr+H1MchfpAw
M6lpWEkzem7bCDxt1zdfAPvFyxkF6wR0UXHUdPdx5sMfyjNxMolrQZQBFSusM8kngLw/ZWp9kONX
GLxdzTzzfLXH93QziiNW2SkIrlLY1DEVL6DraDrR/WgXquisEbCueBxF827deKsoFxwic7dt4dV7
Fp/+UpRAxIebWX3qOenbBbFQSukfKY1YzuM/VjJxX1MESg/0O7xVOZEM+lBK6f1VTAY1YdPP89ue
H1uA2GtvCrqp/+9+UqtQ8L+Cx8awBWXIWvGDruoIB1guLcwI2qHLfQf4HV71Bmh6AywK2m0CN7bW
KAGF+7LFJPH671DDdbSlF1gGK20xdIMCdkeu9gGMQR9JPntuCIAHEiOmdGPg4KaOtE8ieeUG80uR
x6g8SLRClmjWY5K3bqs9WF2/Xx28AMrNpLLCWly/S3VzeZQzQL2c1I/yrqXqOc9mV21KPfJULOLB
bQW1boKo3FVTcLqAnXDiTBl6pBKJEbj713PyNExIj1MZp9QRYHuhqd+ONP24H840EqgTsovNB5Gl
u2V40rpx6ZXo5bOXs50Xn3OMcxaM6h8tJcdBSdFwrYC10v8YEFLyk2mY/fZImnBO7Ys31VRf4XM/
uc157hz24V3Ly1PCheMvbLvb4lLdE52pZv4uphoxViVoVRyA37QldbS7Yl7jvBfKhNmAN5yhDGBM
NLlHXhaH+7/vtTMEnEaRzHo28drVXagafM1hg8U6Q6ObNZq0Zs98NqhCY21DlDCB1SuNIJiE8UCb
xi7AeV9A0K1k4YiifiAh/e04ouXXGQdq68FdXhwoHKXmHbz93svx+qOhiPCJI65Z2UoYsAdN/30C
OGc0p6vLR76FCdv3u2yVCsibmS0jSg1hob/O5ncNzAbe6AEyNnx2IU2paFFgyjwZCb8bfmztq7cz
teoGNJfJ7e1H/gTPLZo+PO+b79j1a6gvLwrLA2I0mOkJT0qSQnvmMffdIJh8K0cmmGMpRCaHp5FQ
rN0ScaRiyqWeQzsSXYeIL/YrDVvVA2vF/XhCrfB5HH/K6sqOIaDbe17fHqgYO7RGkppYBqMKKNqq
+1EqdwySJNOdI62C0E9q76FT53keDaQB1iyFbS4y9Jfh7cZPpQA7SeT2kgJRTfon/4Q652CZ3J7B
dWuOHVgeLHXLexv4swWW7czDZjKuS/6XCEt8l1cza5Qt4cL4VvGiDBx7jVVEl14Ep5Svgko1E5LF
ZZ8b1nOLTkYifT/kaDVfm61JQmwRlXTFOs7T7JFw8JEGy4GpqyEtrPI4lrK4EZplhK+oj/vWu65t
dVW1QepPCKmaWVDcJ7LADYMwt9s9gS0yVJ7AHI0MRCY0IF8boERW8xQAoNklEs1pkzg+h6WiVYXa
WKfpnokHkHkd2Qnq/BBuRxkZ0CebKzMDP1diYQH0Sa3nQ/Ro5Bf1bPl+fG9z+3pwY3GBLq/+HeZH
NjxaABn+Ld2j+XnFC/fQYkkFokJuvX3mEBu2V2G/95Btv26aIRHRgjWFPE5joOEcwDDuATzoWTRw
EIupaUd9jF37vxHDPU45QWrI+QFSWDE0i3XftUE3dEceApU0W/gojGaFun9CsgFCT1uUsOTUHGiU
eYDgq+bUUzAuxLpXErF5Sh4uIfr+7H+LCFYwnQe9OHOmzCsV6hLGgtyM7/pqdM/CfhZeByD4LfhJ
h5TyJQ1DTD42Fmy0WHacI5X7XMLTgRbrdqOxIxIXxMWbY6Vc0YQqhoU3KdHfQQwxEP0ta93vBvNF
BpPEO6hPzVDgFS8O/Q/iVYfPmTm+4QPBhHGDYRfj92yRosk9fBCqH+NwKTFV21yDhSTZIfrHs92H
A0vW8Xm9VqohuarU9D/gXOwERHuYrRI6iyJ1AeqEyKseZTh0OA3sfIN0mPFouS77jAQ1ZoY7OWzK
DJUlTi0Cm4SjeFT7Jp2uCZ1EIKt++CvKAyx5ZyemyIGtnb8Dy4aRlghyh3S+vHaMxloLQpVfqyvp
jWTdXXGN3ABYihI4Y/v/G2+d8yAD03MksgU3RS3aEN4wROMhl2M5Fo/9NeSfJrPrtOo+osFxZylt
ZXXxDqyhhUnixuNRPaDQyTjTkzOiqErM2gHejIZ1a1gs4NWag97DohejYOz/4LVKS45GjG39uSvn
k3w9agDaPd4kgen0uBMKLIGbFbcvKRMO4/Aho3pynx7BgrlSomgBayTG9qDH6cpdKiKwQmS68x2L
4x0+5xpzqZjfPV9TrQKq+mKuRJt9XGhbwWj3PW1URaB6PV0wkjwRvIB+q1q4O8RrSf5oyjx9K1S+
yYMQhBwePDBP2BJHNUO5x8xZI9bTJo4sGs72kDSlnpO7W27K7YLxLQihG9maxTU/tZQcNljnB4rb
8Q9hdtO0Dvxmcf5+Y73pWQLVQ7AbATiMRDRQtiFy+0Q0zXxJHTLr9VOKIwAlOvGyjt7ZWqH2x4p5
pQ/qM6odTrrs/3gZ2NR1tJmDjdgYeG9N9Eu2NyEENTWCO32Y0K7fqDs1cFlTU553XlonrPft2jRC
3RkwgwPOG0UrMzN9UWCyBRwWN1bE2Wyhc6E0dYnNo3PkFQz9DFf/iZgHEBzGqeD9NhEXwVZcgsmG
vKhKg9SoBWoQPDeMvFeOEYyUuZgTzPhMRwGnEI00cGPV2qV8kpsZd9ATxJZhAq4iMBm8L7/KaEhF
cipA5hEIParPHXLYLSwbpAsDmJFjfN208c/kQEh1TV583pKHwJzNR4/d+1ZnALuyV/EIV9bt9EU1
v0fZzOq0hm/MNf/HkPah/M/DCpFbiG0WKitR5F7fM4Z3EYeEHGSOYEsNZ9dod88O9KBa07isfmbf
Cf5ZyQPYh+TEWvgOTmhPkYZUpdsPnmQfnxozq+N9jDge2YxhKrmJNO5nAcpmtJYbiJDWeUoA+zF3
vwI8k1dhH3Dt7M14hk2ZggjEU4cUt5hj0PoTEkzuRlzSZElLilMK3rZyjPbAxYC7XD+G+yZJDYgu
gtawBuz3xdOVPpV15yjIJsohJtAdoSCnFgeutXNHezplSZ3/tyBaJdaCngx7B/1z5WKri/Q0gRfU
RZLuCtjfSswhEnNUqWuAoclVC+KC4z5sN+CLcci58igy1S+gTK8OekjMWjS/WTbLdJyW0ZnHcAHm
XpRge08sc+S2abFbuJUUGGk5bYP5bKFIsVCocLStcjb0gyHNxQlK2Q2iHthiYzc1gyAt8sDvVpzd
hpiJWgqqx4WMTMg9xL0AvqWxlbpYSFIVS+QtWoq3xnunmKFr7itL4Mm3TRggH4noE1nVfU083S6F
UXyPtwtQUffuncRoxv1j29bxlTgtccBJYFszgfFKPHWHzBMq4sFIm4/+4aDOFGlWzy5YmqEm7eMX
pR/Jh1PgO01PdpkLzAW9DoVf6IE8QoiB9kPPbZEkTjh/Oqs5BgrdhRiVStnd6X4NFznueJVvlCLT
dwsHrXfogH/5Gr5fAlqQquuogzDe2Zgosc0UOmHT/ohlvP1NMq0nqGnsOeocdatEA2Wh0Griigwk
bu4zBH5/nA/KsTp8pt3dyIVzH1frHfqV/domFa6SmV2x8lPDn5LqDySPYBeQYDc84kjT7JV/sPbq
XvUB8uRIqtsWWwGV32TQmMyXm526C379+staGKf5WHlg5NPppIG2m9pUVd3t4I3Z7fnrnohPq5J/
PcFnsTNTmq3d62/dH9sBKzIb+Wb7Q7ui8lhkCRtlbEM6xK+NAoO5CfKU0P9jx0oaifuMHP1G5yQm
+oXmFTHvWQMn9PmZ6DoZjn6D3x46MLzGlHOXYHcKi5Gl1ouYX2BN2QX9k4r4UAhzFC/ZeDFsY2GY
w6IseXk3MTo/sgD2QIyY95rtweOiHyxzRf+iHlSNvMfSSHwUH5oKJKkTqGReYW1bENb+y+nd4KIo
1Q3pqeDsbxaDwFp2uV/yNFkN1xOIgHiEfxJWkRIB/5GzDwaLKaC9viAV8C+q/r5RK4EvaBRd/7lt
MJ4W1XyIqhs0xltSkh4xWChsCHUwf2e+st9leAhaeQT+IRBNpdrU5awCHZOHdi9zCeLNABpFVj0G
rJMS5aV8R+jXVink/+Su58d9gKONXN3pzbRG9mjErc/5DToZDFs7W1TpDx66lhzsCSFQOnXRcXoC
nRJ2qgQ68FqNnOAALu+Tc3DbqWt6U5a0Pm7AymHsB6eTtftJDL9OoYzdEEsz8iiXJ0JvY0fl9BmJ
RPxR/1hO+d8OO/o4j6GeJgNKHyFDVlKQJsFRlnyMhJTKuIOKQ1kjKsjKoMIA40t8slg91EnG/gP6
I+ZVavp9d+7UhV2oF631Ux/2djHTwGq67+1qWFKO6lgjSWfzr/SGXLeG/9h95/LIzbymVDiVbav0
eFz9J73a25fgnM6hiBiZInctSZHUM+PtiJ2oTAlAQVILu3VtzeNrMBHXe4CLAr/SRg1EtSHzG2d3
VFsblMKOfh0GCJmvAF4MN7Y8FwcyPoV3/5CX+EEZ4CdXot/+MgcTyrtB6SMnxyiBZpcPJPhGgSk8
3OU+9moQNS8CXQ64WwfE3pEX8e71gSLMReQnG1XsQcPCDlG0gvrwaRwvg2/sw4KZqo6r2yd+/pgm
j5IJ1CiCFgbdkM2iAfAoc6iMbr/wEJ4qfP6YUCn6uu7IkRNrpTGXyEM3qG0RMwy2eUbOlHQJnH73
haTv96VAMJioXxMgB9VP9LJh5IEQs2+jufe6BPxjXRItmLK4KauqEBycFGNgrDJprCMvuugWUQro
ObgtQbNRhdldv/zHb81s9vB5IlYg3Pyyg2XAhRAbCxqP/hWNI09dN0upi43EbXibnZNeIwY/IZuO
ySZG0B0sG13eT3gdPzUXit5hKGFHxnA5YDAfLnzXVvNOY+rh4sgf6CqmS9u3n7jWJXGcs0GGfKhW
fWTI7MHJVArzEN0r9rRn7aK4cygcSngWHBnA5CC//wjUYK9E6znwqaQhrqjw3IsbwPNGUexibKqR
Lbm/A2Wbh6E2Ksrzdilpq94da2jIIiZTFggc3Xx82/4YVxEzyUAoR6nbBliMsh6CUjX2oN5D6P/6
YtboqYhhTk1HDJ6Fjmn5c4oHHDG+6n0DoNF8q3i25fqXsgt194U0gGUnZsXQeli4ZdAQsM6FjPHZ
jJ4Bb1h+0JtJpwj2d57qOkfcz/wwUykMJAMYttnY9cqYiLV7jtOoJ25uidyLOCKaN+YRtoVH+oER
ciFT7jU7+4Aap+uMG4LrHv6uFf93mBZDaZHzmE3LgssjBHRup/JFvDV6NzFKG8g8RmDZe9y2xj2F
TddpdEegQbDrDTRq2maZ4BPyy2lpwSndBIV1oKSGPKVKT6fRWYjrIcWi30WbdpwLowsCxNx9EE0U
5ml1dhqCOrHAyKjY6Rr4FeJxBN0uJFw/k0/YSfUvMeParfgKaaZcd/TVjSSOrwI3NGSfeHXIZyQy
mEATzneyQh9Qhh4lzkLaloeYAl1QPTx+iAd5WpyDSqikAI3e7u+GjTTyejpr29ilLOqhTBolX8Ly
Ah+Rwf06raT+5QDcXZ2nk+luAR01bMlS4wyawLImGPIEwUxho9CbtrzDnmDf/5p+DwlreXSZoeaa
mqq6DUE9oqkYXK09N03k/PW2w4Yc+on7H/LrFojYGN9lsUB5oiccYsoA11JEE2115+jz4Jqtdvt0
cJVmQtz3E17nfeVhSjO/sUou6CWGOFN9gX7WgJ5yzbZZWX/eaYiDHJcmedemiIkwuURGS8XePgOF
40sBfZ0J9ZCkyBEDyyHgOfLdscRL2jgvLWis4/LTuJkdmkHX3DLscBmK0l/rotfGBtHKVOq97a3d
d4ajzstvCVXcEG00Cqi6tkDGVEk1eopgcroUN/eyvw8Lu9xfMTxSup63wOTiZZx7kdejR8JAIFxY
k4fQZH/xPJV8D7/yx6suyUyYF3n+JkpGPeLPGHORgO6PHjg8gWdTvRUu8yhI58ySq5Yhq1wkZgKN
cVg3lF6aG9ssK35C65F+fHlY6ps3q5kmleI0lM4wl9Wc+OZvxsIWWMiqJ6mjQCTLDIc7Q6pbRFcD
Kki+6sJTz7rfgQeAof+ZMt/97yEmHWLdrq2hrxglKt4nLlmvKbEJ30uW0q4g8Tme2+Jxariy08Eu
iuDBD9eae65zh4HPuK5COMz8f7J6zqlh8MBMOjH7nJaLSv6XxnUckS9HJQ1XrwHwZvn+zEXq5sMK
cbw+sa/fTfnTnQFnwS6AjK8MwjkH6Hmo65Gt3z2olwQwc1bfDJDVSb/ilnlPSfAVPeQBPvtrfw40
k49aIPhPC4SW8W3zrXmCesqulY/j10jXKwCf+GuQYvVT2S/n44DbaHMP7mNc5Kc4iBjRInri6vDe
Sm3Uy8rmZ7x8RyNBvIgGK0DyFKi1dXvQcyoJTlnmOwW6Efy4AJdYg9Z5CSgogAoDcruMaiSHqGeQ
KITwv3/3+sa//S91bik+gpvBGBsalxO9PU0wkxe/cc382ae4nsqV++EB2nXr3NvvFvFh6sGFTx2m
7rJrm+6rJfUvjPTPJWhUf/TCqNDA0s/+V9wQ+DyjpNzHAfO6dqk+ehflVrKQeMzI5DaqUpoX/4xr
CfGgSpMf3SDXtNb5IU+gewoZ9DvuNYXSM3YkhH6EAI0836jh4orQtIT060eQCLyTmcgv4SHpcnV7
8dRzj0wuF94qCinnKSs0PJ/XEr87FVJ0jYlD5qM3Hq02cSXT5LjAur7JmDslUh+xx8v9PCSnqL0J
k8EjOg3yQEbgX30Xl3hrLv5Npt6W+x96xjeUR6fNH8/O6eDl/5TYdnjYtrorSXUPc8CyKH6OlO+7
HTSUrnWP1F+5+gG04ju3NMhxc/89D2++yVVovCXnfM5+fNMYQrcL3tW9L3FcmIXqE93mcbgDd5U/
ngya+7km2g/8A5K5ZhaLId1p875RgXQZQdQuvo7EaFqIZmMqdG0R1WxYYnPFirACtw/PEWsqU6hw
OHC8ZfPQryhCxBUGc0r8/TaSdh3d2d+RDwO/es8oSOeQnPCaqyRX99HAOMpH9yNdOoqvIbJsRCxU
2jnNj6ulIMccy6lEjkqUsJxxpW/WaocDcNqcQ7dsJr0eFTIOWuLw4KUgQ2dluqCCdUu9FeMjxX1R
eNfbYh59SyQusoa7R5QcuHfe/MAWOtr+v6T6s+mMCXqW69qodI3JbKhQfWhW+3QINA+1v/WBkfgp
+Izm65clUSiuXHvPqKXumN6udELdotxTepyjYLfQLuldFQO7Gzb1YS39/HCNrdMdhOOY6xeQCfHU
tvrFDE2ns2LKbxCH9D1zFOlOfshlgCY+yoC4L5R180iOu5CAZtBk2AolQ38pakzK+8RylmEXgFFT
xPXltn6OZRZD9SbII6+iX4KD2I3EzxYRZ0QYrULGSp6ZRveA2hxO9li594KNUv3Wt7aTwEtU1zkx
krUhiQqMlhh2BPjp3M23mTDoOUWQhUbFYQH4hoOX5UnlYyGntgIzTfzYPYUz7k985NZnv4RkLl6S
FQZk4unqR0jDlzeKMsPL0PnEWHDe5FZ/SVgWkwg4o7ACTop2FsigMyN2kslfbh2Lx5F43aBOnNwP
EImuPzCdH+YSZNMBYcuilYFFyjHSOv3ihD+wETApfKO8k3IjgFJZ3LVTQrHDDsG3+BTr89nwKI4W
2aMzhVnxjHmMpdSNVnXtH9KMSnEAgf8fGY7Rvn/9jw5M34Hn6x02flVtmS/Ij7boGW9wDu8TuiRN
KT2N9ruuqKWC3jzRkr7arqQ4uXG+OoSe/TcDNLFpEoKHDByOI/7UpUlLvUCaOaMB2/fOun+aeigp
1OhITVKvggKBSTf7U8IfXVmUdLE4JwPa7kz/JR1QhrPJNsS10EwNDYTKVozYTSn3CLV3slY+ou0j
3Y7nqttWKDGNIM9iycHkMFqZb1s+0KTLUN+ZCWwxXOJ8MQCZDDxEU+k6BWyl8q1BOcOUc1SpF/yY
H+B6pz/1Gv9HbPp75X1aStiOYpDhOZ0I5vJNzcgSWMlVZpHZdT0e2LfMXfW0m0k1H4T6f0hdNSei
DgrComZ/ulXGhSbDFI0LbfUC9t/+UNizJgt1N/x5FmsdNvresXiDsg5kAgYFVX/go9KCbnqmeSUT
SVFX16bbbtRamlCiXkBZpg3OrLycPtsU11qsxQ0YGlcqBdxbUGiiZBpwwcVk0voNDM4K1fPYPS3I
Fh3ySUYxCCDNR/Ye7e0R9ebZ7FVFbjzcu/ZOiiiMNCfIqirTUU3siuuu9RV0LfEetQh/T7Dn/zgy
GxpqK/9+/BuHKz3BTz0a2VgerGT8mBi9+6nlu58lsF2GHfO97/qVU6EUzZchSiDAsvZKs8GU/OPa
c299TcxX0abTgUu1xs0p33zx5sYZ3cpEpygX3ZUsW3pe0zocpvjj9f+12Gjz/fmMSk/tMmEOIcPZ
TLDdYKuemY75EvsgsTfd0TDY6P9gb+qNEjY/wrm2MchavidVxeBXVGjYF34xnWRpVwBqbrdGtdeO
148Urj3KJ9H+RarbR0g9ewKnWjz1/a3dH1KPhDI6zmCDsZul7xZIS9gpNQBXA6SJ4rWhODEKHgo3
tbhT+/7bLXzPy9gyV1i7Bue571M2VTx36SGz6WLUPZA+HJ6t0l/cbneGO8QbJ7UGoqCsKWfoSRQY
OutCZR2jCNvYw1QH3fJcValitZgXxo70bY2ctgBDPpl7xB1SikyYPodiaDgGJUVKFaOtvUUnQNdb
Hat49QzL76j8alIKN73IIZziiN2vtdKoVOZ/6GSWzs7l5sPlpwbjAaJ72J2Ny98GKjF9zEQrj3O5
Fzx3HDZS1DcyLIuZxzOVVl0aIkL+1qA+nYXyw7thG/1giNdrIcQ4ubokJz5rpBAZxcUdZAFPcE3F
iwiyJu1qVOF5DWNHfQDerSdCkG4wOlEI4hAUnFd3wXotJ+AsiA2QnOHdsqg0gCRi/U7Pyw141RxA
YANXwbgMXGObwXJI7YRRFHxUCpqdShLjiNTSNerTw30URqsXjIAEfc3edGdSg01dx6wH9bIIpfq1
J1Y8vNNjt4Gv5jY1CdF/l+4uZYQs8JfjABQYTm3p/WxFnW0cTyCnZr7zl8ETditocaFvlwUfWf87
B8XFI7paeWHMvs8BZxJtNvMpdS7wu91onCrJg1nSB3EOiiAaVc1XhyLHbiFmRZ3WVM7u3acxW7ws
H6bh+H30jv3dZu53p6Vw97Henh5hYaCh67J3n8eGXtg/trP1d6V/JM7HHCgZlm20pu3Z3ftWh8Lf
UwwkyWCuBEW/I2qMdUjnT28TNEMRIDKShjkLb8e+g8PS12IRgRu8Bw58QCfUbUx+7OgkzEQ9Fuse
ygXJWY6WxIu0w6atUOwUP1vZs1D11j++ful+wyp4lzBJ40VAWuPo6pxuypirReYq5SGZ5a7Xqd2a
p4f2NBEuonjKT77zRFkvRAPSByQjpJipwg8TWtLppQNVeby8hmHIzFHDgDi6lbZ6hIhAZZnDEUmz
6sNNeOGHHwXiPzL1RghztIszoLqiJcsUMA1lcjqHXijbUTdlUFZkg63jZkIJOVd5FiMVvoLw6QjW
XmKPHv11ghAuXeYKzm/+2Ss7za1EXtF0BLUM9OGgqbXEJ3Hj9A/CDin9ziYH+87fk6PfRXEDDu28
8Zro3oVrCvEPkIyjg4nJ6KDkZaOARnrTJ4e5Nm2VYI/nPxAl6e+ZHGP4bL2QV04Dgshwh4iiqWe0
EL7Sb5JGJku8pDKXOhjdXWpGeWI9aW9U/2euBhQT4c7B8fp/EfK6ypuhahfD2PwghOYM39zNsgDl
vK2vHH+Qcrs6m2A0Cu41Ncx2oaNzNGufHZmj8z+/outSsXR6UZpAOqP2/EZ/WhWmcEqv2b1BmF68
o5QLTYU5NZNYVozDbldfMiVRJMxVDyZYgWZP7dCpTRq0RT6BCrOPkybTZScBoyyMbXKzPXR6rGFX
dg9NQefqP0BC1lbdXWK95E8kHUHf7lAXSzyO6/62gkqZrMlui1ZibZC52c7GwuO0L6rhRgwnYxLK
BpuQic6djxL3QIZcqLKuUM1LQp1+CLYBq5g6CHe9bITkJbJ0n0dvzFz97+ejrN0BrjLCUdbHJyZk
QMt4uaeTt5MST8A/TX+ml5EjXAPqfucIL0ZKfaiyX0c0aeLcppF5JxSHbqOrN7Wy4jcVk7TkC51J
ruCQ6F4ZW6Tq9pCdCtonLbSbjDjaHXjE7hFBd/27oap/nAgjK/b+nBr0pFDc+C7taZBcVQcOVoOt
AU6gKVuvWuVv3J8o49rPacJjz4seXYq3KQHf5k4LYKT6yO8XLZ/+g+QINuZ+mFZBrO9RnbSxTwde
fRC0npVkvAO2k2ymUpAzbiIrIXXvh4k+hjpTOwBd4hNnPje2JzUtF/tS3qYgt4I10vMwR6SIpI7I
hFayv0u6CXvmMa29Zip18jIWi4t/dBAqHCNpdazwpuExRN4xrjlGCtS3HePYnO9tX+sfGUtDPQur
ZIf3CwBB6kATU1gyD5N+nLJ05jVqmFkQ9wdZLFjYgTSArt8MHcyhfB9u9AgD20MOKAlimChHSstI
ZcgCxnWOWJFY0VeI/tZfDLSrTnYkcZ3H4Bl2TSBVtvANEiT79bcxdi9kKTPDLAeJ986u22Tj8gov
q6Dvcz1E4rgIeSJunL6k5Hu95wm6sTbjOwDnFZAQZ2OcNYFE8FjLOVBx+qSFTCpZwOTOgam/w77A
psZSytIwvG8+59nywNRP/sKiqtL0UGU2kMZSkXgVKlyS12oQG2LyBlJIdM8XM5u2xPyRcCXjc908
HwnTGGQfpG4CF3NpVM3eaptYAHuJVqEVaioCgEj7NJsTBPzfUCqK0a2WeUivz+DnZ6s2wxWYjYfx
4YqsIlbzPzemTqNR8iQjyqGLBO12f9pb6a0JW4TtEkdDTgneE2fo63EKMpUHzdSkYPc7NP/EtkpG
UOPkbHi+6J8bZ1dDKqi7mRZB0v6vArTxQf83AwNKIs3G/USD0djU1BR3TM976PN77ikxyXpmwPBn
jVY+BRYYW9q5ZNLA73vT8RUCH4wCfjGClWiUPpblq3EiFnkx8/IeAF7rDbTnR7REgviHoxeShI6X
mu4gPsJyfAzRgCRF8fWRf8+72d230bHV+0LPiMU2LFoQu2eVzUg1WDiY9uSsdR3rpH282+UkRReA
NQLPnhneQ87H8yXRrbDloUvSoN40ATZP+R/98I7JYWbI3D5faoUwA06sK2h5muTMN7wXkEkF8Igs
zHSnPUVTBHQU2L3CgZjh5qvKL2CVzjSSZKRwvyH4TH91zC754g2cxbFLFP2zHzXcehzNGtFGR8g5
DqN4Tx4+aqafsU1HqStMHQG3mfrb1Y+2WDEGqIxeJZbetCvHarHnkQ+t/lfykybHOR8byMwoopAf
oaxfvEPolhZMco1MAWP66UkZFwGoKg8SiLmAAlAuBBWDZCiLchI5OxUyR7kTG5ByaEuRH+btJt/Y
PwgmhntBLJ7abmoPs33pMdVPvCbF4SRTdX/Vdxh/JLGNwHVHvt/9W7xUrbnAktOkQAhZSUCsL7dQ
LlodXuP6CNgGED8uYru+X3FqAlxt8cV3Ta353VZL8frWA1BgJVDmWcyL9bGEHEXIkYa1dBQZxZyM
yX9g6LaGRdTqiSfCZ5UdIgXGz62ZN4BQCkxSsj7kNmMBNpv7hXvJNVkYm4uBZWPNgTRKqxyd7OPL
iwbatAx0fquRArzzDd02j6Fd6g7dRhYsKmh2yuGI4LbM135DBIGE5OEOcy2NdHSwLhwUXSh2DKF+
0J0C35WXr/qyLMavArv4hk4uOAhS2iKoe3qU++8wTgjPSC0ITJ21FOOTm50WKFrhfHuc90RndIyF
nvuKosyqKD5GJGu6nAE7spGahdd5fsewH43T1z5C18nGVTVxXGnNP8Zpk8WNjbPWYHTiUUeHREPY
vtsrOzrtyEue/owefjm0TSKek6kPDNJL+usrYU50hMZeW0yT5bXD2NEhoavBrzzhbzVLp1CW6ZcF
L7b92w0q4/IdYJOuNkQeDQDezMZyKtaF4DRjt2CGEIWiIA+DBFXd1NJzxTbpCEXdZV4EWZEcQQkI
K1O8dinSsZbNYbsRyHIcceNbvT5GMsCctatIJxvTEm1NDf4ffp/0uzsNKSuRZh8x15kB3Ccbmrnm
OhvbHPLvfxFfWznSCnKkQ3tTBkR94AXJiZ5rN0fx3jscZRPtnVKAGjdC7bFlzV9C+SkQgijfxeoE
lIyzBJ/NbfLjgX0wOe4luoIn3d6upW0DtrNykQib9KHLhhMDFOvZ0+nia9kZMiINEdjXrgTyX/rk
D0kIMs71zjyCR9bqfteHKOEhMZCVaVlCd8EQ90YSPrY583gwI3ca1MI2vuI4I4AWt3Im62qdkkKi
zxnB5/8jvqwJj3gVDFAVl0/2d1Tvmxp5xY/ZYL6qu6a3ZR6LIfk9Ki055XWKjzQ6rAij6pf6r9lw
5HNOWuHG+OjH7pZc/UTcVcR9EJOy6Z+vrTWFFeSq4KF/OTm8xeOgMDn5yJ3wTTpqXUvBKxzcedif
gHYez+D8j4DZr/wbncSWpV6Fb1cSUlD0ZRsPrxp0DD/zE4Zo9rY1KnMEkV1ClGwwmOIuMJbsg4dC
d/pPXXU9VpblBBJosnIYtUeKZtIlb/Sunn0VnZn+kHQZQwQTviyr9xEKIfBK9tEm9GMbedfY87kI
fejrVd0A0dpVHKU1LtfK4gXYpHSW5/eaxlfAVp76kAJz6a4aBBxsvSPcEwZCN6RrZDW4usn9c2ur
b217wPaG0UFiUbpUTlq7/luaFYvB72X2TYXTp+04pYuq2+KYzE1eUXIkQDohdRmqolvLyLu4gfDX
O0/8aqWfE/2fAQ7+7WPsTu4UhGKLHHK5+GI/JXLOPDY0k2WLFaZ4Dkp5nPdVayIVSPEiJnpgn1Bn
l6+a/5trzSbTuaa5Cpjme0m+zZQBu6MR0ZUIPhgW/W8dXeOaAV5oUSJ3ZzBeL8E/3lvFBps7OrgH
DcfrZe2c97VSK/sMttD9j3iShBXDpysnTITO6OOiI9R2cSQ36DS5LcL7ecI0AKKnxRL5+8KKA4Pl
BX9P5XpMw4hD+oUgm/YQ8wORkwg6J2kT6KhuCfLYRJKtbL8YBy2ZyfaZNWT3oKYLYFaD1xPKufv9
o0mKQhCoiZrm1+oLfdvGW3ga3iV3YoRhtostbi6Wd82F1zf1w4XI/WrjtzsTQKpjDotxZ8yeH9FM
IuO3dvkAS1y9PAmCGSeRF7VqMLI0/fKVfTHiCePmMwAHYFKB06t99j7QL9Fvnll49oASRQ42nZaN
GF7oLxgpfy6LNN0jkzY/hN6sKmMkQwtr2SvPdsPtAEhr39aHbFc0pWIaRoSgxSArMlQV6fraBH3l
HKjKpwjzQWK2lAEA6u5+SPDK07bEo2RYzOwA8xzV7oF4Lp2ZGwMJevC3kWW7yREhI5Yp0aTdWOIM
lmEvKw2fUGp/Ii5EmC2KWz5F8z8WIJZLXWYR5z6Z+Eq/QDik4O5bO+m1FcZ0EqCNioMRAIYVVOJh
DGp0o40lr6bCTsFjCU2fEhkLwpZEEGev1NOOYA+Fwbdz7MrGR4NEP5aYbgw01HxKQpY7leUq5XTC
Wgu/zGjnaDBc7+bRzPOzVQ5iOq32UDrJfDtCXECeZOKO87PyQ3Fl+cGviEXglxPzKHmQLQG2xOJq
LB65EdxmIWruBPGKZopuNhcPhx1KdotF4ZPyCI+zs1Zxo0pORYS7l1SYZsRu+XDV7s3eKIGYA8/g
S9CEfkMtuXeRml7jk9aJunIbVVOLUrmPEs0QVJYodqmJX2piGQN5Fdqm7ZRo4S4mz9+1458Zao0d
gEfz+hL9QW3nC+0/2Q02pNoSVF24C2Xhu3ltUiHCh2mUVo7tD/dsfFJS6RmkLSTHBnd3eW2kBamY
lJt7Y12pCmTsLn+VWuCLUtVf4siYQPlgwA0k7hhJAQvtfhpio6V+41oSSY4suk+RyjqfY1OQUIdu
rj/CMueWoptrYoNlGGUy31EqGSC3Pl7VS25UtjqINlT0oA2aFYet55vm+u0y5SLRXB3+4Wyw4t4M
CPReHU2hjJLlhuMsXeUBCRwJxTSUpIPZNdYvmy8TyuabwvR3hS/BY2f82aDHIOyZRpZF8LrbhbZT
oSxyzNZe0VEP3ozVrURM1CRh9jX2jsXr2VP5UBVqFESfY/3igYfDWXCU+/iIhafZajOcpGgcJZyf
qonhCluNOc0h5a/RF0YovIpJSK75KdSs9laYoEXubieo3+H1neHfzty69q1BQzLIh+bR4QS64YwX
8XQ5iBNnhsNf2c/hnwK6OW/fPBGbpBdYwoDtbMVTnnIh91F5NUHUM2CeLh+rdAWWM+OpoPMwA6vY
rxFjr9TBPW4SYPTTj80pI0fXroAYZGBPcoRBHBO327LtMa26TCxMdMxnI6wr87peg4xnmav1c3Z6
OMbqsu2qDyIZfx9Pg5CCdD3Z9XpLZRwxlamnllrRlbFpk9PCygCiWFCHpyFJ8sVGtOx/RInvM0yJ
JofDGjaA/s9cUcECL0NfLQI0ealK1H6voqQgrl8YQ+LcZZzdtUHcg32M+cLvH5Tr+rI+17Bev9ka
jb4HOT33zYTx/6xf1otlQk1nd6dYb8M9CboKqkGZLiWvaLJOe/y6THk7UKJR8tFMS851HHrM4box
dEqyvthkMBt3OhOcLo05EbVFZ1dN4qOzvDQBCNb+EkSXbuBgKb/ryO09LYjrxpydbrJYPwsttil2
qXA1PRX3U49SzBBQKcOSMdr8vIlSOoBiN4cF2fp7OXcL8qiKteiKwwPrSsQ3zaBhuy6YzSNuh0mf
annN+mUTcQOjxOlhLymk06gLJpyZSHbHpbsspWEBcjA240vIYN/NZqvxbcTwBGZ7+FncfhHWyVf3
td3s6ALB2TVZ7i/oXEKTk+Dk6g89uqaNI5upVt99VM16+XGirVQtxvgfeefM9qfA/LNrNirKSB9C
+NH0jvJxZIWdb4BlQR5rEHoc1Im1djeGaFD3u8e8EI+I/ES+Jmr4cTAGJULBVWriwQVmI8no/+Dj
ikm2R7cvAuD3TFkrRKk0Vl2zODqAO4GULQGMK+7nqYUXxVzEYbprFQTzGqpdDgfXfQwkUYARtM9c
L9fPTrLMJ72UqaTgEBjGRbLIilTZwSCKw80+yri+LThNNyTXzfAnv44jK/OFHzLGZfZAs3v/tpX/
NEyUeQbLZmrJyx74+uoYJpr9uykwt0QZWKHNttUI/0r58Dmkbiu/fRPC2l9yo/q3C+Xdx0byabgt
Kk4hUOa3R58zUkKK1boypkcwBEhXJcPhKbDOIXFOGcWTaN0DlUDqrKb+hBlss9lTmUAGKMlBPt8J
zaTSBTolQ8JC1pX7I0o0ZBVUHv6gd1ViIjCrhDZPfRa3gWSqnUsvrn1vdk/wuqIZk4njIRhHPiFn
iIl/VIjZ177iPjVHisyyJfzOGZerHrSuNszFeE5O+7wi0uXFe598yPQ8IpFGQqwvHAnMMoQ6NdYX
lGnESAn7ZJZrEdfLCDwsyPo7uC1v4MOVx0KdEor35Y2Ye2rpqDY5FW7lnTIvQjhF4+/AbKYeXsvd
HJTzi1Hy5D4MUl+M0IbsvTBi4MwQvLnCDSUQJm/IfPL1HW71vbK1Q1WwxJilrkqTCAkcnJjfWMsN
QmQdM9aFYkHpTDpP8eD/aizYQzelaRUo8WMWz11vNHJAz7zkkDBCFFV8Di9qn8u1PRHycTXM3ky1
4HrQeWd5mfCr3PsdRCZMxyq9P8E58QUhiKzDBUDX+deI/8wnNyjh5JGO8Xi4vY4glY+L/wy/tRl6
1sPoe5fbk4f/v2NWJDoPkSPRWZNOvaDIrCDQCtNxv/Z/lRmhew4QoS9myyUx5Kuumdiu8Ep7qKBc
U2jpBYDn+N40e5AjHPQ7rMgbl2eUAmEo/bKC1T2OuZqNpW585YM+v+Et9KoNHLfr71pUQISgocmH
hGsJDZOXKgaiJ0HcvKS7daIF2hwXVNjnr3SdTjexUcSl0KSSbf+mJggPw8pOhkrZlls5MvqUBy+K
pZPn/9kVN1CMcPkbttBSog1q+o1BUtArdc29N4+MSK+Q3a898TIg8b37QHHl6yENTY45wnO1gxK5
GyksQtRWZ1ZnroIWZqRK1lUxliVWsHjVmqMSSdYAMnd6+u7ImvSESmzgsHipFYdIsg51DQgjC2EY
VxCP54kuML4FbD64Xu+JggPA+EZvPU5dIxiPY7HXFlVzFDGyM4zG6t6ByJV3pmOAahTII69lAKXi
tHpRrfdNE/I8Oo6iYDwjmY7W3MndpSJ1/vQeejSzYc94eziWShpZMS0wBlxIzs2byk78ioD0JaUH
I4tFfJ4VZqFVlHSlJSbNU6RA0eYQD1VCq7zghSaI+7m7NyitoMZpxtL3xMO34FdBiaTSUt3VRfjw
ep5RnKyPJUSf1Ologox/lcJNFcu4h1a808FYFB8HHNWkdl7dppnIGRYQdsTMSl5pOJf/5I3IXOEZ
L8UuEOBNefFrk3b8d1Ow+woOQ7+OUp7EhsYb8WqZcL4tiVrRG+pVuUg1HNcXLvG2eAvg9YApjD3c
TasAFNSbqSmlgfTVkrmMsz8ImRmZX8BMudN09pO6i1mT5OfYR/xkRHz+Jn2w14QOeLOfzOlzrSPk
sIeoGWxW+VJkKXHqHNHtwZiotFZIBqkNXdcSiE1NlPc3VRschVVupe6wiZ9E1J2V1wC1iUXjapKE
CxYLJ4fhQHDa4njzfQn4kefqOa8sv6M3cojyNJQ5axrJT76J+5bYYjWMOVq5AldfE9TEnpbvnmxu
ZkFwUhf7Rd5yzSi4w+PIp1r6m/SrECW8bFHQXXuG+oy8Loy3crFIDL+fgYHpJ9bo8Q5tMaYGUwzT
n+DuhwCLX5CC8WdjReOmwCCYmYanWvxxyrA/JYcRGdbGwKS35I5pfrFvAS4hYtHhZpqrGEGn8U05
eRtnpVOX5prKjkCOwCsphi6/vSVoGHAgbhkSC+ld25KVqu7SLSW6BpvlaWPT51hbLwcp6EqKm9Zt
7coDzxJjmSbyXNd+xqtn+aJlhZNNiygsJ7i0sLRIUYIuf58l6iUArvDES7bDl4ZQhw/SmRmLDTeW
Tqm08F3uwilpsRrO6egJKdNFNZhUm3NfJZ5Wax8xnCXZHpsQRuF2YowhJ7+luK+FNKoQPZ2HKZlV
uns4B/rtuxqY/4x0KsLJAejeD7rP0OGoZyYVrFHYyAA9rQuRF12EpMW75LaO8mWTKHsf73nYEXvs
cCJ88kaWICGOFm8K7Aluqkc/913sW13XKcqEaDakjm2Ge+TolIqw3T9cA1KrZp6+pqD6Cq4lfbE6
SqRLj8hrkXCKLYXI5OrmbKVyCRT9LHngIIsVWGVaurE1lYM6dqh2mldcgTkAGqKT+aKmw8LYq7y1
wvf5PjKSvjtKu5Z5ybmoD7gnuKLKh8njPWhgq5lnQeCK2a9sRmAeQlr4wmOsOoyOa/BeH1WovSHu
xvrl7aqlHSrREIIDCpXaNt3QZFPc7HXdmYtkWizhRmZK2kYE1BynrG0xyP4bSfXoopLUy1srl+9G
UVWqp1MYF1FZGnWcnYU7hSALbe3ygMZ5lu9RGSNLloWA5FfzflYHwJqSQaboLoVR+i0FsrFjiFBV
jMHYQIsCn4LfLvOYQZ91+2Z0q87h2UKOS5on7L6eW/OB4wpG9mqglgfxEouPXDg9i1tVt1PR/tL/
Fb35xPDunkMoG7l41H3XgS0UWgne+9LG/UGzzbTqAqInUoMmjwM9zXTNITVSxDtBH0lhOl4PjV3H
WvdL8O9GG1SMkI54n68alU1oWV2HwYjroP2vK97HA8dg1APLKKuo2BfschD8NdwklwAbnQfbotlR
gJcdCnPog+xa7NKhDGrfY2tcZodnujDRwqpuv/P/XT6qmNzQ6c/75wHCWM0IYM6ZDceSBzpOT1P3
7VT56heS2CbgenCQ3iAGLRVbnivvAmx7E2UW211RulB3Qq7Ujy164qu955vNJfOjWgztGa6OxE/5
y/PJeJw7stFfDCjyz5VVF7r6TcQ58bYzBnzaXhiQOJSyiNWyhTYnl14giBhE/7ONAf07h6qRphU2
+uzGLV0wPLqf++wZGxD/COKXy3oTdOD5fbEHruru6KAIBlM+Ru9G+yCnNZsns2J6rrQf+CUuNYlL
a5cNFv8Tyc1mwSfENJhYDucE58KqdJCsWlLJJFT51n+5tqDQCvW+hrzmo5Egk+xLODE0VVqS44FV
Px343st2sqGA+hSvjvrD/6njEk8jDSJQ7+lXvBQXEdeh9ypC6X9XJV5IG++7XlZ94Imj79QRFRx0
mrivqESgbN1jtYHWLCefBpSp4xKmSwUtbjN7FQwgOhSYHjPiDcEhf8A6Ji5cMsDDC1xy5VufBY4n
fQMKv/z5/A5K7vidjf41Rx51pxogpXCjaqnZcgbnVFffnHAYw/rvAwIdTkZWJcl9de6niV23mmgc
queaOGeVaH0oMs76w5Wu8LAuFfIe+eLK4PoFcpESTrWv3sojdDgHK3UtVNyz7Ckg3sbaHRNrnvWf
o83toyF7gLrDtxqu8mgUEkkDnPVNzWHcpOKSUOstMnEgiNWcTapc0g6MEYDwisyy1FsJjfhidqeJ
xkp9Ix6kQ3pVXIzDae/snhAA9ON/MumqANNU2ZQs5QlGdGsZq40T4szZqM4zLLKfgA3HsDpuAYf9
XYM2jX0vbrZgjbz0bxaM/GdCpnnBiuOnhhg7UaZa9//6YEPxd8jryLFmPmawewPubTUMVr1JkmR+
T2pQENHIBKvaquzfE2MRE9VigpZLFq4S4kFxgC6MrYwiXpvZXq931RJHjmWdKf/gLacjC0jNt9fu
VTcAldYLARF1oLWh65OlbNvHcE2A/MVjK41aH+XEk2vskiDsIaQdAhfD33oo8uvXieyMOnPBwHUR
7cBEG2PsqYL5Lrzed+MzawGrjoReWm2Tp9+YhdO5K2BQHdatRzmDyh2T4VXKt2eVWwJMmUgC7nQS
IqUl9NIkRmjiG0FnmhdY6SK90rg6Hnb54mwmeeQ/xOiOCIuuVysTp7HCXl+buNVpPEo4+bazCJCL
fTzN3Voyam3UGzr56+7P6bXvigaFsES2fqYRoMyDm+pzmyywj+xLfjqBjcsyOD+FYWI/eyiMSwY/
t0D1KyWupIcs01rbUtv0ZChgUwdaoYBAN0MhN8Yk9SsE998m4EZ3d/UOEPiaA+kPI3vsggZ0h00Q
u/wkolmBOnPcUsmee3Sdwv/Cu5M8O5qK7VpPYzCdbE/pFA8gD1MSNtRW1+ins14ZMpgFnTgN7mdP
9brrgPkGmBboNc7MiZcdvBTbvwFNPq9rPz5zyvcsREq/SjWZhVUI8qbvxBrDPIzEYya3aSJtaJnB
lINprNlzf7WtuOEO/+reuWqYmIWCBs3G1oRZ0d/GsDA/tHGWG3OmLRgPhEm9LJg0p/KpDlF8Vhth
s7STalyj/9gn0Wxmd+Yber8n+JXQ9keuUgqbUz6hcdANDBI0BHhw+t7leXv/85Rd3YArO2631J4V
xvlrYaI7B4+QU2x2einWG+XN5kqk+jhjsCy3ICySye9rUNyHfOfuqM/M4ucTSqHQ86z+b97ETJDP
+h6RlQudZ4bRuTFuvTbB8Exfh9cPE7Z8gllMV6/MntYqb+OsiTONvYfmApCHp4qAMxBrpIKpDsx7
/zihnYEs22pI3RAB18ul6/TFDqUBuL56cHbN2hiOAv/GfKftICJ7Qc1NYCntCUKq2ApN6GHAFokn
5ygPkyY9LDcf73XJuqjb/ZfppurrUI8pasJgKNIabzNi8Fp4zG130yCf1DbqIuFVSjnWUYBI8sZI
SEBcjnG44DUk1wElrxz7c1OhzULQjqQ+oqIQBVEGJ3miRHfsfB/8eHoSmCkCibIMi5SQUqmANQAQ
f8SxlhwNuKW1inPAe1to/x3KPRBvMYoD1symYKm5eLLyFr8+hZ4Kbs5uN5Cny9/Cq8yjFTC1Lrbw
ivbSHFCjrOAv3aX4+BfnOsFp2eFyxGCa91It4Y9Gw7W1rKEwLEoVqU9/KuMLdWGkSF3aPsLak/38
ZxmcV4PHtI2r3Pwy6CN+n/G1DMyvVfOY3wZ54nJdlrUH3dP1YD0ePxzu4o8sLM0M6CYy01kaKBdF
cEB4tE3vdWHwtQf7LktNZ3yhkPDp+61XBdO8etqwkO4or0ipIfFS/h8451HPHvqoeFZmZcuLYota
HAvxRQbSNyRb2tWDb53fGY1CEqm7kE/A9UGVawQzDMkyvoSqg1vpl0Mbz/dGwG2im5vwfPfQRBWP
t5AdZeUTJEcQcQhDBVvIHD/xa+R5EqNB17lQ4SJWsef0WkD5FmnxbULrBs0eI6hUf+bYxzpTGnmL
kfIGhkfyNPHLhbgRSHKkw4wXRkrD1LMV091xN9wKkfcoMHbL/vnETvYgYwnJxU+xMqzlBwaKX/b9
MmhmE06qngzZLWNaYHFWi/rbKdOtzwxlqVqVLlFD8hGiqB9YBZFEtYRB0PT2X6HmfdmolQNx7I/A
MN0uJVIDV9hOrxFCBsFiFpv1jtXfDNA7vkLixhSxV0rPvtRNJYNzrjwFbJ5NBIPesEgVZdOpS334
ZbZyO815rA2VPrfCWtuxEs3KCdRP6s5bKIQD2L2CsyUke5NbQ8lWuHzQwAkZJDmhS37lL0yCIKfv
iCWIuLUfJjpj3EKcNKYEtsrKBsNnMEZvCmAFFp6tp0Q4BzdM+Oe+w3JA1QorWB7u5RJScVp1BR2Q
vok/Jxg7GyyR5xP2tdE3tE0FtD0SkBpAWATt4By0Cla/4+rJlP1Fvrt1LidgIKPj/oxv447J790y
CWAijacNurWpdqwYU1jMbkfDdwnfWM5aTSt3F50uvlB+BYxUBy4l5Qiq5ACLvbzn3ChoeAckKPRL
NdpdLFV99hbWDD159y97zM05oMIZmtMj17+/qu+FiGAyTRdzbt2hAgRs5OHnPkDLJItITGRDs5M4
akvQm6E50xOB2RammBhOgBPjetnt1FwFT4ahGsIAos0JzNw3OOH5+L8fkkr3amLIRjCPHoTrPI5B
rxgW5CNm9bY3Tc/w7Pb+lcI1SLCkBSTzMcmU3cznGqKiTkeBWQs3FlMiGyB8oMzv5kkbaA7qiQVr
4ltTQmakwIX25I66YR08LTwqhf5VBli/r/E9rmIzVReSIR/BqUE1I8owCUn8bFuQeP5cePn13Fzs
k0QgxYgODl0NUOoDAt9FuASlj0rB1e3v2w+w8M+zQIKxgCUb+EAaHK24bm0T7L92wXv3LImwD8YH
OMTFpciECVQdnQSY1MlZW0R4EL3GIThCt3a5vgbpI7sEBAPILQl2zpMwTUcoPFtd/Rqyg2LcOq/N
3qFooTg4IgoSQdXBFyrDLPP0tP2LHuDkuJamQG7aQZ/SFeM6QKeb3CG6wbG/JP17B/AvpdSEG3f1
dzwC1FQQcIEDdGnZX2srt3/B19U8kOOQdat0MHRWJ7eZX1rV2dkmaqNPkIg4zE3/WH/GQkFedUJ8
5/MWjGyJh+Y+tcdtG5VCE9yjyG3fXO65deLhYmXwpQXM1ZKjaFzLmqZiqdDTQPORIb5ghNr3PLLZ
RM/KGNXvnm23JpltOBPZMmW22D+FXn78Kn8rQiDnXsnLyCg/CUPhrvrysX/80xOdgskXHSFzBPWf
cXTSaxrzVSwxPRjVKr7Bk7FsXbCrCZp0vBqfGw3P4dvOJ6InSe2/T2m9e2+x1PjRRmFcy+rN97yX
tiejzsp3z17B6QVmYh6zrBAp8Hc1Ce4eQkcFJQbfO1eueHXv3htsuYNfLhVAtiQjNitvT2ik/FUt
qUPI1u8mjZIliOS6TDRAQ9ku2povqub20YXzrLmdGNP0186Xw7azZIg03vMh7tvLmsf/w2LlnKji
wBf+Xdo2WhcRfi62vrNzCfn6m9SMQoDMKG8Mowi1l2clzvCkkrQgCFQ6QqD9c+1UPhKVs3XfRH/n
zRWf06LOq1j+vCUC9WYkFAhuup6MsSyQ8N7vLu2SsPCWBJgGFrBNTKCuJ4XE3JXwBVR4LjWhznFB
acrji3AkTii+Nq0TiTbD/WS21dzb43u7SkmN6TC3KFnOuvCLTCYSmT+d5xvYVnFoBi3csU7sfw2H
QVzPJtzcmSp/GnewSyHfawj3fam7XtJROGUS3NmeU/THIheR+ia25ym0wtpH5sjaYy/53o4EV49m
SWRAeJcFCi6JS3oDZ18O8hefLZucUgkEQm86IDtxouKFfASE/3hEeC0Lot7t8Y2jtD+9WhSFWXg1
RtjNDtqer5uVX7L9HqH/yk251gxqKwGhEvujK28r0ZMi50TI/xWEBPGt/6ymPHXqRSJOw7eL5q3e
vdDI9IKiSGtT3JIrEAYTFv4oPTgdRgPtefrCaj/PI0XP8b6Ht+vV7BQD0uko6Zfsaor53vTBRQM0
1pYlatIIHAqJ4cUYIvdwWMSM/2cC1sKKq8nV/HRAqLD0VCxCzx/PCFRBd6RPeMcNbHov5DkWJprG
pPBfrAovu0FoiAKYMMosDbG34FCQqRKedF+T34MYZPbcpntgsH3OqZfwZtpJLRKl4KNHDi11Xi4t
OnIwo1FoJbIET+kh45ANa6UjlraVd6+ZSJfdUQsD33Wxj07SejkRI/4T7GhYXB4VocdHrpuaMSkt
PlkwacQCfXlGCUtUi7m6B9GGU4Mx8SosHryFZgQTZbXtuCBHMYW2ecKlutqjxYt+mcxRA91K/mYX
JHhMyHPk1XlFDdbIL+sPe9ylCKfgMhku6fRpTtKd2RWv9VBlotjAwtSOvCXwaexNpG+kTT8sUQOs
uJaNcA/odURtb+6Jz8rSFkEzyAM9yEko5j7o4vxjloKOeV6055pE/bGdaFURdFtWHteIonA0KUXB
ItUnN/u/W5OgnKUpc5zOx+W7EysAT8pbaHI/mW862P+jPsP3Z2vw6Fbipp9ZXw1yTYSwIg1UtrUx
FzRwsk4UCIlgSXLvG8OEnE8Qf/AqTMY5vgtMOw2b1N/KcSF9QHZYWjnJHla9E/74Q60x8rtTS/n5
ZlcBWLG7NIEhZ828qnMzhD9I2qRgVkUi99f61GY8ww/krDhivjcCYKwtyGkv7iZceDoe0eXiDjGY
5ONM351n+rpsrMCM7YPY0qy/HfXqj6kjRSxtgZOgKcYLrZlVPPKXV9kJ3IMFMUwstwSh2XLoi1Tz
aHg5PNqkWoJQIPVHq+IXy2NPeyhff81fscrrj3u+WtdEjEcpLh1CMOPqOCIxwEH7xGJcyoI6ORFS
WvLOiKXKLoG1eVTKSyv9bT8BRJxRzTiT6k+akDzCz3zhPZycDshunorMAG0WzuQNzsZFYrrBT/qz
6VCuMf117W4X+7dHhu0etLkGcrP7E7ihuf86A7XimuVRGMxmwQHmkF/thKJ8HZSCk4Ni9C1TWlc+
7Nxr0ImZzLWCWNqpIP4Yt9LZfjLo3D65SieplzjU4qpqveSbDn7pUIQMlZpg74kq0p0dWuAc5X0f
8ESdO3qQ1eO4blUxQ/6y0ibcqMCQxIFIXp2QiGs7o88pytAf8EU1mFho7zRSTzUuV5cUCGyE+SNX
Dymy1NFdxya+25tEMgHVRnQPmcgbo1Gm5z4CTEgkNwjhs5ekpkem/Er1eaLszlMlqy7JlYhB2q2S
LayQ4FQrAcXzdcZI9wdLqRDoFBfBy0RT4MZnkFZeRCNPn0YYW3MferFfiJp8xI1VzKkTWzCoXZTh
7RrOHep9R307T4E02tjpdIDXk8sR0BPo9i+QmcuOpXtNfMRxhjLuUWYqgqrN3uwtf07341Mh1Akb
8nD9YOZY0FRRMGczscJjiNJZhodjf5IOKHZ/5XOF/urvhISe4TM+jF81Y1PcZs+7iO7Im5NEIf0D
psHwcV6r6gzidhkEzo59T1oRdzcPa5lpwpvU7EX+M6Y72UfGuYQOoTZ2lAG3TiCjj73xVqJhs4vn
5UtSvA45pKgxXiTZGjKbaY+3uNztS/i9m6W3y8b1BH4MElSWREv1PpMPqlHm3lErYLqq9big+PAT
bGDBVnxjSBxeMLnD51Lru3Ti8jrATjVSCyilXLr9CcmwUClQVpAJE8EeS1bNPsTfgRrUfcBO7Hbh
6TiOqUNqkPVEAMGqUsG9F7gJPlH1fIaOe0V45xIe/SpECUXGMFpP9UXol28lU7GjI/k/PLEkaeWQ
n6txCJcqOkxNrLu3hGKCAFNoBMwNgD56fhQpjVQZ7VM12bIslQMfNt7jIFW8LQxLL9qvJlARQZrV
lOi5Re9EVqmh8yLO1IWOvY8nIHoR9AJmjlryEi2nooGS1boAeelc4lY8/GWrO4Nchnx9uRydYsnx
rSwdI8vZQB95WM+gM05XzchJVeDeN6cg1UnsYfyjvfSlcNkB/TU0QysuoFDy3fHTF3YJ9OTzKji2
x2OeoaLisTrLitOgmQneN3x+BoyJBh6lLgKp4T0MuTZCxHzEWQLeY7/aA5Bl12RcxuqFKXEMINtY
UDFxg/MpQnkyNIu1w5ML+HzS3s9x9V6bRt/qJ0XAqi7SDOdjcnCaImuDDEpfAaLcvgydj92vhSb7
mQd6rSoj1gFKowSak8D68cye9rF+RuDFLEaUP/fR0cEDogYCVjH9Y48a0UJxGbydxvOStHZA9ZXY
n2T0qhYrM+psBIXZlxFFHn14XIdY8982KyIn5x0AU5JEcIry6ZCs+IMuExOqlGawCj3wMKaeqE3H
RYKfrCs18IicKBxo3iWa4Qtuc4k9KuNXVkjGbaVm9Yur1CggZOA7pzbhJuJCViT00FYy5hqIngBn
qPYsENSqbo4I9g6OCFlvhpYvP3sqvUVxuL10YBa2giLbBWebEO4cn+yQ/xeILp0djmFxIim8cuUs
ASVZio2JTzLLl6CkhLqN0i1fuM1ZvGGSwY7hW194sgDDj3AUNE7UV4EKT2PdnmrSrsJCm9EFANxu
q32OK5VJOEGF7ghCJxMoqk8nWPMrOJ++aXviCe3NJ0mzjQIHSludb4rm2dXaRZwcliN7FWyrs7mM
L9p1/ZGTSDocfPjoYQaoxJLM8C/ifK+z0xa0wN1w2sC7vIt93gEw1BVIHqJRpUHTElwDvphQ9KsB
aGa2k3ThMHcY5868dTPapJy4w7F0Vjfmsjh4rMuPvplrQrub8xINDIG6KgNdhzP9qBw9LQEO+Jt6
8b95myFRlgN1NwkXat3ZO09KfGWshbz3JFWa2+njwdkEvEHXzCfR9TqHiMCMiieXIBTzkXZMoWA7
qN2ATueg+O7cSquLCEJM/q9StzkdMWM+vokBJj9NXuEveMW4MvZ3lLeAmyYnT1Fi6c2/IR8+MIGG
IUgAmU0VJTMCAH8cKITuxChFzBHZBjewKWjNe7qiboN693uw7B8uNRYI2PR6wXly5E30MZLZTZaV
HSniPwi+u4LC0LV6ILDWwtksJyOua2YllEBZA7W+Pw0feWXIgV8wDY8n69zwv4ztK7boMrWFNam5
bXCNAE/hbOpQ1hCQr5bx77q8f3nasE7MhTYoe5Nk6zVPcrB8fk7THj/3ug1j2x45hPPLpSld6zcR
xuQ2/aamMj0OVladaznWQvQQN9U9NR6I5UUvX0TzlFkv/jmk/istjzmfpIy0sblVprC7FwnpHlJN
Kncg9E0/ZSQH+jp5ESLRofKwCC7puR+9gqCPHsnRaROGTgLI3Wh3UFI9vROIwvdHdBsgdieBzJ5e
ojCIBA/sHRP4QjG9WBR2hJLEU5/SdkZ1ikiY3RE6PUGXjHTnC55mWWauHu90u96GOz/UJx5zvBnU
jRpC+8Da0UwkGqjdTTSf6DkJB1m/lyIjBuOk5bJ9p31q7OMTu7nJBzIPEnpktadxio8dRN59ngVQ
RbW972ADq8K4ju8FPkxlTSJptTvqaldCRnddIsftUfxRjB+owoCheg1umiwmsOAXtkZ5SUJ7erU7
58KS9GSGGGuGdJ5dxpEEc9UazFDximw4nek3pmmM08j8IBDCWK8G4D8gWPERwhvdL6AsDokhtHF5
RKm5G7QPlKd4C9Xn7BhoGJKjTHe7V3Umt0vPmNiL8k1tUWF4EnuUw+R/XVic3UtGPFIRxZ3y2Vg/
54jIMou5Ka9Uw+VzfNOL6xGrqLTWEWNOHZI/yhoV/x5yxZzFkIEt1/qzRBw9rMKDo/UF4WhAHKha
7/1nV7Tq0Y9mdHo99KHYHngPnz39rjKxPsmndSRavG6ErwN51V1UThIBo8vGqCa1sUM0KHWqEhJ4
L0347+l22RidDBXeNS8KmQ6GZK5VZVStXiBjj5n6T3GJcvLjgn2MwvaAM67IhDBKrCoFI3XleVQN
AADtCYqOKnzidQOm1AfiK2I7fIAcHanm2KWtqgwKP3DbEKDtfgwgyeTCRzNgmx7O1g+eMXisrbyn
ngWtMAtlsAQv4xlZBD/MVCbZwIOKPPXIWLlPlNVof5AuADLFf0B4DsxIgLZ28poIBb8wSu4/eR2n
J1ZPSKx28+gF0b3cqpi3vD1kaKkXrMQtjaT0GKKm9wdikf1rEE+UJZ8IDWd0oyLpcMBJbGjPrKKC
ay7GFTqQa8TmYWCuEfsXUYxjb44Za2LxpHnEDkLMZDZ53o3BHyLSAzKmC8UgJEjqdRwIdqfGQnVp
DVAHck3qzStsB4WFJa/6s4m26Xq6vv+HWO4SonsW+kx4OfldIo0e9nRiV+UzC71xOBoK3fmwuzpD
08tOu+8HZZxeJveSBfnwCUAf5t9lLsk8Nnh+khvakdBvtFsjMgz5mxqkiNGAPSIRHaz8rC8on8mf
x5RooOBq3S2WmLlSEReQUNe3CIL8HOmWPv9wZJTTFPsMVz2A1Lb7vqT3Gcz/icSM+FJSjaWsKOjR
Cpcj684070jIkwBHaKa8TMqXcunfIVYqtP8UsU0+0/bq4zFP0ZZujxm22oIWWBLZuysbjEmg4L51
9KpQYCG6oDb+Xmu8OXDs6q2xFiIVLHsY3xdrV7xQuq561nZ3TMSsP1fkIduN/5b3FUvmOJTqU7/C
sY7zv4NxsxgPPIGQi6snaLUyahpW+Sz8esTd3dbbYWYT9g1Xcu4I4QMVDGCmg6q+Mid58loJsBsP
DwVbFn7UJKdzrRfg1qzJ7biS2aJR91kUsz2fsPHsq6ZMs16XpYozfJPs7XxGlPPMz15ycFVJHmzd
SRkhIQh+KgJllHXVNDNJ0S+B3UvtD33MNbB9EQ3zj+KzbrRl4Oeev6ohh9kKuoPq/H2FWK6suDF5
viMlF54ph//x3E2v49LKrL7hMC8psPyvvxvts+Ye8K5IO1CRcOBkVI/N9yqycM66NWuofCkB4WQJ
3LUoxdFrUMWGXWURC8dfQuVg5IC4RE7TmSbArOW3fMCLivDYUhSsQoTk0EhwxS+rsao92LkdqoZw
nw/otKASBlP2U4g+qRplxqFsb8+KMtDwo/KWBvOfOJpOOC8ZZgXz7SBC2RNzIgpho+HVrCJWBWzJ
M1p+emmYVBzqGgBr4/R1P8UokYCfcxCCCmHRY1XF4RfYw1b/tJkSPrLcPidd1UNMroj7r4u7VvPW
m0wsHjEd9bp8NPbfxh7QYSPZ4XubPfGqVf19abA7oPmBBCoKstMyK2fN3qHlNXNoZmwCRDmWVZ25
SKDSkh8eQkv1lhg4Vpr0LIeoMwluXCkLriEtjijJc1GWrF1vgvRlKSEs0GadXh2GliExj18QAPcF
D0CA4Ga2vaXF1n45OY6GwqIFruwrexewraK9eC9fNDT6IdW12a2fKO0Rna5ZYU0B/hixDcarueic
pfm97++mANv9nm+vnKHiCxESxv1QDLmrlOreM0GV90nRCb4a17dq/I6weiovwtITHCWjGizEvQ7F
tKYgdKUbyzh3V7J0oPJZ3sX5K786X3BKllbfN1/M2xiXJ0O/Qw6ngsGKTXaDfZjwUV8MmE+RhWfT
Rb+fCVFF1EAZ2UQEViAaFZotroLtovoASgPrF6NL52xqvLTCuLdSqytJmk7GopyMV//qCUw6whQo
CFk2s7TFIYg7cMnUUVF/z7FwvY5ol90PBCPJaf9q5SXniGtxgaXWqO4zXKCw+UrwmmOL+I7GbIyd
rbEEUyPPE/ZWKF9PEqCNACTLFwqfnJxbapv8HdKLbgnHUAzM2j+0kVii5sSJKGUqtCQts1VtoVVw
96+XQgXJcxV9LGWQlCJMwyuwcwtGcC9lL+kJlirp4i8dp+0uBJtUXSUDzUasr4vUzkICJYZwvr10
ql7tK4zmaJZq0ZILxON+2C1sR+XcZG5bVSu3J7KIcAdy0tfY4fXDhASFOOK/tMqYPbhe1nmQ/0Ts
T409eBsulOf2o13kiTEMuSUiPsXQ9FMwaDz+eDAQHTZwSYaFqLTkLCPSjhcBUwp1mSrzNq2+1HSB
3IHWY1ika9aM3RhxehLW1UeDpCCjw2UG6KDhQebnBo3dA7hvx+oBx3x4MTO/H2tu9LZtDx5j/MaG
Zhh3oAtDA3PcWFjAkiSaOyVHds/XGNw3F89YkGNQR9VyElagSERUYuC47wDuCAuJcjugc+ECXfNX
im2CehF0C+Ur+SN7v5GNmEzzIYKRvr2HWBEa06MGvWxIPRebA7jQVMO5FlrrssVO5Vec6mbg/3zg
EKbm5uJsJ2fsTku2/kPl4oyIW2TJJqFRb2VgdJLKydGxx+hUWi6wcj6jXKFpYxAOr4XwDeUM5GRd
kH6impkDKQdMKymAcwp0eNAC+njRyAB0M+04MOwe+zlsevXxx7WQXG0KwWm1bG7FZXvLmq5wjJC4
gtw2cqDDgT0Y33rBgcnE2bcQzKNWvxifQnnP4WzuzizgvYQcksFFbvj2HmnecBBVKFgr/D/Z3Iu9
UHa6il9oiwFsjcIkS7zjXTj/VuIKCkWNKQrZLOgcOfKx2JRRZiof0EhRRT7HYvTldkSmwQHAdcPj
LAJhMT9xUOkT/gA8NiAHNWWmcXLwYmBjhGG08Zksc4ECPsFV1Qq2mKO0J0JTf3VZ9mF72LKwcJF1
htE/quUy39mzF4H1hvCw1JAui+72W+ClI9T0ed2QhKhDXKsk5fdPe2VScBQa4/ByOXoWhxku+Hkl
aky0SsNEKRuxoOcRRalDlsOauuDVtFIOo6AfkeaZ6f638jxDxRLkahvmcIxN18uXV/9gwDT07Rw+
XZZVYW3GeuEu0gYtGEJyLJO819RpOW8q5f2asMvzQG8dCWkaOZuDLAr6WutL79l27lAiUibDEeL2
zJKe1AjtyRPMF3R3i4fwctWRqgSl3+6FhWxYfomfAHYg95s0P1HXPB2EuFPsdxPjs+WVyB0xqZRO
tXJY8QQhNLmYhFZO+huHyCUngaG8MSBapngivuuUkn1YvsxExJQ9FEjfXha3QKEWEcYBtI+IPfEy
oDDA/yCgCQrWw9iY869/Bpgl5ynRZFBbxW5CnLJ0NYWo/3DaD4RHUYk84jN0OGG5PTenkvqGXy6B
sqqgFQBjj5+PyZrWB+NeFyfGuNadB2AxHfmZuKgZBNTKTTCMpLeMYZw91JTiwnk6mDZpt7yB0RDe
askxlxs1XfImoaJnesmCvEduvOcQUS16KPR9ERJeiR6Jg7gsOgwXa4HnEWqAAPublNk+3xhebPzZ
gj/aPKUUrrx6eQHl5Vy8vVjFIt0BWrHebpKCuEoX/iEDYyYkKYio/SZIoAgBFJ0C//i59hk5Yfa8
YjLsMA1y7Hi9Tc6ZcXKADXwIX9Km/okW2ms8mbpO8r5X9PShOkpWJIL/BRQi2kTWuiM33T94TTbG
AS/q1+wCYskSTwpi1OJJ6VCWcwI1LzX4CXWru2i+fD2MfPje9HbtHnlxL8N2Tbxx78jtHNg2ywM0
IviPBpl49yT+gxN1ncMuMTAQn0wZflpgz6ItR+R62ZPc0gJuSdv2RPsTm/SVZ19FbImv+HTGiSLL
TBIFegcIQIVDWb5XauKf6+I2TSafCwE8PQa10QldguOW6jCH23bC+Jvtn21hpQ+riFqxCneVBYsx
HIrXxZBKAuTQ3IlhtGTppAmTYFj7fxIFuCdv6elH2k+eiqPNC6srQIjuFOL+u9HRZDeBY9F3fg6U
mevTxZGFxBTFkaqP3mCHOlM4EGPGU31NrMUGu6fqVBCdUR2lZ+2RukW983wkiiVOh6CXn5McH19x
Sht6NeYmipB2yKpRSmb48LekQccJFJhTsxIOi/N0h/qb6GXWLL9PUCj3VHbvnStTLmDYRMX/EMEM
M+NrxyegHijlyllj4RPqeFE+vIA72LMkpawfm7+/wJijmQ3sv6z/1u+MCuYh0MWy1fBlzVqjdSbR
ncy4Ca3ns1EgqrM2NAJBfTs6qsGyRH4GTvokvQgR7OL7WUOqDdgK8ogxcPEYhI2cyKIkz0AZpkQT
ykIoZMnvo6cfYtWvVrL6oFiDgZjytHdo9RNYzF5hOF6wsuNF4hnAAmQIwsgu/RrkjBd2/zS4w9HZ
yl5Ok/LgWOwj8P6GM3TdgOybgIHW8swYTtbgX77PlhOR4XjE+SLdOEGq/UkBpBzm0nvENMbnuUU2
+zPfKsqTV566SPvCLSp1VMayS+UEgrU0oaFbQU+h72ynWOgf0RsyuZSJHCTDZoNG0QdZkPhUENbe
kUIfqv0ubSHYfnHUh/hAbKs+Ww7UeQ1ERIh679UVmymoVGR7eL5E3nXqim+l+taTvRko6lEFs2JC
wy3BwdSWFGz1Cgg21L2yUG++EavFSri1aagGJ94WQ5a2N1dE+gUABaMjPnQipuCMEsf6CR8LQfLD
RA4hG78Q6s0DszcQINLnZG8u3ctmDj9HPcgrmuL1Bz+ZDpvYTWQpPULxoljK8edDcCEQXQrVt8sM
8eNvUGRzagRlWQgleWMmb+AVwdQu4KpmwDhdq9DX/UkTzdaK1kJ8poVsI4CKbPl1H91q6MW6qlLD
Mx2FJ6U+7+JdSThMzuVVJZeN06JcVWF8SL6hI6ShmxUZ42piqbgQfqkBk8buuTZMkJ+MGzTT3RFM
qI5dHtQtXIbWeJWZuOwmHYXYon+nLcIbW+AjPrUEpZbjOECBkDKmTjLcE/z6DZk41uVDlfKrglph
jRpgHrRxiu/NnEELFidgEZuc+Yzv/nbZVW04al0e8I6oJ+J6ck+N0S2lHuGjK2EKAIny3yO6FCE8
ZtPsWEMm8jlwJy6gZgRo7ANL53e/D707vBBiR7z9Aqjm6E7scxKtMZdqSv8dyJ7nkxHt4bn47Vtx
uGIdsj4lXkY/iIAGgznHZlzbs8zxN8PZZn8A5hPU03mmkSdH+TTNRUOqDQPlbBZnk8iSggelclTt
3Ri7+4N0kjyAo3/RRh563tNz2EIgpzhJEZeB2CiovezRAtt6FjBuaHEOAivxdyKg5DjOEpmB39gW
dDK2dTjU3IAqhpISpwQXNuTAadDl8Q4UqBcbdhtsAONEwXzP23LVlMif/XEW4I6eQCTnwzdOmc2B
pFZf6pKwZyKvhPi5UTrKbCi+/jZl1zp8pF3bOLZ63lwnM0KTHEss1fx9O0+1g9OEH2nAXXD1G8oe
YesTZennSOLugBD1NnfyNDl5/xWSVV0AhP09Fh5tCNFb2EG/a/mAQCQeRMcqwvJG868fKcT2Aga0
pm+gDZ4gCM27DH9JZK7PBcz93+IGDvkUR1hAuLNAxfvJLKOIN3tAjoTyHAkAxHONXXT9XnXplc5o
usakz1Ba1L3BsdUWYBcpqyE2f+MdtjWBQMMXKk2WYmMtlouq/eRkI4ZM5o6DXj7VTPOknuhspEjM
lrRScZwU1qwdDOb8mNRGCkMuojE6I17ZzHb8VUfCW6wmWOav4s0qhycnzSDo/uHEtBUBZtSIOIDZ
fLK3p93sJuEqv8ZMqQnvtNveXVzQUzQ6t6Lr5EGt0WykGR5TDDhEVIM2pJifX2XQSRsdxDFeKWPS
bj/wkZCUHGFWqlIg8gy9pnt9ggIorlpjLFo9yXz3+ng/LY4OjGaJ6ys2srtaLN39mlbV97o3BNOL
XEzyW1PMJ6MMMIBLVxxE9nE7q2KiUwx53+JQ3u09pVgaZzvbhPKMzvwVAZxBiTg+NHgswk4K1/Fm
Ik5ltLTcjpvXhrkYHVs9vqpXHgYmSiGD/+p56rZLGYMBpsCZsquuq07WVc79/49JJe5nvMrlt32M
n3vKLh4v0U4u3Hs4iU5A3eO4oMG4CfuzpuT7sMnn/Nf53/Py4cf3GMyfJSXsh+jflA6KwQbXZYpq
KmaLPp3vZdLZwCnd97hkwqzzoQc0h2ts6R8rylfzbxlJdrzIkftzETL+oMljdZAMakBIU2bZKnWd
9m6dvJWfWilz8Of7AUCv4Sr6qMTw35Y1o/MpiXQdbGvwpbiOr2VzpIb+Ds0erR/5WZm+yLuLREua
S40R38paHlD0zCbtiIPbAPBTeXPuOTTs8YGDcwQyidaVqPhGKb8EGFzjgMGwZN1etoO7HflA+wF0
4e0oFjiTn+UBDkIJsrvaKu+L5/UExRP4duTqUA5cEV2k2NqX2N8ZcFdOgMd/JcEw4C6YxBP7I4ur
4KTKp3ooxdNOdub6gV3+KskgjmHKcJA6JNLx8o2/+cOjIl3gOaTNTxlArHBMhgRpzvj0c4/dGlEo
d3J3KBWflvpkl14Da53O9wlD4WuwxPjz8t4bdkuE+9sbE+58m8txAaE2+ZHqgiucWVtuwPCnZzbh
oWHhdTBjJnIXyQkMuNh7dVgfFOSOiQ50WRWIrA/GbgDGMl7kchem3KB9A7p8LLqbhbLIuk4XMawQ
Hxquo7qx72GbBJ+FzrzwmU3b0vRqpVjNzNkvAMKBTjYyi+VAYIqKiBUUX8NqMglZMFzjzyWN9HGR
BShnJD/5KbS7ycVr1Q+kKXYrj42jrGmCzVI1h6NDFhIUf7sNQ6ka9jEVpxDumxG/id/gbnrFD9fi
GOCeAVN53JHzvinSArRNTCo71rFwXvmgwQSKyNRrccbwXz/bIapASjUkEZAjZndrg+qt4+fw72rx
l/ianpVazDIboyBPfCPNdtOXVcPRgQWxA8L6qvRAoHGeXXfQBWMFH0d7rDrbds6caTyLUFN+Tz0a
XYT+s91BHdrLZIGCTS7in9vPvVOyNpv78GZtvVqNPr/DXqQBavuK0nlmVxZBm580gk1/x0/LvwTw
leTiFrYLKxqoBkfljfgnfqeH7bFULkExpUlNplHji0xGUwJ6xv6Nrd9n/ZcOOwdl4yTVI7a2Et6F
K4WeifgUqef6J0n/KwakGvAybacv6TO3nYB8js3zGgvKvAFKrj0SlU2gtue/Mh1lPAeknDnMNj+4
hrTH+0zUVzNzDxIzZHOPTWJvYnqwQMCSt7ER0e9NmEWbgKWjbLqEPH8ORVLWyuLwJUxgCN0v7rm5
ksfIQw49WTXO+DuN1j+tfKD9iFSlv93IIDfcqVT4q+3ADN1qBhmOU2BKwO9/4gCMSAQk/2WYb9e5
Qtx2tZ3fuC+pNvet51AD15PiG53PxH6y7mcNjcJ7mf7441qsJTc2+beV3PIRYEaLkBuicSk3yPBP
fQV2MwaptO3l5HIiTXn46iD8f5o6wUxdmwwhCZwjnzy8lFcDfVhg6frI7DMUFjAozPDF8refNwZe
ydDCLasEv5j40yEC5DuSt3zDEMYkBCaGYBmHMfJkVk3rpPULKQCEK2JWbd87P1i5WolplUfw55O4
mzmMLmLFrX0tum8M5Yjy8vGP/1Mbjz14H7Rf0GcEkr4r1EEtEzu5vK+jZDJPoza8CxtfuiltbGSP
qSAqzBZsRKHMCQpy9TYsUc5QKE1MiAckmXq0uVv5VsUYmEKU21OdF08CokXAQ5iF/KBTddRbom9r
cbCEAYKR5aFeFVls9XzVrHu3F4kI43C7QcZOxIlTK42eDJn5BnQmTSpCKU1YKKlyllqYYrOfLMXp
XRYITWl/kYDibREIXTzX/ricS0U+UN11Q2dj3KqZ9vvmwvarSG0BCoT0lgFMIjsf+xy3cTCXG2qx
jEMGDjG1fx+bQR/w7j5a8+UrI/SsLe3qzrQEQU75JejZG4aAmct53vLQbS0C4E8T2TzZcISjnsL1
mbGGT3SNGkaM0uYq1yu2jDfcgXUV1lw3hPLY+zvPU7mp3kNrj5ExiyM89PIkyZRHa/+9v+H1DhOw
WSTRa+vhvSRldTsf3cQ2duCwq1CAEH0bZ082+UppSh9t9Um0OsYU3di1Pyudxdiuo86MGOzrA2au
UPFyGVPxG/YdRF5Sw5p15rIhPYzMVOyHS4HEPbfihiz3x/i4IfE2P7+QvjAAU0usu7ACU+OZCfHW
K2vV7M14D1F1az25yXOIEbCiclAUJsK9M6kCLxnUcKqn63mr61PCnjxNM0oqNBNMEVcSUfp4Fomz
HfaPbyQgDcI8YcsVvk921X0/TfLuBUcL8Gy3+hYix44VMvgJZnP/9niqToU1ocs4OjBjiWMSuuXF
CQoV/25Ml4vupRYyq8kMA58Y8yCIrm6fjvhbbuRZ1biw94tEOu8dZXCc8+06DLbgXIETv7KzbZ83
+bPAPawwrl8rgjSTu3duCdsYgXcffpzor3ed2X/wdXewPVC1fBhT0JEXvqbYgQ20kOfExxKoBgqH
7Hn/jnAFRCnawgXkDG0/RMbNRBSyn89ROL02W9wOY1Lnl2peEF/uy9IjeE1rMtmk9kBoioDlLRdW
Byy8qnA7w9ixTospxC+2PLNZh7LcB6XqUbf4o/PSh4zv9p4Px0YtGEQSkOrtrIYDRDbXysU80F4L
fq9YqLd4ILyA40rkhKpnMt6xo84g34DhJVr91pJCofhc3Td3ZDuyD9z5ZkqPU6FZTK5U8O3ZBpHj
8eMyBNrlp0M7OU7fplemGRSpAT3KcZir2oLYSZhmylRLeNw6FTqQOKggpwe2/iDOW1V13SE2dKcj
cV87sRPGOAseJ+0/PuDC0mlR8l7MfoYlx4LtmKTijlkDXZU4mXbMoKhze/W/W0BvJ+UFXL66XCz4
dyFduPeWnI7B603FPObVGKasrzmMaJVBu2hC2Y6uPDB5pIw3DBPd8untvEq6jgtYAIGHIi/+jyTK
rzQYjdBUfy2975mH1iO+vcZMLixAVhq/wRrZCb666ZuRxfL7yz0Jqxc/JQP8dC9YkxJtDoMrMZ6I
EGB2+h6pMl9NpWQymCZNDmHjIooUgs69n88VvogUDvY/DuCpjoid3WBtDUegIG43PyD8Jxv7kRYf
mNmoEox+5JdKD6fufYUg1GxblYxFWU02PmEQZ4D3Tu4k4Roh0bTEss5mPk5V5odMceHAlJOCUM9v
BQYUZ+B7dePnFdRZTiel8DQcgRIFuPBErdy7PX0jy1pDmlaw5L1bY7byCG7e60SfkcN5RrhQ8+lk
IFaNdrcSpaBr5KcdtJD5TCLkHqooEIVD9nNDxRlshyWNR8eoo9jFBzwna5JFqR8sizfTwmgByPAq
pjhsK0HJ2M4NFEq9CmdKajZjM9K+BS3SQiHN1/pp75EYvmCb8s/IAnWhUhzcNNW1hPoiPVKYVn94
Db16ZtAHbAcIchUHmEspHIl+d9RlBrYT9exRhKaFHe2w+OcjKX3lQEnAlFGQ0KvAgeSXO0qCv2Q4
8J8dwxkw/0qbsaUXyoHZbiFh8RUpbGhtzAi60MRdQjLZu2OPKbLbNdOwuX233YYV6tPwfWIomcXu
su2RMsFLW2vw9J75XFucQPxpJ7P8F8obSAmIX+lxxDtielhT6bTR/mgMlNWvYFa+qZTduxt+030p
Rx5TN11UZ821xj2CzhhDzzavqZ2S44195rz4SVKYUb/KirNx1fcODxlFMBjVk+o3yunlLOtapVEf
/0lkwb7+TUJig3e27NM8lTlU8m7lJjR3fck/ava7D75E3O8r3Jyt7LCp78fLI0E28gDTOXjpL0wR
DQCJkjV7nF1FFEMx/ZgN455HBOkWmy/hrBs66e/ZUESayxwt9zbFtE8z2TY/f6gSwbo2q1SHgriS
p43D5LjaGoERWGRR15VQJJWJenhbKGiZo94zro1Dqq/dYprC2IDmraeC1Jsm/4Y3GL04PbWCjOkU
a2jT5jc4MqCtEzKXWrvh/223f7wwU2BUZj6hh4dPAmLxXxRr7AGCHbZxzGasVpE+xMConenst0Rz
7QWJiW/4R7GzL4RCB2R13kfreZjEq4splGmIvnb77rv1DQ63Ojq9kGId8CeA7rgv3fjoFDGnlFf9
8QjKW8Ttl+G0zL678ZO2nobLeT4MMtbwawi/f1T6v4UjrDNAvZt2QChDAOAqrVKizORRSgB97Kl+
KJRD+uO+wfZVb9WFk6OCr55rY1OKczi8CwozLv+SaUrK+ILqXWGIhEWwGeIVNZy1gMBoXSuYJaFy
alkrgXTNl6auL9l8VlZzDDWt7oPVGqamIyppBWwnUs/jr1Td3fHgLI/VipD+lrJTQoM0PHpRWuQ+
veXpqel+0t91t95E6CUmA/QB5D4IpH9SgLpyF427JeNP4Ym0MUGHKVZ3xkrWlL6KamUYZ3Gb2u0W
LyfYu9ZufzD4scXxH42JijBvS6SpfHUZilwRxyE/sVghUBoqPWktVX2lxlWahjw2/O6dDB45b++d
FPGCv2Vv4eNrRW18Pcv+j3yqCb9tnXlqkRY6x3eMrMiO+lN/0rOUpFOr7J+0YJO5rADsx/hyDI2r
ZyJ+YwH78rQQ5nfFfEGIka5Emb4TT2T1Zf5W4lCo7uNkcpfrKcVs727GQSYMKyPya+RpvLuhDy6H
BkezBqb7yx6dYCyO7DJkX/A7bD60BVeAuhDA7TK9JOFS+9KjYMz3/jk2uzN7tJ1Vt8kmkPn9CiOi
zUXQ0Nc1+WuhDdwxwY0UcmajfoznM4QLMNkFkRwiHNsX4VFXZu79mYmpbkXsLtfTeAimumxZjhwl
/5c33/kJBJRqccerBGzLgDPyQzKGvvH4kqopIWkKc6GQkDZT0luXPJCl472bclm7N5wAullkmx9R
m9BHrgF0yB9hTsl1aGdRm4aiCTwbWuNtUfdZrhEa1Qy2qEpxLui59O7ii7+fF1Wh6v7H0KLf8EkZ
6C4F1i8LBstvgiFw9tYrzYXzEOw+/iDZPMOHNJVs17Xlds5AwgEp9I9yAfAv4aLcD+hCwEW85bqa
Kun6PsYi4QLCYkuHeRPKp4KVGZSIDWB28sdM/Qw26GrV7ekLRyiqwjgQYcSqcrBvK+Qwl2j3ubvt
sSjl7EAFWxAdf3pKi21/y2Te2UGNFxMonA+BKmw+VeYKxB4KoulNul9s9oNLIgiupSlS0YtwFuHD
x/tLb+DJJFRpCZKr9fKNOOGDGF/FT1JtYHx2HEg5QSqsVRd7cLq06n4/92VScRoWRTkdySdwzud0
nNtVKu6aUltFkdcs+HoVNGsbYfu/U5yHUWvSV2i5f6Ek1c6QF0eQ3hp49vf3i5266sd/blsonNOV
eRSiwZrak6AXlyuCD17UZcB1GS9IkZLPoITF6Pdqvd8Z0Kj1QIBebD1mE3sa9A1B6FQGHYsDQbi5
6G0WGq9eKtkt0mdW5riAbBRRQga9/3aaLSSONG32wuu3CD1ZKDfSUsQShgMboMH18NtcIGYF1+nu
rpzKqu0VMtjMWHOvATQOCN52YrA3TTrWf0JITKOMtW/tZcOQebaRYnWi4mrJCEkVqJdPNcd8YH8v
Z7sOVu/vreeZSO96VlqBY0seeGbZrdAKMFgQYZ7bnpmj7x3qknO+B5r8WSPL62NNs9mm3EZrvB1T
Glf2YKjWSuZqpJ0WdWLjAPtsOH4q4zMCjlQLo1/JcI9KaD6vURoHh9X7+XCdVveiNdYb5WivhbQP
SUMNuSSY/9+A9LhuJoKy4Cwf6r1aruk7xOlulqD84bne78WcfeRDRTdA221+41nhvVMgPVJ8ej5u
uscQsw4v+IOXPVeFlcCrt4/Sgzrp/3sI4i2KphJOCIyLzLSYX3ASRkzTlVsItIpm/ZCeXgbny5aw
ZVXviNLIsvs1fdBPnlSmo46uwEkQAAYyTqPXmxCMTYsdDLTK+WwbY/aHbwjhs4wTJ5Qmhak6gDwg
A8fwEpnAN+TOofqkN1W0ipe/lJFFJDvWKuYMd4NH0jeZXgcMzc+FMhXyT5vNRkkanPO6QYw8Lzqp
0OytHkJLANTaVO83Le6WIcQ1jFSSIafVd79kdepNWO0jSPcQa1gyA47/aNIE8Xvuj93j97npuRdb
lfgIwvScKgNyr8PNmhcvV/Mw1FcD0rP2+lV1YRkmxhgYyZQbdtIGH+mDr9RWi1HyGTDXladlo5dk
gGME/kVM69B0mF4eUx8EYWHvYt5hUWI+p8aoFSD2W3f57Ti+UxBPL1eyYvfGhUUKTLw+nxLeoTaI
1IIFMGaCnIxDat13TQCBofFdE+ECKu9YMCbDDUPLRZftxHSdLPAk9ZVqfjmia61vPsKhZayBdTmL
muwEiRcgNlWMJXZkAOaUpgBHzYju7ti1Azkf5t+OmR188F7VG3Dnq3x6d6TI36WuNzJOq6AB2F0i
suZZ76mPqxtbfhfjMV3SRNKw5cXnXn/DZ7mdZKNj0qXusTa8NNUrwQpWkpqMz1ptaoyNjYD12Uus
IMSTLa8Q9QV7BeEjqe+syV2BbHo6oI/HoGpBUqN3KfZkFimD9dzB3aitbhADz9RR8+01ndvNsLnj
H6imM+LdDn6U7PMbpN3My1tscv7u5gM1nTJ28AekCNc8w9cvr+L69rbvWo0TyQKN3OFS+VH2LtiY
g9zvjt0mwzkGZMPOJa4lUFEMSudXwgJ14l2hFvcez15/5hoVBybfOi5liDb6Ll/w4DRN0mwjmokW
IwzViebX0jNwvDVvOXK4Gw8A/35X4Dn86P0ec3VUHWm7Bzrm53J3je3evHukq/UQw51Zj8VIo98Y
cZ/TfvvR58zV5Bq5HKvFDcGRtUg1Q8AkI/bzGk/Vyr89ltL8mHmCeGUVcB+KQ+hrXvUEZdEg+Oaq
qqSeJo/a6exHLKoWuS6ANITxgrlJjcc22FWdki9RyqZuwE4nCyvmSJfQtb2ixzwjOX8iYdzSCut1
sDMLyvaokCqjrSOEKX/rMpILTPt28qV6w8llnUtreMXlN1yOQHugtQoSJpY+faIAnIWsPikBcGiF
cL2Wpz8FAmJdLL9rji930MZ/9u7T2aUG7feYjKw7X0r5Y6iYS2ooxoQ7ntWjZgbzvHHtoX1fI6/B
79ibaaY1JJQTlx3Vc4ruEw+tyK75Ky/xI5SxeYYJom9DniMVyb9fy8tJOn9QQ1Obqf9L3ugxO0Qb
lpN7CvMur2qOzVu2EXJhU48JpCx+r8Nz3+1xMLj8sw7SStHuxotDRueVW4YvQcPzSPaokl6K2Tzg
U0vLJOBtnpaF1hcoL6oOJ7LijC5kux0CsfTcBvVGt540BTEmKMz6hxLorF332CXpBV2BqlwJiI4o
jb9gWKj9C3V3b4qTaF/5SNL61Hk/ia1nSTRtHKdMPRWrD9HyfSl8xlOPRJSl7MGUCqWnFWC0tlmT
XRko7twqRQmhEcsbJMiYGtnw61V6QIIvCd5rfx6AA4pgLF2mLb6UibgD0r1Ndk970G6+I7a+fGgJ
xYiwsSIYbK1kEtc0cRgoD/07RLrSo1Y0YGtdYWlv04GTBNJ1XOBI6aYfPzqnphbBvmnNX6WH6/2s
XM3bVasfMBjzOkq5E4NnxbUbYW0a7o4JzQLLEFCvgUXFQN+CUzVZsTqUxZ9pfiNy/gb/TV15+s1J
SxWvEa4WW7RndKc7AVxDEtv6jK6QInCp3y8KSC8CvsjckF0WYPLh3G6iXA1Xqi61aDDdM8TuGYqX
070Eyok7Ped2ob//ZYzvg8+2cbRhHJ21DZM+8J/wvp44zUiDDaXMqJJuBzBgoZsBCyTaVJTDRrFv
e+IxiZIhw4qZLqMr7qTzhN7uZrAQs9dNh0Iup8Wa059TcwOWI5xObiaaTxQrroF42EaduPWluqwe
eAKjP+Syh3WBxbTo61bRRUwoEDl+Kqvh6x4LluEwWWi1dVc3fV9WhDPxq1uv3EnXfS3c/NSZfp6U
bZgrHM+JGTE0Or/uTa3+vdiUShxyk4WhZLDx8dfX26qhdxZ+Mi725AeFVT6guQpFjuJ5Ep4fZq6j
IXEDQDfLy5YiVCMl1NPYlXvVCFpFqvFEG7GcIpJaVfpQ2ql5Atl/nApt/gdqrk9T60gHqPWDCwte
I2tHg8eDqWPJZTwIw4TJK9LdkBFDKitlSWXoEUhs/iiQdRhU4kqd3v7KKw5NjkqM4NwEMxEqnq1x
WA6I/yZeWkyIDgjDaNKJhUktdJT9bfkr293B8fj3UQsBJWoydm8uVIhCh4uuP8KE0+vuxcmJCmgB
kUU9ibHV3LxsBhNVit/nAUyt71ONGrq7IcdcS9fw0hOhj0nU9y7zzhiibvWX8iF4qG1AK/kyDs2M
7X9f4lguJsqrJRKzBLO/avxoK9hV2ueSKsBGW5uHKTzwJM3Qghtx2zlsPtrHmoKOYsnym/uhA8f4
k5OWP4GIKTthDZNmBSwT4D9BawF9EsG2BjT9YvUQl34wBlDHsVh6fBpvcVGhLyhrxKffz5a1vCfM
J4oA94v9cUXcbZscx0HcVAxRafazKEh7OFhOuujGGuq+1X2e+Y2XKH0tee6T8xINWx8+2DvARk+y
phUgE3F5ekqGhu8d7Twr8XUzg4wiPONs79qeWrureFwpWQm2PFLGhRLFbsmfNbrMtSJ5sfNyl3Nt
MQAddr7C4M8DDiUoURJhCQOH9mN7CSAPxN4YSWptQw+n5tgG+5yJwzJRSYODoigh1hdy8S8ZgTOz
vCoasDCsdeOH/35g52AnfbpUfpQvgVGvvSLLsIKnj1eXhoS6LjPIuFcaW8fJ2aiB3ES/cDdGcUN9
lcCUEFDXqBKPB81kw2ygnl0QoZUA/qQYGKBhjkBUEKjxFdBiMDJ2LPuYTU+7vknjiqcq+wiHnAlB
rpHXQzYZvubjWl6mtyNw+1+5mEXneYFPuQsE+XiE6zDJ7yf+WnR/CFzL1pqUMBZj8MbzJ8DmSZsJ
HuK6aGSSppsQQFZejxkuHDnIjz5YyhJN00A25kyOzxU8BjZKd+c0ptUgE+rMmZYMcGTKsNCJZ1od
kvH0xsM6qARG00lq5F1wktVt35fhiqUE0mKXBbB4aZ4JD5l1tMvWFcJ7YL/9O4+utTZ+NdU3TiJ/
180L0N7E28eU/wDcb7h0BToq/rAlkY1q+2/EIOsBrdPYumzLy9cllyvE2Bh3QrfhOPVe+t2ZzeNR
tHCXF2vadqcTgg4nslJ1YAEPwJ6INMs/jIVE56h3LmpSczMkxMqa5k82nXDwojcj24AGMRTySH9q
P2UVTtCruv4OUIPdv2ohvrJ7EiGeZp2puH8ulaUKx50njFihQPrcEfiVDbIGMzlsXiOHJbVRAvlr
GnrpPVMXNor7l9gAf5juE+CGC0CV81UIES8xsCJ6Nj65bRoqeO3tTKbu3ZPip0qA0Rnc3dUqJxi6
HcJOh9uPsrx72s3BnbcIqMohFGfoQXSjWJaV6GHjhK8QHRH9Fb/37pKPBZEdLft3sSwKSjiqz193
fIJ83kyHEvlF6pN2yAradxR68NTkrU8SutfQ7quuXLlensHJ2nITgStv0J2z6HWvxAKOOWVyHalc
YgFlnMzxTC3GhMnNXNbtFTG9Sl98c98TtAqX7h15M3ASRXGhl+lv25nVYKCLfB/J44o9nWJGtnBM
2TOePRLvzzCL8n/yRlfHoJ983ZIUsvWsQQ9Or9WOcQIPyAIXbxBCqZObRXgJaZwhk6+O+aZ0PWst
Ws0fju4UA/n3AMFUr9/R4LxX591rzuKQM4bMPURoUAsYlHvqTNuMS5mM+++OmUWxmvWbWK/06XIq
9u7HmkrpEB7PnLsFsa6S/xkfPjDPfgIDeWAjnOzgj/STVUXF3TXusdigSqLfFPz4wh4pOhsJt1rX
oDJayRP4cadxyZ1txGLK7ddE67dFmoCRw/dg0NQjFFXS6P992n/ftQaZKptCuS/YQABedpTN7IHH
ntsjTX9QObPhZU6J59EfRTCI7yvzLi6U+kAw1JRpaOxZvtY4PTPI+ND8RCp3aIwGl6Up7WejOidr
gCXQcc3RZ+/X2s9HxTsQG63fNTmU5HuOhUn9uLFqC4QDXqzsZAhfesGthYXMGRu1Vu5ao+4PYr/6
nunag5Tu5p4v9R7wQAOzbS5bmsF1H9M6jJyuIBGBpRhLFhmdCAD4ea8GIwAVIAkBiKSp48Kj4YhL
EtS9xC3DPachvTVnGHsN6LIMMGiqH40DXfyMeRpdE5ZZcsZKfeS0piqRmZRa4d633zbH06JNQnr4
yaByQICjfIfIYeiK05zKN+5W6/UjbptU3uqXDwW4F3EN4thmHgP5cYKe7wx2UewY+LkpjKTzegWa
2QvbsRRR90lddlf72scnpuzng5VnX1GRKrJfGwsJvW2J+TlAsuNvss1wWWSf2P/mX9mf5Po46r96
zpnprfSeFRJ9lGB5/ke64qZ/bugGWKmDi+pBTIFrqxunztF7W/z6xnXkXd4EMdkZ4DSlsSBHecRe
SBu9I3AEuI/DqX84gVpGB8LdknF7zcPUbS85pcm18lIsTbgikcB8bUoJJYLgO+nMgwXqZ1yoysTg
SARnop5xlKyxbnTh2bZQSP6Sf6WkCXv8Pf3AfGubag33Aw4h5cv8Gn8+tL2uKI3c6HkIgVp/Ymei
9xj6CWMWQN6zQNmtadIJRnFUQ1ns4CFRym0xwp3Geua4XLAXZWonN/qbZhCHyOohSipyN6I7PXEX
z1kxp1ouwzDnlQ15d9kAGkE+Lmipcma4UHUvyPPStuk+UEpg0eaoFnhwm04oylawwnL66g0ydRGq
VXp9vdbC8bzU1Ti9pHS/PgAFhdd+LbQTaJeJuKM3yLgyjZ/G8ZvgrtREc/Z+1IIaiJeKU4A3F1bX
cOtEzsKiUFb/ewMU9yTqMyNBfYfRUwiHJ0n9OoYuZwLnt1wNo0l3juSx+iTn1ojEpKw+tSr1Cb6/
Wzq6XlowFY2m34XYeIGynQelKijPlB4U0jMHrEXy2uxyAXXJYi3JKLjz2sC3o9TS4Q1esl8buqNB
5fLTHnpc6pf2H+cC35/qCrYO+tLUSRDN9vM/IUEsCQr7lLGBSzV+zd6Ihrt5s0xwlbFxx3jb0Z+5
3YSgilEq/1AT841fEHGXjx0qFSt4br9OHekWpR6lH4+Wrggi4S5mJMV/ZirI0jqN/uDjadtsFy1Z
5tCJFSpby7TdglJPsoEHoZJ50VRNPYcaiI28AQkSf83y2SaCsAuRl7OwS3puEPo7CEKP3FhJzzn3
72bqKAHXrTVGq+oqsCYAaGQnOV5AeWQRKPls+q8MyFIx6zzRP/ApAvNaxJb99W3nP7eNA0cjrKcp
d6+87JHbJmV1zBPzAUqrjETExNn16iP+VKrGd/xCb/2lCh/615/g1G1rmHURuy22B7ZrDuYiskpm
6gyhg1I4/LKTPPEfAsoyAwrc76hXBk6gxWn6iyAdxUK0f6mPOrfSLrr6iticoJiDQdExDYFeumRK
l/0dW9X3ffYzFxNHx6SE6RUQIeP1krbA/DpSyr9+Yz5Uhrs8vBWmQGzdW/PbK08pcLs+Ild+mRAQ
6N5uipl6Nx3nHFD2IdCcFmiYpuXDZcibVNNkxTXjMqG+m1lBhhKYLa2j+S1ntnWrHjiyBBxTCa37
T1MvQkuU7oM2Oug4NlhzqcjXBXinXOnezVI+0pfg/W9ySywaesU1WEg3td9uEFynq2aaj+gyvElq
1R7hCfOV1EkJk4XZQztTmLBsjkp0uvvchJv2HEbQ8U/SlRvgqaOzeZ4JePkV77v7cX4vpCaX5LSd
eHQBFdvWv5WMXRnkd5DOxRPkMRasWnUH7zcODc3AKtC6rUx5zl8izycB29ZCyHeWfcV6H/vEVsWS
hCDgqt1cI8njybD1e36hNHgFMtFNaV5rDoZAuMRJL8K98uuuqZwIu6lSAgrcR8X2nlSrmp1M3JKi
IMwkSt6VNjc3E/z4cUsthtJXVHv8oMbXfPLsl2lwXKKdxyxD5/+PXCF9a0D3jMWacKmIgN++Jo1N
FEYtsIPmrfepeDbC9tYLSXVCpN6e/YEUiBSEI661demu4uYiuaeeEAF1+Vm68YaluDFRc8VuPSm8
DfcTsDOX037d6vhS0lr6wUuD0N27I9XLuvLvMBDi+kEf9ICP4sal2MwYXSrSJ5w9CTSqRsQQBwUV
156alaQKyZV15kADwuVqOKl+lPzAl1mefRHgu3TwWc3irsf3umtxpcsoEl5ZksP4YD2ed7/9EtAe
i3H+oLdryB2wUbe0y3sG140CNvb/RInWUTtnrF19nxvdk2I/7Aubcx2THCq9fXlAqZa8hw28FWz6
WsVeDU6fXY8PBCSF96rosEKXLmXVwUaFKHJ1u8n5qMitexG5oMrDEhSeGplWaBXb3g+nxvwi983t
Y3yg8fY4vzgNqd5kNppui4xdJYI06J1cPA3KNlkhVC4/AL42okcOEbuZuQm8n81oqmT3RdfHCPt9
N9sE2ThlxmgQVnNDo9QKcR27ZCRXk1MiDlrwFh8IAnhaKE4b840eWj9M7r3evxXRCJSxa6rKToL0
llwXma4TXe+6wf7RTa9euHyz5TT8Pb6iy1efbf19BJ2PtpYV/kTUK2z/g819RuAZkxlzQPXxRm3A
2W7ApIVUuiar/UTt5NYie1s9Z2T8lumOhOqKcuBzpevkQ8C75f4xwNO2ShFfAgY8HLSv+i2b7Xse
rowOvpAfsMRQwLalKpG1vAh2F50fpUp4VWV2KPyzx32Sio+R4wZZVh/CsoC/Qd9WWuNsLiZb/P69
XnsDhCNN3KMG9UkBtBoe8pr/5yjcQssB3OZgIW8UNK0DDZZh7US6W84p+yRzbIzW4QIMzmPpz6nc
QFx5YJCet3gCmtgr3Pddeuy0SijG+Dwmk3c2Yz1jgjYLagT0etqDjkesnK/43y8/uRukmXgaRZNS
gzpYUQ7dGmMR7HPflO9Xg/0x5OCCddvX/knGhs1Uobbk5Yi4byli35OfTdsoO+gKdJkKJPr1vtTu
zXYe2edo5jiKoawrIZxMxgC6u5km8aC6SJTqNauA3g4hTNwXQe1bY1TShdNf3d/FTvrC1+qUdI5P
zzFSXhDe0s6QTq1xiAeHvqsGejOcte9ScNxZaUam/OZldsWLP6ndZQhQQMW+3Y8XysHwzyR9oElC
6MhCCrIXaCz55MQWVQ33F2ykcO/LS8a0b3bgxhqh0vQP9X5eWqOxzAFR56q3dP4bp6JaDa6ausWZ
GhKtyOh9S/xOAwRoUrywey+WXbQsXwDKitOPZ4PkO8OyU8rrrQ2b2uLRJl/rHbg7AHYYbvEKJs4L
Xy/xe79Kf8AoLNZGpL3cF3iXh+xeurQq6HPAxDgAVoEGggj4yFD0/3w753u1z7xQLIVmp0QaqXGb
Wy3qBKm8DIGIPM7onyyyxQEtgHVH1a9bmEcqLijnKEEm0uyj0PyF3HKGplRKxz2ORJ9fcCPjp5ii
VWxRmNNwyXLyaGA7rKJQBbiiB8sNRwIvsv6tPsP5w17LbqY+fH3wxQP0B+613BWpbpCuz1KQMgmh
+Xyg8sbHNahGjEyGqgQiRwuB8gxIXi7/yhVCm72sUOJTfToIekd5ihr3Zbaa34YOJfDdUghccLqz
yMjr4YZVR9xgvIsu9fgryXdKyJDjCEiH2JOOcPS+PNCFBtLEU+iPUGTm1sx1se+CZqu7MHnVhuWF
FSlil3Whv1BUz3HmCC9H1NgCrTv4SriYplQrukRs7ScDcBvocLZuHFEq2hl4Mwlyf7uWsJwFc+Vx
cKt/LHmiEfwXkIjflanLQ+V1kPDis+OjCEPNL/cPV+FAlialNJ94Ip+IUH2AyuOgeVIqrgrEwcXR
7CHbTUOQwz9KeghfKMVVGg3Z7IL9wTRqRIckiJ5RVlzF+k8Urte+jR8vP8C+8SzQMdptBtmiAaus
Fay3zq1ZixxqHplfTNJY3wDgHNMZNZiBVJ/cTjFdZUihwuc2hHj2jHTIK8Dw+q/OI3iFzZPJN7R0
I6RGjFrlNu4uuOwXqtpD/4zruRVE9yh/H/c6TLw+olmi6qpBA6UXJngtzjtjSrhYjZoe/5DSkD7b
DGKqYlA9QwF13Noz/LpecBHenylwfTD/wSUq/q7jUKu/EYghHWp1Td+KYkSwS4enPKvlTPp3CLW1
eLm1w/xf71Lno/QHMfaVbOqNF3VAPec+ZTtAx/P32g/K7GZoYVpZ3/xSmY2s/qqmIKInwqkTgsgR
1rAmC6PEgjfUa/HC7Pzc1eAe7XNxa2Sc+MFq+Nk9OBt1cyoIiKzht+hX+bQ8UnvPRd1Eg1WUuKzt
eFd6utKOn1kU1TVxoKfAlFxGtdBl94adGYp6Y8IgI7Ia5M5f4qtBkPhVHgPgCJ75EjGhzSWELQVr
0VuZWkLyXTrunMABG6HJLZz3Ai/PWk/h9/V2e4nDGP7FNcTmmNYVhGrh9PTqIxM+20Ff4ILBlYK7
A/G97gofVMsZM4esz9AFL0XdA0ElO/oeGHbCveYtijU2KVkg3LjQWrhcrbgRfpyFP7TlSm222+/h
HwASFb3kDKe9hhZFOdDq//CWGFga2hqm2E8XItFHv83NB+mk0B+TqgpzxUmf8iL5TxsfEnKAEG2n
M0X6alr9OtrYSwi2Mfo5ZUtlGA0ZCF4vzSswL1fBMUnHIzu2+GImQRKXkxjT8HGQ3thyYIkYd8lT
7M+x11VL8HYhdnvsV7c8wUw+6uYcQUkNMwm2OO94BQ/p7wnQMPGviQl1xqQdCIStulX89jYq97r2
uBbncp6dRsCVnbe5adibJoAav1fwP4PHDNk5Jo5Beuw4jkEmCwkxw0S96HUCogCwlEBry3o3U280
aEXIJQEc0TicJnHUM3aJmaQ83Ofdw6INuq09zvLdP/340HQJA0sv7keWHIUm0KcBQOTHLOqz0BRY
bd0F99tlf0Gekd8Mm+EoQXK2bqhxtTiHTgDmuW8Yz1JSLZdRcwhFADQ1gdessxU9eOp94T1lyQ2C
G/YLoEZFLb8nFFIYhQ9wnwS23Nbb2u/imm+1nimod8KemRNQhhSVPmgPRbnd9SA7/NEyHz/na9ua
JCf2ThEGiCs+RmxnsRQzbsCCwmS9DDSHNhIWBCbsn/6DC1ZW8bXkLVX9B0/EvnVSoyjZUBDWie6S
onCJZYH7LvhFiW1eyT9dROxnj37wXnRlLA6qbpKZFCsUMTXX6ihMRO4rpHusDFy3n1uyOc4npS4b
KwoFEJ9EyaeajE6BzaJp1Op8HzBXOsHRpiG4wLab1RK5fxJktardlE9g7jg10O8mIrH1nf8iA3jz
OWLM5bLe99FrKyQtStMOqaIBNH8PggoJ8vFnyQ0I+urIvMbc2MMKFo/UlkgVKSi6inddWUYjG2GB
L6j4emWAuGABiOxdwcHVorJuA4wItKVUsDDJ1aZbkQlEZoipks2uTCSK1VzVVD2AmDVxN+7L2zTV
C51l9ac/44i4BDCqRy2e7pk81SbStKsbQNPzrJze/52Sm/0r81GTNVyiy2BinZLAvhczUgQ0U+Vs
vVlrGQ/qqnIV6ohADnZ4f3pWBzSeCeF6HkgzbE43++26v80XveqW60Qe4/cREwdv+kuxkYui6hlt
125C8EMR5a2suD9gK9yOdOCazXjJd+e2Gr9kf7RIDislBwxIJwjFKV1y0qYv7yFrktriBKmtc/p4
i8C52Z3QfBJhkMCsXmQ24fBp91xkqruvmGNrgyaTuKg0ZyJ7I4unY28Y0QdRmBQXNwWv94qqO0dY
7RGzPbddXxA2z/nF/WaeSWW4enwP1ZIPiv50aiA3KrgEDG5BU8ItBJu5fBGAYUKpQHZB5jUyDbAv
jxyL7/QhsAJCDJZoupCZYd92QcqKrAhSM62fH3cE2wR9ijLMq++yklrJd6cvyBPTWGmD8zblzmAx
g8tuUeU5QZz+qHgtwDjnY5aKsjUV6nY1IO7J6mowBNemHJszLsmntdGX+lPd607yVUPi6aXj29Px
nMcUeJOcVo3t+JnPCpqxCtQi7DD2M6x0rPJzrTb0YGyLyIbbf9D++T8/nPMoPlKKsZTeiEchRC7f
KlN9O4h1YwWGR7+6yGeTkUeotO8b0V14fNlUDmeIz+PKCFeySBFIghemceXHOHMS6zzPFx20Lr2e
/ag5s/jniVLngXffsjaRYCIfCwnmzEcxOGCLO1WE6AYzQx9nRU5MfITB5VuH/iimd+iEznh8g7ud
6xZ1GnCysItoCkNc+ADo1XAm2jWUOz/mwqMr5rm0occmzfCdlvnHt03/+g18y6ZX5ySSxAuPSPtR
SQMTZeodRuoANWCiE93Y8zha0i7aspBZ+WlIwAZ46USVi80faYMGRD7j6oxYAkBF8qXmpYEABJxB
gMevpBa3LjemXnLOJVrGvDeVG/ipBdkGg8qiaPnInL5KZbrRaDo4zpPd95F0gNSHygiN6zJTIdyl
+ZB0r9Wdtb3qj3nJFGFgC/wpIccA0hwKr9y1YQxe051zoDKK96qNJn0vBewkpVNdnfbN+6cdaY4a
pB67UarfjgrXL17iPM89TJOqS7WM9dnMWJWeHYSGaKE4uzi145ByWREYcIjObuZhgdFqOELw0/RB
hGL1f768hHmd1zfpM+Viljcc71gY7UjjdK9JrUrIIJ9aWD1hu/m55WLj8aI5LQ0Qc/nWsBoklMq4
n+rgFtvpSlp99PNJA2S+SXsOLyPrKOCvifLGuj2WLE/hZtcBJZBs68v2znNuFW89BLmesXGzNMl8
S80y5/WzAC8QOmygF4qpjKVWcWFghM4uzTjuMtrbwiABdLZ5JoSFYBXl1jX9Phq8mj1EeoexcUHg
XeTVJa4boQbf3czH/AAT5xCIYXZPe8Hy3xs/hVSDfu0f3/cb6tAh9Amf4PfuCDT0qlxlPWfq0vNZ
Jm904wgwPQpoj38B/V8BPq4yi/UcW81wUBGkzdKkScI9imPUk7ucg3zrYa06YSbCb/X11Dwstxvf
/YzUhRsyU56MEZZZpBKyeSc3+QFb/oMtXAMCyLej+xAS4R+dRYEACw4h5udCXrDMjN459Lau6RqL
pvmHC1C5bGv9hyDuzQy27v4YrNojDP/uUkTyLZXaw9gpV4RGwxJ7QmOcH5mrPpjpuBE0r9KNhstx
AYJNiz7Xi5MJ17tftPmzl2W0+0kX360ZZg+y9WomFbJE7jrvoPV36uGFGfUnbUHUkZXbs10FMlgb
A8RwAsU0+uBKDnMtIbCTJnAqoUu1z6GMnAycBqhuY3xkJkwnYwAQNKg6ND5rKP37O1RNWUyKw5FM
81QrEvdpcvyF8H1rVUPHEa+TLsa5dovlBfT9bPvJF67MaUapVrynueVIcua3e3FGpLVjOKRNl80U
ax1Xyfu+ISbAk8/xU2PSyqq6bfvVQ4qL8cFpMD910hUQfQoI6aIiDa8wx09BWx3KQUEc79s+tyIF
ie6Nau/rTa29qTCWkdzW8QciFRjjf8B67g8PmQnQJ4Q/SLWMx+xfHJ+YY1jMxBc+5wrb59rNSink
NleIw91BX0WiHPJgo69CnZ9/hvvij/b0S/isJgMN5AUJJ+bE9+1QCUt2Ez7BXOevhggT3AMlrlB8
dZgE+HQpwGbAzeWqtcaz/ghPYSRNgL0uWwlSgyV923QiyQe9WIha9r9rsd2hJUKiNFFLE+Y/B0hD
rz93KPZXfH6ukqPNu9ND32mrB3A0XNUOjBU4ztH5giFpV5ok5TK3blNwQDhvvZ6n5hsvM4Yf3wGU
kKhQVYf0ISQ5V0JYhUCR+MJ5XwHu/j42DGb5EX9o3sxiK0316NIet7E8FyOtTkD/FeMU4SPAHG1X
l0Ne6x2HoS1/OWCZSoV3EXF9ZNI1QGLpXH1cXWofXb3H28jCywIKciE8Pc+pOJO+d8KHEtajECXj
ty4LFe3aSQWK8K1JC5MYyZxoa1Joa7Bi54yujviPbEHJ/5rDzMWb1CQayhOcpaiCn31umOdVlMn6
YU8mcWw27sCtPnQEMHk6Hn8U3xLrX+cf4adEtUIvKw2X/zuPLeVqNBsYIDRkIV4k6lpVb4LoO5px
rV4igKHv1/C1AZHmrPkawZT4eJm129HuLT+D5R1C168GL7jy2jiA2SZd5N+J/uFuNyh11mE87Jsz
b7gjwKHBwI8zuT4ePNC4BlmA3iEvuEUEtaujBy9YiOWGpHbtB7tRjCPq63z4DCmk4IyPDPSH9B8b
u7V00C7Qpvdx+2s7oqmJdgWYA5+hZTO5QLYTrf4vd/apD5jW6eFeeQkUrbZ57POPQ/7RmHtHrx08
lWwf8QXMyYNB+tNeLMPmVCW3DduR0fozqzNjw27whUuQIYdDpfSxijLUUrj7+46rn+ZxWQeoqvR+
T2DnaV+kXlrEAy/vjoiu/gfOpgEetkFr8sayiS9JT8IUFT8Uu4YnZlhFTFbThabDjSwucyBsWrYE
zLI93sOEj2C3wtcKtwm6N6UxgYHKHlXGIn4ArSemRXN7A4n1o2BBnHNLiCzqPjjSoOO5MUnEVzs5
p/XqaFCPopgDuVApneB/0wLs1Zf7k6Al1Yv8JObJp7ykQARtH52zp8oAEcY2EGrGYr+c7qoVcSoR
4UQPtdqde2IwWd6PrNVntBsWYtaDMVUVQ/3Accaa0RN+3my1SipVXyX1+pkADezL6ZeNp/QYMWpT
Ell00v0ESMmNv3REJFuU1lJJYr0VqMED5FiFrY45QpQuNZ3nNnidrgrZpJ5xnPviGNR41JtZCY1m
VRmpoCI2QNgcP2JfaMfUznq8DMgHlKZmo8SzpAKXDK4Y3KlKK5MPVV4Ks4uiOmmdLidsWmTDtOH0
+p6YuX7L5LwVhHJFdKdGQvoFJZwdPMzvfz32k9Ft9tU10GipcbX3L9mR9gsBcJnxkzdzxujUIDzw
q07/WCRRLj9OHIsYGeE4DJekjoJ9z3ILhSst5gDXaBQWpitVM+g5hGAzp3VBkhl/tUnUBK5CXH6X
9WQieN8oWJFFep7hQYv4JUaKMGUtuPc9xTeEj0xdXFwOiFiY8nFibCtQQvf415xfW0DtI7mvgvF1
VJjPhcq3Zmxp1ivcXtf/ymnhjbXWpYiJTLxUoHVh3cazjv+9q04v+5v+FCLWNIuheQ/vdPRt7QZU
3sZTaah8AAAku37Uja0z81h0COY5kg5VvmvgObiPpBkuHRuI+PBz4TZDJE6Z4a/99QkRPvbE7MLk
J876PHgYyFAls3aGd4R4pgBe1sKLkCo0lAbvGHYQcc8XPtbO0fX5GNpce9motug//TpMbIWZLQyO
nH/q3jXC/yPMOtXEZkRch1hFfSAVHIKCTq4Sj78Eb3xElOe5yc98PYdMNC3hTwJ2tiuspHOZWPtf
jNotLBaHqqTJMb+cGKdZlxN+2z2aucOEyTDzWfdBhOZ5x0ibsfcOiHvWipug66RcMpLHkSCFWVEI
BmAmzMpvTTU4JF9qXnC+K3JsZ/qF1jU7DTmtx5P0i1iatmiGyELDotF4VPZ6ZuYuuuQfkqRuCxvO
cbTE3+HtNQSjOCZrfof2oeuIbBGp8u1kjjKZKZQnqtGw40ECK9OpQAouuabIy/lZ2n2vrR+H4xVp
wEu81TV0VshMWIWgFVGufYnsP2Qq505wO+E/Rw4cI9ChQyY1HPqyQ2wgFO79DIbz6nLK00jlxLCz
RoxTNKhSadY7UegUG1zA9nWX7smQQdgpzZNVxZ2Ih0ngtog2tp3fMrUUzzRVRRsyPzQ1DSZ7dHZ8
sL2LjQGOoTbGAGo2WnM4TNN11gnsF64sWS1v/JIfMuSpnAr/NXPGGY8xMZ9ESfmyNm+DACMuxr/w
crScc0UN/9YsDvAl8hpbzLYqzi6gOdHElcksJFitsi+XoJgmUJp2QAsuAe798zTL9624wTVseHjv
YNT7YGN3xnDoczdxZ/Nwi4zY4aOTqLeUcpvRllIxYFoYOBhuOBa7N8/ffVZ/V7PVofBcCNRvV8bM
pvSBoSBMcSzB7tzbM+UX6SHV7F38uTvagjoKJHzfNALJVWDmsaqDnzdNN56HeCkfaLG83OMxTYk1
M1i9j+w8Cv9DAN50i1eFwWYHnr5FYP4vxi76Pm0cGksDjUSYvEmCltKrh6DOK1pMy5qUz5LJliGY
VjGixQA2KyFFk/mXOqC6ydhM+OCBVCzHp1nKSY4U9iKackt04dn4qckbNtv6S7MNDY8m+/w4Nwcp
8NdFo+VXv+l0z55RoYayQmW9LJ2U3wyw79st+upGeHsqXgzem/Nn6YydyUS0S/yBfM4TfWls548U
ppR4an3apGXY/EOwgs6ay24kNOpkba0IFAiisvWWxiERIA1NsUz5yxHa1wmrfZCBeXNG2tlqdIo4
nY7WdbRUFnlAgpJz3wYLZ1hV7X17tsx3ZP5Rxn+PYQ/RdtKkOgbsl3jLvWZIFUhT5AaXroX+/W78
tui6juCwHEKY+K1AsRIUJDJRaykERuSBsXbBW1BJplZdMtlpwuZ8uXuvWenHmr8DRVMm3vkTOPoG
+kPZEfXZ5kUwklF+xQwEkXwufqupPY/iCqQniZ74i3vltWMSol0NuTAnI28lm5epZctEBP3LKT0R
P6PlTEFXgTwlajzchqKlF4RqrUg8w/7SdxHOKUoN4HzeQTcac2CdhQYQQ6rwq4OyfAO1MvvCsF4L
nrOnkHwlKeeHxevbLjJqDXWwMU0Ef5gtYL9Wcw4EieZZ+JMG1Mh9Aauvr6Lq8Ox/74KS+0VSN4Qr
g2lR+QQrYRpzKRtqeVyHauh003+ZZLraRGkuThvjjPfr+TkxcLo7qrYPIj34g4keM8JN6cvq1cUc
rUxHvsNSlT3z4wthtUoriH10Bo4soxwVV/4Qz+ft9OwdLhygDozycjj+jWkubZHgmMfZWeMpTCfk
Hlo6/f4IIAb9SdQuCqGXxK1cQ7G9DGrh5u4lBUMWxH2/Jxyx8Efn9ohzKIyeN+x4JhQEpED7VsN9
oZHP2bRYS7YfkkIb1gXJ9THR8sHJVmSpvJkEu30MwerMEQ3b8IyaL/PnRDNcuPr1HgYaSR4yp+Pl
4dVzcjZVRMFY3XD4/GKtstNfP/zTGSG9UHEpp74VD/7/HNDg7QIycUihlqZiPKQftMBAKiNhgmle
Z3JvKoDiJsY63UwIQeNFOF4LTJUCOrc752O0mW3WkbETp9f6Et6Tx1qUkKDk5vjWbnp6ORS0Kavh
ypVs6vOKQGVUpJFT16os8mZzgcMWDAyh0U72yDiR7bTsr0HJYClw7FYzwdoRqswhy8KcA7rcmCNw
RTJo0ay0oBxrK1LOWAb597OxWpho9zcn5HRUK1u3Uy0DLZ7Jz+W7Ff5PphHQwt0qQiQc2cu1JNlp
BXp/DajOSWtIgc5m/zMMf//olMVD4+B6po7H9QdlMSyE2JXcvvgNDqCZ41SD8dplG4RrECd08h90
6gAdRngvLplm8zokcO6boYQcXPR5uDuBNd4oJrpt+B22JwtXoQwO2ETQRqZ7zn7KkGInJi+m9hYx
cTOCiOkOUsQSkGPEu623l+0N72gvgl6zLL+lmqxIyCBP+9ehAyLk/+RYdKQ83LI3NgdYHyF2f4DH
5BwMTeRTbgdoF8WPe4v8C4zD/O0Jp0LG2yPb+bcyEmnxSKZAf3oVGUTTjZw1BzokM856VqOmHT1N
6EqXnDgbg13h6eH0clYByu17Z0wYFMAz0GnJs70vAQt7tI/OCWrJLxIJo8yQ6CTqnuCK8KMySuLG
zu6FpTPIa9ELgKYEEW8dV4yDnpcg18RFJRJQpkKOzeG9lJs0ywFGuX3IGcfH7utjTlUAHk4pFrbd
iTWF23MtrWjPWUwKWN2g4NfWmAW4GrLtEE/SbCw0xnAf/cbAzoFm3vYPbp4fBhFhi2MguvAAx5lT
vSDnL5Ks+oHCPLvyTkAKA11KpdyzjNrDW5fpo6v6BCeO1I0ukNRF/nyenG1LCDmQdKCa5+tS1Z96
uD1WgC7wGTlo2d+zg4MRDxlaEsi3ovr3JAuVhvqExnygxOTKLGoa2Hy3Td1WpGWVba6Dbl6muE85
LbLHZlA2vBIOhCXDM/A01C9KMnBNbAMQLQn22HGkSzMbDfK3MzoehHUeT11PGSiE/gear563vZv4
jvmJrd44uPiAqDy3Y/3lKO2AM0SqnYhF0WCGreHpVglbPz88P1qmMsF2Q6jbJO8nueHaiP/PHjMR
DUhQ1LhNW1m1egSHTEjz9Na+iWsG5vOtmZZHUniu19xMLqH6VVsP73+RdwD4DethKD/DgHrhH8lc
LAKyQFy/3wp0xOtVz1WHpfqNjauLFvpH712TNhJJnnIv8w3LUrQvO8Uix0WtDQotGALCjsspMpV3
YYyS8Tl4wQtf+WMZ3tHIbq8225RiC5qlJk98EJcN/E2sLq1rqqH2GB1HUmX9xAlM/yV27UyBOX5s
l/cbU2UduTs4GdVf08xmAeOMCpAZANhf+8jDm7jKn+ZjzZUUlYjyYM/w3w1ekF4KP0yo9GY8s7fZ
q2M75t+wYaPQtItkx6vxZBfPzWG6Ed5/oymil2APOjLYFPAYQiKazjTZadPGULiqFrD9pOcxnosr
aDH/WDiZfNrzOqZLSKmjctLVqbW5Al0nilozIkEbnHOxT0498l6QXFYDIFGqd7B47fuGxjLTzV6q
rn8op00yXYURcY8KSNiXjWsAbqDQ9qXPILN+vOmapCcc4egWXh5K4WHtaQ/jNQ4emXcjTdfWCITv
EtESVZPsU+Ex/6uzhLW7UvyaIGxx+n7ZUFj47750tW4C/GduX0/pnSKa7Y65vEb/TTBbSWRgWwQr
Atg5LQY+gLb6lwCWMeUeD8ijQC98jnkdr1PhzWoCE5z7ovRi4Z1KNKX3SvDbWPm5qMJbneR6gcVo
0Ch0WAO+SGpXwFu0s+WeKt3hIQgTiIbcE0EtF8YPe75vI4KmQhEfTEWCcoLtXtxpxDaWZgYyfkrU
Tkx6bbUNMwk/e+QrNsAc/+BWn0hMwZYsuypiJsfZeXzcaUZdAY1dm2dnedcP2ig7JX17YNUsDyBu
qEfk8GAS8CVjfqsiI3o8fiow9s1gKMqYsMeicx2WY13X/XyRSlvfRFdOXiJ1EDCW41c+fGrcqdFc
O0douzM+xS16s3ye3O6sQ7Vf1Bc5T3AsXknXGq38gk0alDtPnOJQzpIWiHf/KaDUagxvnQHd09Zs
6yXjMCOuDDOBTNUscw/Q51z1+wJnvshIaKsinkhF92HijHe/O2awy7t9HFs4NlT0keDKpCnFD1bT
X1n1C7gdTSmYwMRAveiljQgo9KriCKdM6LQJXBpChAR/inOnndVHw2YAn4K0sWlw6/8GdJj24lC+
mF1Qo6FtXdWiduNBAtIhAmbCOCYux35fPkD31Xc3fX2AnJHjyzRIowh3cz8RcZvaeuUtuMEwmVd5
O0kJdWU5qopR5elKNSTPoQMqI/yy9kRFClkfNy0OW7jRxBfk7byM1j1avgWpJaP4/SG+Z9tmbj+K
V2urkfSEkFjTiTCay9yKIoQcM0lBXrJU97LLrz0Z4fBGc+XUvu+t5IQ4LlOvZF0GQJHbBNJXU9lL
PG8Jwn+pD7O5PcrjyQDEm3oT/AQm4Tfr/3ayFgCG4UEG8r8vRvRfQR5pmPT7NPtvR6uDcoLSHPS3
DzqFYG8cDEdMj2ClubpNi0QsrDFIw5xbxLgDPT16f304YM0eHwxDkt+FiryfbVE2mpXUtYanKaqS
85OOImkkvT98E90vq8EB5rn1pgEFQqiuw/OzXAk+oJsVcCaiehSEwUc/rg6i8dqL44KISvoH8z69
edDMJQ3TFlbRjqR+j47wsdSc0udCIaIbObOTGvJ6uUy+kso2DGUdPJrU2LgsqFepy+cGfsqnNUyv
7K79wr6N18N3ngTJGScAY9XG89GFVKvjkL9AoSr48n715EZtm0W0n4LDcQCGeCnvk4qotTGbhY3X
cSp+kyfN2HIEaFggLwDjsjFd1oZQjsOYBv1O6QyqA1UvK1sT10eQ1GQFm9DmHGTwEAYNlpUBEiYn
KgfGx2LJOHJiTzd2pHGZ2YNMWGtcVOBV2hXfKTXRFH7Ku4MPZnkPBT4Ruo/npeP8FOAmRhFvh7VO
7jX0K0iJHamNSPsWmFbLIQq1xmIgPSC2k5Xan6i2BuADA+jxWph/QbHrWmN6glMYhETz1dzloduj
HjhVOaaB0N2lBYlwoGBrI43+2eTD2o38C7T10YzxD0uunVlZZWuJxPXyKzqUI5tebMKH4AKKfRky
ZkkP5azbPCYgL57oEcsYioA777zleN5EoGmyfuuDa99BR13NMg1e7oUmFTwcJDpWeAMDkbZSt5tV
CPW29eTklgsOCu/XXayWAczadBc8zH7q7yDjO9H/NeY6aaA7d5ArmM0NGpKpYGoKxEDnxxjTTEUo
G1KBKqAYNwQoKaMH0XRI11aJaespeN4c0ZDhCIU02LfSCa50EPzsQhQ4g8JkDnViLEhOxYVNVWua
KwtHFiaANolp1bXScc1yLAlDNwsVHvzsPQQ/sxqo2vBNXXAfcFqJFwJFUHrh7HcRdpjGlnv4DkxC
BnykU1utoXsPeAm6FPKvZLBNlH5A5JByLPjsf+AHRuKOU4OBFZCmmFHyl3CnGp5aN+VcU9K0QlQ9
U9DicZWFynJ0+b49XckUB0CBbEfpo38ggETkLMAoGl1mlQOQHgTMkpqSsguswlsY+Og0Vb+mPJsn
SU5/UdOe89Q7vhe/rqO/iGl/0zDWYvB9ZJYXPeNNQaHw5GDZ1dBrSxDeFc5KSS0mcQQ2IwZJvvTw
mdu353GaCuwaMhke1s1jYqoHl0KAly8stxGlmHHh6heG9W1h8nfMH++gWhAvQU6IJwMFFrcjUgR7
nj7/l0Z4eITMpbSk1WxP6LH9BvmF+FH9XSG0K4xaZhBtRNnqULzZPk//rajAdfB6lLkGS2n3mKEO
8Fnd0rYQ1ktDoUIga2URJ3SW5oQQrrO4nhcJr1wbY8iFxMsjSL+nG3qAMw2fiZv0xdUw6ZuzvvF/
BtbcvRsCHVjX13tAEf42cevoVRUnN4u9gVVd4Q9m6/7TiRohnM+8VAojxRD122orGcdmfIAXQbfu
NNzAwtUdBDoac2pRZtZRNAfEMAPkr/+GOlNKj7IcyDdBivcIAo8o5hh559lJrNZJziBnc23y2Jes
NBOb/aFTIBs065kPv8ywZdfSaF9vLJaxC/IhaV64SXS8GfK5u6vihGC6SG160cdyTKtk6zXU0Slb
S2IqAAajyisI3GbecqWs3Mn5h1ljRApULoy7+a8pDJCa8sRoz3HFOcKmRIh917cyOoXs7ceo1Cbp
Q6gxCXeIcJFCEe2HCdsiKne5wHPoNUtecXl1pQPzH8ziuO0e8Bstl009ecAH1axyP1DiNgCYIY4h
f+nGwunvgP1ix7RKOInDaLOTtYx9Dv5kPbMvwLDKWpuwWBV2Ss7KOFCQQM165KCKGvhGJcPO+JsM
CHK4HwgOygHWJ8yDF+adlaSHjXzlRxfzERuUPyHPVVr8fRpxSN/iPHxVmQs5b9Fv6gSf4OL/SLAX
1VdWDI7mQARKuyxQt2RWbHge/9fxvJR7sowIYj8W+aeIdGbhE2BaXaCHJItzEyEaDY2tsO8KHWtG
ryyUuj8udt3fDYolgl+cpmrUznf3MNKOX40xAUgCWiN21dlGWWhKhBuCOB692jCgqEVanJsEmLgk
xCfLwW93odeW+2xeqY3JrKtWYs7cNNHLQBxHepJZovP+c3OZHYoe6Zvk3CZMOXdAzPTCAH7dmCDz
gFpS9CT27KrBM+k1odt3M/alStM61WewQp4Mk2d/SXT/+OWbCGWy+7vFEFbb+5X9j4Jnabdi74G0
8X88qtfynLfUCO9kqLjD+MpkBrGouB4jf8lRvCaD7mOSWx3OeOEUIMsDs77hjTBsRkmlGZyaZ1ME
NGoPgd4TA1q+PLopv39kTJJdjailsvMmaU+LbSKX9AOLL1al6L2O37IPuJVMQSY3c+ep9PaQyvXX
O7KqCc7EtNGMKrqL5oBW2vJa+srwNnkLPsicr6wl76JvBKmPa+8zp9lRCcuPsJV8l+kcyu7Wp2YA
avNZqLcR6aVTI3i1a+xhF4QCAwhRXPbm1EVBk8cTcA4OudPIhtdkUmLcFEdwF8ikKniNYI/Wva+N
J5jpfBAufyhzFDELx6CjtlDuPoVNWOww5RwQoewCs78IP7N1zV9vF2erLrkmBdksktVyhEaig95h
99I/kAJBgOkY88AcSHX7q9U34Qej/SL85JxhpvfFfkzhEvJXMxE7HWoSro3E4s0L86zZa/KgcNDa
pVqEnC7ZOeTADwh95LD9frGkb0GbflXIHpFAS6d73qNUs/piy497t4grC2xeCrAe8GCyWt7ydEU1
F4CIHrj/gnp/Q8uyy/tBKP0tH46ZC1XmkVQftbO1nw1SUFNo55zWygNxAenwuo9Jd3YFj48F80zN
92nxz5GKWrp4aGdkWV0MhDC/TAfym1NvxJ66VxypS4+A92c9puSk4ybvLPvCK3tJKMH1h2FVkrJy
cDgib0jm3uwTyfGB9+4Z/YLbvdFuOQa7hHI4dQ3ASGK4ykthc9OW4XvIZI2w4jcmDSXXtmRbLn4o
PlV8oZfZEBaePgrTuB7X3ZddZZHHjjLW4iUBoNQ4g+xJG5BeV82TL5zWloOVfxHO6RrFaMjVBBDn
v7BWiv878p9SxXIQucWsijPRbqRoE80ubf/vX1PlmCU+R4qe8VDJt+0guInQLmCuKZKBLluw7M1y
NK+1OYC9GZmQhbGuJ0Y6MEvmCqh8um1jV32I6ihMFJQq6Q9HT3JvkBtokTpPl3lE7hReKxy/TTgq
Y/0X4IcYGBOwBEFkYajWkG/rbGGqW8Rk//UuSMa2YvMAZEWl9IWv9JL0ApGFV1m6TpZUrnA8Olgc
Xo2vBfmT08Yc/VknPosT6wTE5C7tT6One401DJVtwf1FZzrRRD2l4BJVwkHSL4E+AO/EC9M3WJia
jkaSvcc9wFVU471GC/HqAcDQC29i6eMm8hyDsZFp8du1UGvq0Odx1x4vfqXWeqVfVARV6PfbJjx8
f7kQj6CmZgXYYA3HyeKy236UM4BaQD1LS7sUHLADOTzxW7Av66X6Pbd/Tg4ZJjcrFYwNzIqOEDQM
yd2StnUt8RqTSohKd8ZEBtmjKr67fKvkqiI5XXJrOrgpLi61SdqBEippTPwFW+EiqPMZsjAHM88B
sZhp12IbVT4HpX/n40QDeu8SGb4y1P+xZgW+6SpjLx9XptXv6YEcbB4STyYyitV1sAFkXfDW9CTM
pga+kN07977KnyOJwrSDjzUqkPFi+PUspc6BYe7JlnCtHCDdenHa8i27fDuCZ+9JfZISJCK9aIUC
gOD9z3anccOTiqRlpxz7sOa+O8nZYhIt8OqbRADcBrSu5v+EBAb2+tN3CdBBFhPLxR9m9eWv2MR6
UmYoYelHIm8r2aONEyYje3oNkRgB7VSX1xvnL5+mEEIvpv6vlfK6VGg9WAblR4iHOjSBT73xLJ9l
YEyqj6WmuQPlPwR1huLtHiaQYB602by3Dvp2LQpTfRh7gte/Wl2Y2v0NeGO7IPky6kgM5757WL2Y
gR4+EqJhcCPKbOkxhQbradX/+MAlx2/eeZCLB7FQZASXGuaOclkpxLn9L8ZU3uabdCEBtt1dMLHT
2iHEX+FpJIxBct8GN5DWVEVYe9lzh7TLMiDeiBHZsZyz+oENclx+oxlCPaaNu/0B/XA68Bn/m39h
5h6ATJwT3NRIOcT+AaT/SIzdS2A6bBln5sAvD1wHvtoh9rPP2k5ycLYT9T3fkYj6bgLg8qIQ4/oE
FMeOt527pZwbZZIM/gNKEjw7IKimYMZWfeNh3sDo1HZ8tPzAfdPYCHIlSD9Kbb8L/6/EeMA1usk5
BKbl5ER9kWRIKQXfeP0XG0oYUazdTArgrpBuE4xp4JHAb7IYaLY6D0mIP9FCCofGysf4wWAsNQiW
Jp8ZHon62IF7WBtlBTYf2XuTBrbmSRHqHoVjjygZkTqGahC5ux0IwOfQ681oEtAW4uRTfTq68CoA
aY4Q6mIXH9/xAV4UwX981FxWel+KIQ/JSY67BXfZSLtS7VNf8CYoUwIx+I4KOmnYZjZ6dIhIU5uf
LTwcQ8oqNndPMWPgcmj37SttRHfzRG1xaP2AV0ZNDhtzQx0dg7A08SdGp0psnwLSj9VE3tkUOtaj
/0GCq5Jn+VGa/e2qtVs2KB4aIm84AKW17XA38GQnxXiyUMbs1LonbJE2owtO7q4VXWSuaT3+QJ45
m7LOd5THVXqveUOCoEKFhQN+Y2+rlWn0IT5xh9tMlQwBHfgPG4a/YvsqSen065wqtXhsA0mZO41Q
j+KXVArKrzl6Lw07JA8KACMejI7q+eZIodVI6C2Eye1GhuXcwenSYlZbDC/bzZ4+nnoCWoPxMxnN
wE5rO9pWKE/qIoqlUfO1CybVHwJ22kWarQcF/C7Dgw5iOWxk6wXuDhlM9C9DOmrGnleBbEgjv9Bn
RWVhtWKe7NOG5g83YhueWNyC0NXfiRAVMCuf6V1bBcE2F5b6QatM+oW7opabm3JcHt/tDiDwnwn7
mlS73GbtAgt6lxOrXRXg5ao/nkAFp//r1WE7EbZ1emV7P7m5efQ+T62kHSToJqU0sea1iuEPsRUe
4uyv3Jq7zZWjhYlcKQsNmR62Qvcz0KYLfBwc7VWFaKLvuzMCPy9Rk+L57A0EdloL0YxaI8NOAmPL
t+Octhvy+TommdDwUQdUtPkBhXvqLV6C+TPeT+RuRiJ6x4oT3WHsUWEzVzCpS1TcOcu/e4UMw2AD
vJ+WwwNph+jiv2tBp/7ou/lsmTtzsVhL/5+mb5biD9/lGf18kUv1Zx6QWvWSnqRh5KEE5/icZGvh
BcZXVSNwqNYLAHvbJwJ4QgOIMP4yJiThONJADH9HzzhpadFOTuEcgPmP0jC5/DKwMoXIstkZf1Sw
bxm7oTS/FEMQrvyvR6tXrKMJBOlDfY7+59kQSDlyrgA156u/AUqlJPzi9o7lG4XAoQWR+o3jXre0
RdPaVuVPlk0y2QxgN7tU7kcuDYVwkMwDe39n9lvj3OqtHS8f74HPjbEUmBfJvoG7JPqQ8M8CUDv8
LPw1F2qTj24N0OqfiaTb692iAvEF79Ty7hqHBHW8SEWaZMwHfmdEmLIcJzqxBL/ByAlYhX+mcHr4
RuS+JSgyIjUmevLOEbhWGIcSsvdcyijkY15y+6bD6WWYRYQhTshdWk1XkFs3PEGBSBzkw3ZvrbZy
WMw4daKVg0tq1oOwBqYrcWpAut2H7YdKcNp7nZ7YHLxPo6pymFCyfHZNoJrWRds5YSmUVIMbHeKc
SfdRuF9fbWvMBabxb+389zv8kisF4mCrzstUDdLmDmImUlMJXh6ilDOJ2PNbMwaTyEvN0IOYxFzl
d1cNWgrqn/Yl8aRaBNYRmJB7P8EJDQGKDJNpIdEUGpQSTzz8MUtb39dcrlLQSlnATxNCXS1rrwkf
c1uWkZ0+xUK+0rQLRO6I+MVUbshnvxmwrmH17rx+Sg3OWp99j4xreCdcyXoY+cn7UUG+BQiqsbC3
taINr8xW2m1mcciv5KDKsgBg3iOG4SCZCEzVKmVzLJgmmiCBeQyweu8gb48reSHNITNpI0Q35ajm
lxzfe6rCJPwkubNYMXwGfpFaR0W7S9yO+iZEdTeXAhz7eUxBXKWNTcZIXMVShqEUfAk4h1Nmi8Dt
od6GVEMHytQASIYZrbrwN9FmHX5jDY45OdUS8stbkZMzkUtHnkWbYhWyG6dWyjnfMgOuZayOdyDz
HGxiz2uyg8e2v6ME1G4d51aWj7ZRLRvtyeWpVip89KQ2FHnpebvCJRrAgPaMRxc5v+cUW+ZuR5Lq
1fqH3X7tomzQ9W378gL5hPJlefUjdnvcRRBVu88KDs/byVdugc+2/NMRpTqfOUXrH4c92BX0+OvE
rqaV9Cc80iydFqBW96HPfXeemM2X/sLBCcaAYA1NfLahFyygDhgPaQUrh1oO7rOtida5/oyra8fc
TiSvsojAHZW1gNY3cWMOqWattDCT4W/EhD0dPcqeKRPgG/yJ2ZBytOFbZ60KDj2jWSnT2C7HDrpy
ZF1fTgmyBf6T+CVYl8YIO/2a17Fa/3/TzMd2ZYSMUeHkB+RVXCKruC+Hv/IYMDhcAXMSuB2HLeuh
eidpXW7OuQ7ACofQOUNv1L48TjFpC07N1EUZK76pIBM3ekNtddREhXB7KXt0Q4Nx4gCGXJH44Rrb
24hcFWexp9bh9Or89YfQS7qlE++95rwPFgj6KZ2hrbQaw2JL6TxNwxUpSV9QSKBraYISgJAw3oa0
9pZLrfXMre4ZMA1tg90Jz5KlV+Te2N1UalXVwCwbpbqGjgcz5lhpWSy3tYKNfeHfruCZPHOn1C+z
RsxMmplD+QdQ8j8WKCpGCT+zxCBlQe8dN7C4DejdgX29CB/jP70i7XtsKNMvvGoH6pJeWrXOctxa
TaST86iEwCrrakOAcPgEefRwJhIzONQ4e4zZLzL6pedDp9Kh4xAw8PLFbQAuYgIyjJtg7C/h4Ej1
rN96yBhkh5zMaBPFRxDgArbVuyfdu3fX3lpLEEtCmI0XpHEIOWg6gSgyPutz2LAsj8DT4legVeYy
XzqvPJebP+h6jIl3wQiuDv154RzujROFtaoiUoD2LLPMMBxSR/e9KG6sAfac8hYj0Afj5fscsRzj
OWkh/sjY7G+5d7U3xlSWauEspgv1moCHSN6VYxbAODHAGJl6jSCXiSUkxKXRNiLZ/qN+a9iGdbWp
Dk2kKg97TwDQtk10I7nX4iRRVzQVicEOSPTcxqrNhULvqLZo1EeWKGSUOBsYYnpQmIWGMb7Mzr0K
3eVQ6XO/tOaMtYG/gbzz4oKFULuNaWdBiJTYDYvddpXn8WQzRA+ri6UhOhhG2vCoanfYmnXqLCYt
qoDn770XWhMmDc+PUpriKdFZWW1SFzahoc+BQaNB/zX77P9yk/S6qT9h7l+JHtge8dLNw9x5Qx6C
NTNl/2DVQOZu3Km6m7k7YqxKMJGLDnUSAAra0DWIprrTLceDiftf7gZA4lZQvD5E9SV7VekhYoVZ
f2W/ROuaadhYLq/YcYicN99O9yWb5oByo1VyfXEm87I85NLX6elV1oyHZu0ISTXHNRcEkE7pfEq1
Yg3Xy+ZclfSay2G/vNQBt4n8WHRyj4c9pirxHeCDL/5jF13y+VjOu4/FfFK1aKw68GIu77kCAc6m
NjIJ3dgKXzuDg9p42cv4YzntQWFyzI/MpFcHVV7vZ254+txnh3KY9qXuc0vkH7/wmnpgmb92l5UD
30mDtwCAixLeGrobLbYFjkoluTM7N3b4T0rt0UZSQaGb9Bsfdptb0ajzpD3GnBTEXv6iW/5IeSB2
4DKmJWXNldDJLqIFBOVnqdkuEHgwx7xpBnWSDcLUYVcuHKBsVtRRd/NPMY1HsI8ZF/Jp5SqKV5To
Kx1H27m4++O7AkO3fEQAwk5Lbuz0Q+1ySelqayQSNCUTDZAD24M2TMpfkooKj5atPZI10BWuFfnR
YRPs5rLpDkywfMU7KtGhhJyyWlTjs4dWFfutnQTREN26PNcjQPJmjhhPZyhiRjm4BTMm1fd3xMPt
gq0aj0cQZihjWspQAFCqiKkSYMtIt9ZkPl1bvxtsbjGtzd0JdsWz8X5GIeEAc2GGo7Jr92ZF39G7
0/jEPz+ll4suDXIUlvbW8M5Imgpybz85eLlxRlbJLos5nIcQ3iPE2tAfdkefWzwQgk6cuCmxP5DK
kuvmqT5kqsAGqHMnxcaMDE2sY6yolb6LP5uhye9mCsdQJbQ9AL3EVE8Ll+qpVAyw4wYBSx5GaxsT
hs2DVmK0MhwaAbtFRv2do7dzRrXcxKR1eEmhX+6rXqtzJtteTzirI+Rm8qx1EwCXPmpCUJdv/H5s
dazhPB3HpznJqFJF4CcI5O5rWG9RCeLHr0BOGvS7sLDkPzph3cp5DfWL2hqWWGyMxobhlBuhg2DQ
CZRpWEMDc3q6BF3rEJjKwKRGmK3RwXvdPYBJ0JXcbv84YMd3ptF2CNGLEPKH99ODN5LGMgjFF45s
OEsKvqp2KdWim2t3ZmZv9nULwdK7hrcY1xr4WU5td1//6goxzAXTxClu0CHY8gxlvW++aCM3qAho
mP7s78+eTQG+IrgvqSUICVW9RyKOMUmYQBcch8nxxZe+totzHSa4IfIB18pX2H54KT6inUz6p4RZ
35RIkT2xSYZsZRfhNTFQEE9gWXvPWx7eXkvQGNSU7uNVxefhz+XxnZGOBW7Ptb0V41CgJp/5Tqn5
HtjEyrt7wEzge6LqS4YTg5pLna9SAXtgTjj5Wc82ztsYtJZcSmPTcssNJMwcixB1I0hx/4sU4yq5
R0BdZOLIoCmkckf5oN9bacKGSQUtRbeW0uoYn17JwfaTakNvloH5H76B00sSCNS0N4s11KkvfVUF
0n0hZt+Tsp4XkIWIYfqlO6Ostcl0C9W1t9B4U5mvTQHbMjq6PIODlM/t2THONttim191NpiSJXXN
ytJwIuDngjMLw4SbEUphCFowi0kWlAGs7FzqemZZZRNSFWjanUgqOGvzekybCOm5eM6P+ttzoly8
70uxQ++0bxgwqc7YytI/4P5AYBv5TK0xmpwJKB5kF3RHS+OjLFxWIyBrbzEMaq/lX76LzbzktyB+
Cmypb0GEZVJXD/RR2JlS+Z2ivxkuVxq13DH7P2kRAnsxJjXLFXpA1/aZk7riHVLpOPC3c9nQ1KNy
Lrgr5WasCiv0mdo5ewYC9oUVAGyK20wu5Yk11/ByWKusTf/1l7fI2v+4S5O5eawu9XfJzcdD6df1
SXGCX6s26LHP21yWufyT1MFyxPydO3McpXSHXhdmLzWxAP+sGlc6Vx9mzRpXX7KTcgFP5ygtqV87
h3VV7OUh568LXi0dlP6lLTPdf8AOkL8H8I+s+Aonk5fqhvNy3cah9KDYq4n+PVy32gXxdOgmzlLf
1k205km8JdM23Rnjjbz+a50XZnCdseOKETtzyahaPwi3GGcoN6N6yQD7QQhXadu53Us6qrHZmbbS
qffZAGTfxR1NQrUswiX7bxb1fw7WIUB+EOOYtaF2Rn1o2ThadE2HalNSIGbRz658hcuBhMFiMScj
f9AmO8GPfF+iDXg9/OjkIlavXhpA+FXS6ijDEegnQzmYEMMRPBmNlwZP0K3y5u6I1oeNU/PJbVhx
EzofPJpiYCY0ni+Q2y1zKqEqV2UThYMbarLrfg8Ottu3XDiLw54x+WGwbtvg9TirIWUJ2b5oTt/4
EzqTbJ2gweJVufhI9EJn0Esz6uv3boq1pB9WUzGC0uqijXDNgGeIkKGn+F7WWm1uWBhd+/Dtyp4u
m2KUN6DzBSmCWZQSAgRWGgA+0yIaVxELICW5Vzbm6VfiZijKE6WREFEszZIfoJtMX8xR1AHXdIB+
AZWtY/1UtxlIfETD+aCJYKiZ7Jf5GeQg1ghFbfGosBG4d4YoL9GtA8GOVjsM6cVB/BzcFvJgjL7W
VVKDk/dWoWK9SnjcPL9hi7IMdmtXddVf3bINnKs5W7CJxCH9M9xlSedNjISoLe1NZ5xzdGxEmG3p
UCFWJcrLgt0/dG2Hzh93zRDEz2nYazv2rftgsiUPQ9wpnzbOjqpTkmDlyeDTcIV5XSvRipiGHl0g
PZgxrJFIlAGVTcrJ6PRmh26lPEFrC8/jvSGhxdz/Qv4yivyV4iE8Pg5QZikBNXZ+b0ZXBFn1mp1q
F5iyd0u2Cpr/PrDz6xnJnZ4t7uEhy462yVU0qc4Xeo+CiqL8qw9T8FwADZ7/f9OU6pLLL0EwuzT/
Og9W+WADlinAK+tqQMJXvIr9rpb6WdGQGdHoWyN8NhYSAJaRzUPCN8sIWFqNeOZRLZrJApGIhuC3
M0Om7CKDTRzxAjwyamn4VHu2I7P7aa9+0z8n1suwNdF3lq1YlZh3TU7hK+6SgE+P6WHAl6JKSwei
DysQlcKibdJsSluLcqpJfWCeY0n8Gjy9Y6RsUiSlvynJfKdLE4jn42MLh2dSqrs7486rUQ0HIqS/
hoIeDCQNorCUS+wLWmWjTMXpTMen7Zo7qpYUC6YXHo2/YOWzfyEacwCdcsXlnmvRLnw5/mvA5WLF
DMLPNYf/DWgHfHmQg+V0WfzUNvW/Tot+r83rmnDaW59q/KQqN3jAekw+FbQoIyuAs8/VgQV/stMb
DVxXBDA7kRKr7G+/CS7MU8yMIOT4as47cQej4XP9t4sxH+96Br2xK7mFbso+xwQqd2GGd/Zz1ME3
28Hfieo0NGcJHQHSwlfLEwL5vVXqm1N0SeSMHwcNxJrquEDMd4jqhSL39GXHNP81yKjmKJZdZqyu
Pe/rvmEWUqj/vtmuQRmbP9AO0Yhe6XcyjBTnEvwJqFMHFU9V8E6hTTNZh07Mso+0+S4m0Zk7L7hb
SbRX5XBRanUOvxeX+Spf13g2R0TYPVgtMwRf3QcxLUnIu5L+KfIWSBADAXWQwDpz1mzkLZOM3Gb0
YUlBT3CInkhbzjpyGIdvkjevny6yLudWiMN2YC+Yo35nq4MzdeYLQfMj+SqgvxinYapRNj5oC4sm
F2Dl2zf9+94Z/MYG5Z5H2jwIO9pkcmPp/wag1oz4o8dV2PrzCQh0+f0MwMvnYYZvqyY4vZ+kl7Zr
1IkyBTn5EongkQM68NkW7BVLL1BpPW60CBVeB0yiT5A94rXWOmI5fQXIdBE59gl9bqcQcqjT6AoW
6ROwcIVmsGEbKJvREIdiDWBgUhVeKJZb8/4D13zUpaGi7QaQ4ktt+K0YpdQfyE/J/UtEbXUBPQv6
6Qeq8iYqWwI17gUSuUVYl1FRIjtp1KZtFQHH0WN8l/64MijtLe6CWkWneaPPhz1k8LPy4ESffNBs
FaEByn5eIEdlVlPEAHPrk91ZyAFX4/Cnncdvk4CkldErF00/3HfL/AkFGWTwF6hhuLiHwxx4DiRK
g1N9KPBAguDD+NWMQrUPy6lKkzarucmLVU8K8pKaUSS5cgKGNTiGkIjCWWgY1KpHRTNfzipNROlX
hSZtYNRebdS7vlotbOTz7tzzqcHElehtJUKIgEEMdaR3rohkyBDAvUaqkcUPB3osN1uuKKWAPG3D
PUM1u3dsAoJMqQRAqVy+vs3mPNz/KR2848yA2516WlNKyL9c/fyufZp19kQQlTdmpDKXW9vYDTK7
xv8V+Sf7ZaWbMb0F/DzEkwmNqGoUxq6JXwLqtXnRanPasaFgs6ztbIHN9psZUyrMlbI+Jp97s3os
g82/ToExbjG8J89dADcYigh7NyDWO+VSR3g3C9QS4HzGCMy913vBJ38dtOh3uHfFI/18Jgl+nYmC
TbUrswTiXe8ahleLvX7yS0nGGrM2IzihckBlsgyyIWCiLF/webCvy/nvObuaFSS+qq7+42rg7EEv
3wv2Xg3VUvA7n73A8cXGburoEmp0Q7UXgwsE/irR4v55Qk9J/CQVyyOXdwsaE5JlveL+NvrfcfMe
fg+KDey2nJa1weLWvAAd9hBEh126X50vqmLJ8C3mlqivaiM5OVbZBFO/woCGMuhoUd9nza3zlQ9a
UGrG6Daojp5V1u3oWIopfpFumu8KcwFUYT5yL4um5yBugwAZpoGkG5z4BKVKLrYJvYf1YY6dndnM
leFc9VzNpuWsuub+HsvrX8OneiWE4efzKz2KPOrJ6QB+fsYxzAs1CHYcVqXgyntcQcPcMlDVfZVe
2h7r7+J9texZ87qPnWcBiZvu7SwyTbq7x4YbCoXO6jdkZ4NJsHPTp6LJKHJXrhTQX371QTS5fu5c
I436CqYI5ilrZ6Lx2GWEYXdCdv9mk9q2ltgBenq46bwQxipeMm37I8Kk82fbbyrl7/W0lwIGh8cC
ms/tam/uAX4NrVUKYTRLvd/sH+28XBDKJXK9t8jhX2A/gBNfJkJJq2H5zatH7/qIYiXDTM1FUPIi
5FiTYNY4ogRfUG5o6z/e87gUh5U92Z+h9bHyzNlKyTlP12lMmu2nEmEOc+NDnTcNugV3KDuAy2R0
QHeUmoA+PCCLTL13wDLapaB63Q/4y0bt9HmrMPewP5v9xsxyF223IE3NEEDvgc3TNCsEfKMJf3SO
SUnxGQHaueBRYqYs1Ap7T3qanyxQST/AkJiqg0ZYE8bTkpbvTnKwAlO+hUjpxU33yxRu1QsnH6LC
I0ew2JYtbFmurSCDsHxP+nTAl7L0QYtq6jOLZ63omfQHVD3KRVLP5ZqkBbMmaWaXobWloZz5HqOR
G3v9Vr9BuoaMsnwcOoEEH4kAinPxuOQEpJlSmxFs0eseJvbTqXJ39r987ZsX9J72Vy96AYTKSzlK
pBuhwR2C4cEdPdjHkfARsc7otLBirHouUvIZgvgebVH5xzckV+/hYsToliM2IiymCr8/zj1qi4Q1
ggVISM4HddxUsQ8vXT2Xmor/ZhxQ/sLOBg6PXg3oLl5IPFLFxlsii6bWG+xUT4/OUik1nIBb7Rqm
ghvkvXLOLnc5Z/+lVPcRV7FpKTgRR6m3Ufs+REPQ+41xQY3x9jRJrJj3cJFZiD06jGFwikptzZ4M
O+gjRpNQhmlGr7JfRlhOFW//0QzQRj+9KGXaTzYDG6dQgWBTwdSqOotiEvPnpO7kSTLYI7kuzAUt
XLTXajbWhbCXo6QikOOC7TxVULPNTL9/tu3GNbZx+50SUkhfDBhL6Cg4QPBPFNos09ExynM0MmMq
t/fRrJeN+QHgiuMqCiRtJ7SKxeB3FvlDt41pbdy8S+1OnmTcEnQ2f2DvMfx7E3dITi0GKH2dSQLG
l4p1xzc0gUSMPQbGLfq+s0fqzPZWs/xcFVo1lKNmcPczfSgmFmYgjfFYh9XVsWx5JzQ482vtfZw9
UPw4tiJAqgyGW5fDDLlYv/enXt6a0InsMgpcJWDKIEyReUhwz4aciQzohpEkcQDDqad6a5CtucRx
pa9Hx4XJPcjBXnfec6CUeqe3xL2/q6kAXkUAK/+pT/TRjMonQMjuH/iAYeNuIsk38yBr8BHyJZgQ
G8gHTyLUw3ZPdToa+M/pb+aXph3L1Cz6xjNWZCGm2UFUPQdRzo3GiZ24RJqGJJxAM7q3UBuZBI6X
cpWhRZIpRqCFnU1N2LP15fjLUYiE3F56V8mAF2iX1RqLoM32pMQPT0kSZvqg5jc6HWKs6WTh1JQ1
cngnWCy+/gZk/J+p53Uc84dMi5eEbbVUj4Ra0rj6C4i8rYX/bEHjUCfHO3bu2/ajfYjsjkzOj/Gt
mktKOzRyK2QeswGYCTt4Tc4RS1BbwVcBXoI3mf6dsJCX3N1yOc0p7gY16ZHBAXYqJ/DCuR0hKwND
bDqQFH3CtXr6/VdwOTK4ddDcJKkxtJ0hDfPxo4C35vI7iwWLMHqNnZyjB+EyWCzh6FD8AcO2K2gS
XjXrPHghupm5sgGxe+s2hZk6gaWFXTua9eJSNi1STEk2mOBVyN3b+r8l4CdQw7kfYbsuk9/gzUFy
GDzoMJyUkYP2EOoO5yY1EL2lxJANwovb+ij5+pcAL32k8Oq4EYpqemDxSIDvfXzdSLkHDYiW9/7z
evdG8jRxLmcrr1tQ+4nzL0lt3r+p3oHUMuseOXnm0koY+8hHfpLLTfKawLnx8oLkTqWXsXizhZ+D
yzJKzaPC596rr65Ow8BIBtrcWd2wDRQCrT3nfznzigOr92c0b31VcSWe5eVvc9Hrh+tW4IjXTcpW
la4wMaCRu2yKEyadCV3EjGjwWPstpW8KgKvXPeOFCDXkV5SzjnS2D7yGn13aeRpV1YqeKdMSe5k1
w9ftjVOvfi9snvV3rhcPo6bdLX0rHYrX2VQOXGmpGV1fvbqtZwOGqDcRIykexi5cdH7QaXovvofQ
ZtovyQfylnWULsBMopZzGwnQSVT7oMOEHgfbL/Qqgr8dzTJ+iN+hyKdULi3Ql+sOrB3GddmFOVml
LIwEd/+O+pxwOd6l6s2F/3O0PSpqPLJAzYZ2yT+FxJeYrQxJJHqimbKVlfAXbnr2/dlKfcuiUP8Z
qQBIASPrMt3dY4g/4DEEsV0Zm5nU4DM2i8dO11IeboHnlC2LNFkjPZ/iVyn6BZP7PiwDmTdtHxWl
M7cUrQP9iXOi07UGAFjOGDIZE/elqsPv0QTZ7EqYxoA6dhtHIyVmQupzG/4ATLK9XAWxFUpOiYd/
1vW8WEAveIo6VSqeEm4C0r6qciKjUXL67lCPPWrs6Vbkx813LCqeXcLSruT+yeJg+Pl4TMCFyqw5
blS3VTJT1kMfV9cmKMBlFlnMvjeLUNIIsLKiOx1QaCk4xbzadtxMgYGUc/AxbT8cr+NAmvW66X0g
MIY0ZtvAPAaafmnhtdRWPmfmmvuFoyjcRujz5nnZ5pm/wE1hto4RiS1cyZP8tmcvShaQtN6tq3Ig
5bD9CfrDB6884mIGYmCuYpJ+e+FsS08GSjo5LVywynKO6mT9kefLNjAMPi2MExbpQLSAEXgCly4L
RO44IYtIyVxU4Eo89XccLPVHcKQ2D1JoN8DhigohJ9M/5N4X9HCQCq0dC/kCwMvAj6aqUWBAbb/R
lnM9Z4VJVGlc8erj3+CXZiRyDnTuf1d0Vmf2Gv7Eg8qMQ5Anawi55owMCCoaze9I7gESHHCtk4YD
2rmpYKf1uHhrq0YXHkw+QQ8m+2C6PSD8PHX0e51pz4ITmtx4L8KIX92XDCMCd3tS4kxd8nDRdU5a
uS5NpyKfacN81PNWYrDAvIUV09ihFgpWkDdHDrU/W5bFM60z6kdo6lyOpLc1oAimVYtyH0qtw8e9
E+PIcqlTnst14hMwfuOJa4gUSJcaxt9RkgyMNRRp7waB6gNEocZYT3Vk5Ey2i0aH3VyHSfASIKKe
q6+0QRHDm62O1+NuIhQsQoOOlgcNe7qmOFPeVrC8cIvOyri5GuAKouUCyRxgN0eofp7EsAoHAcdi
cr5sVy+8uOOGI5OgsNCcfFbWJjRlfrQqgwsfhiFAkMrndZue6JmdZ/++YJGhOe2IfMG2HJN9J8gE
AtaIbBCtOf0v5VFYXnkm9sU/DQSuAc4TDd6z27evnlDjFsyu27YvrOMzb71gxV8lTiJQFSM+y3RV
wA8HNuHM46AgSxtHD7WwqOgz0hQ+lgKakNvnbzdP6MCHX4QYEjhue3gG5wTTw7xqeWauc+3Fg3ct
a7CbRURT8esrF2umfSjZjbt37N4idpT1USzzk62KZKvnuR1GunD9dySgboShGbBuKyTUZ9RoI+uq
h57uC3YkRPzgXzcV5JCcxl12m2yDdK9RNzdDsV3YWwvUoSZgqqCGpoBrnJnxoFqrcRAPh21kF6sy
DUx+HZYelBtpXr/Cb6/uKU0kLpfemym8/34qjYlVfwRMVqQn/8NCopG6M3VgoKfH8/RmV2scfcx/
Lo7QW1MYIWx6Y8GI5fcudTVlGLy/unPIZtCyh6UhfMZcUtrbtVU7m/Y2ZAWSvWeJcJ6VsFPOzx5u
Ai/oJO3aqEod1N5QOerkxqOZlNprDZGlw8xC7l86KXPLiyJyYOlqWtajWZ3iopmkVTig3ZHN3uB0
v8+DsW66sc77GsQUq72UeUJF+CxPj9nzcTGaFtfdTC/wAjcrWSD16CBQORj1wNfC8+Phi4cBM0rC
UeGBSP/HqGjulZg+1iz05PltS7ZboszCMWuOUcq61AofD+pztP/7hY01Js6gqjUPntb0Dw5H5uR1
/8FeP71DDE3Go7VhUiwPHl16H1UK6AuJJkCMNhO92je9ugDtiWw35CgyC08r2JTLY//Io54twkgp
K1JdVv4kcTBcN0ACwuKtwRXOapRBMZp16FttvzIw/3mai/Hv46nfKateoNXyt1csvV94fxttTPiw
fMVWN8DkorRhjUcnbJ4LNaQJeXLESZNP08+5AtMQwpNKaTDcPBV6mTmmz7/UtQpaMFV3VWMK9cRA
OO8pg2gq3saf+yB6ipo522KdWPe9x81NZyvZI1i8lb4xzDZcBrWdWZ6gAAkeaT+KZtRrJTMq/vre
leKelcGg1AvGymvgfP5jKlHqa3gmiYDrcmxxwjWkeyfAM7aSD2vtGeEJc7HYTHkjct5RCD2um4M1
mPxeNfj7YsHSJr3+N1W6/hSAhjyLLsQ5uY72DuE179qOeH4MpnhZbknVcchxNx6m462V2ezA+CXb
X3EtP95QOerJbtAc1U3bhQKQcxJGWNHgdAoER6PAqc8qVPWazSW3v7lxtZ2DRvyYSS98yzB7gi9V
VY9rykLKN4wwDctrnJ4m3bg2bDn92/mEfLnsXA619RspOtqCMRga4KgoT5JCkMoWpWkj3DeWrYwn
SBYYKuF5gkH5ggxBS0llX1Pb6xi16dQz/toeBgi+liIHPzuhGqK2KmTisFDa6hnAm1W0KPERVvIJ
aVk4ikb9Y3rxNiLSDCwr5JmEZ+lE2ct5zunCVm2+TOmnSmWORz+zJzj6DBLId9rXyI4N1kMdyxox
tGMK740qGnX1GwI0AvLGtXEyt18FUtg4TOdUR6WtvU/Wqn4kpjNqTVnanb19XRuyt4XlnrtF3b70
oC6/oguhAUYJWl7B7JbEdvO7OyndmNOW2jb4faGd3gMP5X53hQfuO1Ea4t/wgrP02EX4W0fmOCuh
IlGfeKPeRJf+1j1xQ3hjyv3XgAaHwQIeXd2vntLR8O2aVIeLPfNXHV+egDq9iQpy/JcZR/3RcCtN
Qm8wnvg7lBn3VnjJEDq8bZQZSt+CccSIBPbfq6kD3lcbYh3Kgn7nvb7QnBahI7pY1xsrsvF6Ih2y
A9sSi86gVUTrU2jR9G7Li8qoJRYKj0INsVx9jMYSHIJXQCSyziAZjFYO5tDlySCUl5OUknwRBvB7
wVgR2YZCx4Ed7OpfCthvzHFj7DPv1eFi7M8fEyl0HXSryK2S9bx2/QT2AkRLff+ShFFQOnNcsWt5
gwAOGwDaVBO5/xOWSdxfaWNT3fVBWzQEL6Dz7Uaf5xl1DQnPA80Xqc/KPTKR7NAzMgrqvKImnsK3
Xbsd28KWnAJ5g2Mzbo//bG999ffu6tHKkxWAQP5QJOQW6cxZR2+CTND7S5qTVr3uCmrtVET8rwvB
Iv4cousMkltXw2nhfBLlJtvFAKQea0YZyoJqsvwtZ365Z1nZ2Hq1l7iRHi4pLyiEE3zp6axkkKcN
Ipls2526s6FTIlF9xN11B7xQ3te+yrXEy7qNnQRI9A/oll94HhI3U+jFUsDA4N4W1U09AmViceML
b0VSs9xW3zC8VddptuheB7aP3HnL9i0tEzGt4FTzsN/uttcu+tEKHjPIG1xmSqpAN1vdAlWhuUFt
RDtuv0UHqeDB3EaF/Q8kFT10IpAjMEDq23fII30wjZ8Zd7oOtlKOYZ85ft1046iEhLfe8gMZqq3i
ax8atsXMfixkESIdKwacg7XRBCPkiPr6TABKjRzOo9QRJqU3lJLqA0HrEKcoRLIdvD6h6Hh9L+Pc
RVMOpLpBdpdhG4O27CqcBaIWhmUTRYbAnEQTyLDzkkKctz5bvcX/JGWPs6Ia83aorUZ3bLD8U3xk
3ftYlsTZfwBojQPrGr7upSEIjpUoN8437sQUbc3yxNE9lM7JZ1Z30BoxGjmtP5w3pDVoQCjSY4yZ
h8i/4ROrZTTC9SJfj3HFF3wK7JE+Vcd3sAPwmr9GvsotiqMI11pe2N/JjM4TK4IvvdNNGWI9DfXh
COf0AMNqL+l6FkheCsKA8V1uhhq5vViMsR1OTseRaznnzkkn8iYXsLU/eEdQd4DPrmkZQJkL+fwv
RA7Q7W+O7vhOwUiOo34VKQemel2db/3e780rJyVeCR6ivsOUoLXrTn0I4VfqW0rRSrsvPN7Do5b1
x6CZH2YGQxL3cyU02gLAHLUJFjFsX74nvfkF27/90M4yB1DPMH2OIV/oYW0LNH9ismMO6u2k5Zib
6lzfEZ4OjfKJDDD/5KOiv0vK8JOQwwXOcHBzGps2QZ5rbRft6zBehN9F0KLCn+H9IDCsUXPNfE81
DC3hgGIBhctLrnwbHaPAW9WS7LyXilgcimxS7ElYfef9DZ9wveVY4J/vJ+stXzfzx6NQniMcvGwx
8A+XeED7yXfU3rRdUVDnsUj+Rpy9//z1luuVy67E9qg2x5zPvnhx1tkSBiXBvhK5QSvl1w5OfBAV
BKOcQC47g1L6heuCPkayc8POPFqNff3nlPnC626ROMUF8Q9YAHkDMVqv+AhytEWy8ZNJSaquA8Sh
ZF4rJa9TEmMxR3fqJmXC21RG28PS6IksehK9TmhtoPN+iPy8pDw2Bad59a2/Cs44o+5nRaIPvptf
zeV3mRkKdyucWVWz1MM6D/uFjJF5tbAMSqi/4w5eQl5GnGs8LHmDyR1uVspU4KISRGMREeAtsStv
aC3NtiYwcwpko6tBv5dWzFBESDsV1ETxKE5wqkoE+7CH7sQmxddyXv5mm1+hAZWIrTQ6mdOG/YIn
3WvAKTyLjYMsO8AWBfPiUjCD1ZAzumEIqFix4tcCU9h120+uP60Ig6y373+UY02U69SVBWkTxekJ
YY4QkCPxqewugR39QcEoQei/DTFS0oJnqNRrvzyV9FyRMcNGJsvLsnI0Qf+95Un+vTnsmoUI7VAQ
Zyg4QtJwL6aOe5c7NagwJYQjWnBzUbZog0Wza111d7mmvYxGwmrSwYGsnX6nFdQM3to1CEG0CC01
6VUBum2fwKBjDaqtkLbhgujAlQY4RId983TAJ6is/DOnr5AoxGifN4PkAh3Lxfq6s1sOtalH6KOH
CqzgrcoK0xpSNVgJqvB2DBR5mP5yNCICrZnrix3Opyh8l2dy02zy+/v73S+ccLkgf19tIFTRl+2P
3G7BlHi+GRMk6YB0DiXvT3BssXMGNuTs5BWbWEewaIv21sE09v8CAqwchovzKHP9BFEekeXARdwY
e+INDVdew1PHxZRcyd5yGp2T5VanEHHIsnQ6nkrmzBTQXEHgk+uIbATujQXYYRp8cAZJ7YIWJ93j
uKbdNkRTjwe0XGzbIqDRbELFqToxK7ip5/Wz0KcLtiJRKHvYNebJrj2HxdiGtYb3hlCFtITU5ouV
lR4CE9lFFHQdVWmrKgZypZcEwpOuaVesUkZq9EE68z2lckMmRwGgD2ODqLUyllzzaEWhFPzd4Yes
DRGIH1S/Z3w33Z3sN2Oevs/OhYQ+0HX7Lg5c6ZKcnwpjLfMW88pfyFYacKFlXg+tJBoxY3UlizVN
IEB60EEX0XeXyMPEAbUUsAVJLJ2/KBik4urGF1gYDZh6kAio7T4tlhikZq3BFIimn9SxJIbA2OYQ
v0PCm7YrbnFLVjVHoznbODC2rf9tYMULl5SpzyEEl8DzzOPoWGozSuAtfxNNDOGApYuatiQIUQjZ
JHp7BaOArzDhIdppJ4iRjWOddclmO99bxKadFHsbHWm8D4l7WA7iQ+VrObqm6a9hPqPluVgEFQDV
Wu4MN89/99uoDCDhe5emW0RtOL7sjIFEgNL4btCP8LU/ihSAIpHs9MMwhH2TPrR7M80IqtCuNjBR
5QtGn6QAWyszKIyVp6MoRfB/8WQC2bC+iam+q9PsSFT5eqrGWMdA7kAR51Ha90vQe4J+pTKVWXsp
RKCuka5TJ0YJ8bfmsp5TW01qz8P8LXCT0s5/OISDhVFcZuQgjJN5mKNJ1OmOiKRYly/xVsxu4dpj
QhTzjAqv15ydAIzXrrXoZ/ofF7MWSX9/bTZ3p62HBcNUTT2QxdWIM9bdvRiYhcD5aBLWTw6NKS2F
qxunL2fvCbx4TKtLRsxjybq6axydtoYlJfZQQunDqkEAMJnrSXTJOC1yKleDnqvsPgBgDsQkB0ci
JLKutqf2+1SXy4aOfsJ6grOsOyJpnBmAg+00vBmsZ35NTbKhuYM1cGmaUX5RKehRgEAav7f6ZxVO
Kk7tQO8V035rvPZSxrwX+3emu1SjUkx4F4RtXeu1YIzLEVLZBz7WavdX8De9WiDaFhiLzZhRKgfv
TqnMSyPE/K3taRmF2Q+qmVHT2whkAhxiTn/bFkwJZ7OkAiPWcXgpl3/v3U0EXWc0wR6iBX+jYMo3
D6gul1Ro4SquAQnCqt8EKnvGOaI/zykcCjEmbN1DM8Y9cRftiZyd0WYIEMdditClAmx7XPlRQvEd
gSftXzfzhkHv08RVIqPqq3T93+7PFk8kXix4rjiEy8Lzi+r+qDCcZoOnvBHVq3mNrg4lp07Z0wTa
W5C9DevAUm2nXvPkqcqL4yXUkNLJDGn0EEan8ZOqMEH5V4vwF5zz4qyHwoqmhMf4duxQ6bb5pwtT
ORAU/nk+etLsQ0/9TVonKf8trzI7mXrxv4GMhJMVHt+mwriT7jm1mCCzNs4pC3TVFMOcIj4WNM3L
zSkoEFXBMfkruGM7dJv9x3qRue605At1uP++eWMj8gvre2GBrtkLbWEFNZU//XEnP3K5/EGGDxEA
Nq7CiyYdcCVKnON0MGRpGqs7xrVtvtT8p66Zb+h0Je8Mw03l6mb040Qj/NN58+cXrpiDAwkh3Vim
gz4cX09d7ok8ym45kuMj+IvsQtq7S+YS1283pnkKvqpLPw3F2KjkCnPHXKhGIh+J0dnIu1FFu402
hcpgn3U7KxdPhK4wcJ4fGAPo2hVeM4CgXE2petVj0d7gSfKPgnXcdu40oXQVaTm666YKdH8ezBl3
d2rBCgSbTFhvIdbmpvtBECycgdzv/wW3sy1uiI279G6A0qKXKRhRPrvXF9Va7G8W43tTzgc5RYfQ
o0QrczKOeoBD5R7cv44YHSQXcXznFMtjyTAXvpuT+ozeo2UEWJj8wQJfBSBZRmfyLneXx+plTEUY
N7PhQXStxhZjrJX1NmixFvG8J/DuMd7X/mGu6dONdfdfm4muVuUGSSQcvTXoTl7niroGyhD+NBbq
3J14Tr2CW+4+P329sfjpM33OCzkwLrt3kHGpZXEWzBjYB6pbDIjQX2SIiL4QlVg4fPac9bDD3523
kzvTO4Y7gMRCaKIB3Pfcx7umWDK9eaoVwahng7d5oLb7T4aNXm7BN9ZjSHRFwgyjsFJ6qBX6r8sJ
EF8JP+0JNwI/cRmYDfWcpekm2ItNBoSgDtZR+sn4pao2THoj6xnaBSHmnHsVQqTVBU2PNBmNBSyX
bAgsWW4KHxszxe39gxDBUMcjac7fKRCYF3QNebH2f3VM2TBYRAgP3YW3jfy+GwVo4oZAP/JQlG+P
tvUo+ji80omjjQt56wv0UaXXh2lSQUHRjBkIJ4K0hQMKOp+uyE+9g1jwGgOhnau5FLncaFrv9dDA
mRJP4oBIuYY57spZcfxk6GaR+93MG1Ucph2xqml87xNGq1raQWh6v/qEkM+Uur/v8BQ50LkOi8X/
aGin/iiejO9hc/vYdaC+X9Y4+gI/Q6MsmC/BsOHTyMloHKxogOWbbLiXDj+ITHJuU7p8ZXj2GK1B
SHWVHpwikmN2zbYCLw0291Q+eRaqa4HGxuYDS2ptInq2OeBIAWMzPmFb0Ak8ZJE9nZzgwRHDFrFv
Lku2/rGdxiNMvO4eUr2Sprws+gBidNy4MSCny/PnQsfpg3FisvzRXj2CxCSkxvU37X3G7BKL/fyb
7f0OX4XWf9FlI3W6KSMMbzWq/WPExMAnZtQKC0/ow1a9CCFlh0fjxMZ1na6LSuvy8f/vwZEgJfzx
PtfkwsD8FUrhGiW1pmGDr5Gd+69lAQ/8RtzUae3DFZkRDSgyTD0rjRbSIi/h8dFJF1KM8b2ufqk6
YLQYB0s9vnTf9rKSv+3VgXx1P4hqp2FVVj0TL2QcMdRGiMHgZcFHKvjtK+7WQnDqGn7XdgmV5Uqz
n3+K3qb2O8OPUrGzIs+s5TZWvN/eT+DzfmAtJQy4gsduCXy9uFAo80P4CXj4Z+hxDT9VINycH/YG
rpPmYHaneehC2nBfaEaG1qehDiP2YxvEpKWDq893bfZJJJvs+dHtOlcbwYEr4ShgVZjh9oME23lb
AYEEccTmKXt7B/p0loZ6o8uELtqlXluXqZs0NBWZoBVbtGYhq6+Ux0bDWXxI1KYwdDiZEArDetN/
Pq3C3QeeIs8P0IVhsE71hRIrR+xHW6uKkVkV80EIgcjSxFoSmnIlnehjq/GNC+PYipSgvOklD/Vi
QobEdTGeYvHrtSoxNp+v4szyiKHWABRYF7ivNm4JyKa49SOMDKnOyr2sVqiDygEKgc5dzcIpOPSW
1imx8828HiXclLjQ16KsIkQcSkUwCrzHDLK0wRiljHaRVvMgLD1T/GQiea98gwCSa8L7/r5wdOSI
z0V6q4LHJCvIP2Ub50Cu+fM58kWg4YtgQ83yfbHfjunGz32HeJ6ygXBgiANcBFQ72SJEDTnORSk7
bJQuqWJH3B8B4VIJLYDmYXtIzp3m5WfbC+mLXzIJAbdMWQXlaoEfk/ONavWps/1naiWn9uzSplum
mjA2LzLOlZHZrd+d3OtkgzZmY0VD1WBM9laVr+AshE8ddXCxGVVr3b0dw+h3o7HqxMlIPjZmFrai
8PjQ7BbUhc/4rXmJcAD3xQEFpo70cChPTQEgG5uG7GzrLEXUqSkQApmimlnXxUmqVKouCx4Z8FhO
Pm3rQtHPcKdvMbGdTZPU4Sn8WqNA1VjNiOj+lgou/LbHaVPJUb9VHXhLUEl7ZfSrxeuBpjN/vD+N
bxyw3YH8xJ97azRDfDs+NPavhsdMkosICwXyWdIXxWipGwlhUL1Ilf1yqdzn0GVGRlQhRdRhX3Tn
Ybg3topXlw3JgdhhfLu/fsGbYzf30QayDH+r+qeevnExspZHOyJOi08orNUEyfPGMZp8QWzur7ch
ivYup0j/wmIbliplexPpQYBlGmbawHdAkkUghEX0NYX58lxPnflEzivyOV5sWirQDh7/uNyw873b
QrhH+FM5mlVS1HPlWLcigImsPOpXj/BvM98YuaIcVjjeLjqHfc8pf4RuuENylLBeTieSp4UkH/50
MpbAM+169ixJHYZ4UiaeBmsJS+SXgQ6xywhu86Nj/GUK1M7Sh/4aLgKOSALIBEtwTZ6/DcAg//Ot
cZDblMY7t26ndKyyeSzdBsMTkWTl0YrMiCcOlNurAPZ+yup1mWKoB/Px1HaE6sTclO6/l98IS1/R
f+UrqLq1h4Zkf5uYZMSLtva160dH79brQqEAHJ3vwI71dinyXDCaJZLDDgDHTMvfPfhxAtm6DNdd
RovnY7dj5EyASMeWzk4gk5SVYeJIuyEYoujfmOZLHyPbzEMw85f9/6yaq6pbaZO4ZcfVsow7dDbT
4yBrnYU9a83QaVUcAvKgl1iXdqHyS2a6HcfP7z2f9f2OEM3YoUS0GR4syLtf06lIjPmNHBe+eh/B
O3lsTFUn9xzUbHKcjU4HfgQ2h3fuq7lTLiRgzl09au/zyypDgogwwXd07AlqVyYQejAkZCVWODj6
KAcCHh/xZ+LsCI23w3mFEai9VYLfxmqDltjgZMmvWulIr1tey8Om8hL6Y1xLlpHNwMovYTL4LorH
1i8oLo00/Gs4OWZiPEuunwaPitZvEbYV4pPxxGxIAk9u/HK0jjB01hlCxWl184fpFfj7qTuC6+Ch
zO2VbihiMdu5wyTa3odTbwXWnzgwATm11VUq+inHy1HQv1c6j0uWN8T3NnxA3T8ASHbDadut9d7S
NQiYmrjVbvw2d9JI9sVHO3zQJ1tpkVDvNGuWT1h9MuK4xdZ43bb7BjUulTTiv/cZjyF++Fn/TJvq
BTy0nFLH5LfwQF9CB9z2s/+GRbbx/nOa4uxejA1W0icpdH8PvW0CqUMRGxSaakNlucoVfVMOQV3D
OKGmULPf+rJi/QWDL7ooXOANSIpAbN1Cqh16bIQUK1d+ll1hGlO+fe3KPH6yObEVEpijUXL0fTay
s+hsfCKp73o4MYmNMiImO+UDV/F8VZsYybWp6NDBjFO+SioIHUDmbMoE+el7MHg/N3zP4lKHwTvy
oTG9PbsC0WkzGPDUpo/pshVMEzMryP0QYZ2Byrtx7RCLqVayR5xK+8AeywL768SljrUrv/BKGU+r
ol8LNoDNTVcf/a1eZBz2w3TZgNeXHDmaZ3AzEqrCCHMOA/eeg2nqdroVIa7RrbS2WAhaS/cVCdkk
5+DvXJw6sEC1gGUyKO8kzVpiXWbzRqEaxw4Juj3ztF1GrWnGuEeg3vln5zTlHgTOvqWaH8rGCJ8z
uynS0XIWrKvnZpdJeHkadOiyFMTGGnQEaHLlEr2O88xWxe3IQiIizGGuf4+T4mB96ElXrrnAJjTc
u8jb0ulyYiAr9LC7iNe5wcRlxJ/X7b79YHeZvmzp13I3gfGCfC3NPqoEBuOG/+D9/1m600o3ES4E
Gwjk2RiAMjTCje7jm/mExabod9QfFc9AbSNJacR4zx8Hb5cIGfpg3fCo5JPAQuURivQ/VISLX7MG
d0/FOHlDgLG2twNrGAQzfudRp+/OiR+WTjBfjxJCeMjlxOXqhFLuMakVtJrPc0OKHeTyDu2t4yXm
broq7A9Fk1oBu0bgi1HI8lm48U5zQMv3tH5n9DMc7ZjUQUsNf289awVZfjcTDKQLyotBANqamgCa
gaqx59nK20FXLTEoAGMt45wslATNbHJU1e4l4FGA1f0IZKUCgcehhOK5szjxaGfUTg2sSwGKeXr5
Rf69VksPwvG4GQkwMXkcYPczB4s0xgx3g1sP+vgYwF/whoyktDYh7hBgkrJHU5huhrh2xoib2AwP
sHL/FiLwfT/B8wHsYgYGsxSpobAmv/iB94HkC5Tg+mJcwxHR5bN9yzR8OqYUXlbshnK4OBEL72XH
akMllybL9yPNuJtgOmG5/CvFKoElw3O7X6Rv+4Pi1e8RDbyLE46LIn13AChlRfIer6pdAL1acUFo
STG5ZDoODzihs/7PCYtUzHLSpL8HGxABC5xcI+PE67oXooLZRb4tiNCVpTl/CMSzQdXhbHZ8ceuC
oYCYoyKABvAd/hIN6cW+e5bUYGzf0CR9vPPnWtuQzNJlXIiGAoGFlfub6RiU4A7ub9LhvcYCcCFa
8HBl1aVeAESFN1rxqB45OaOsuR/u0dnpPNBWqzuVcHqzkSFbWNzAaIHevO68DgfsnuHeNfNIuSRk
QwFherh7LQuCN2n3oAlBl00Qhvsg2CzlxTeC03t3K0UxJKCOH5oHTQLZQFqcJAjR+o7VuNGcToU7
7ECQ534Xsm0uxs9bAcrU5GdsZNp8Xoc636biPGpjUrOKF6+mgl0MfZzGMSVuwKg76wdPnX18fA7b
g2W3lbVmBAT9X9og0Uhq9+7y+6UwiWNYdMqM8Bg8ps9rSDKfdVtqT0DFIK0fEo96w3MPTgIn0VeG
ZFjooNw6+SFylqktG59pAKusSWXZJMASJs7HUNty4aq6vPBrJfkb1JlU0Nqu1Y8Ei41a07Qs++CW
1Zf75RIZ6yF2oagyiJJvdUu6uSMhd1IoDirDRKyxHZuT9pcR6Vv/BsySiPjr/0qqV3n8nWLQ44T9
ETY/heNEbkRUvkwi8kgamKmb0JrcbzSlhs2SWOJ2ck0k41flzbHvIL3uG8T15oRxipR9q4W17EH8
03eWRLgTAMWvAj5SrztEqTOoH3c+xyqDNQKRQOZstw+RB5kK2GLrIZ3IQbNUPqMN8ahL0BrEXAKB
IO9Ep1nHqu0yHMQ3QgeXojA4iYce7uJ/tSvo0R9QMIVx1JkfIMuaSMUyTar/lBSBeWO1IX49w5Ob
YWCWCcX+WDxyMkO1Dt7GkcLaZoiMah8npVpxi38AXQY1vKAsWxXrfmvr0QibgYQ+XElCOF8i5joV
IgbaY2c0DF/ZhrCPc+tWss9aUwXywOfoBwDXY78oGoXArS2ZAnL9qmBNQ5Rmdqgupkl1vzO7rDAu
CNP9cTtC3ll9+JnkA4nhgIIAppXxCWDCS8ojKswOidNVZymx3j7ncmhZYDkpBgBXBSkkwPdn+jNg
Fkt/zEkIIgmCp5xyZGbRjpyWz8k6Ra3tWICLcy+vEXODZFyiw+o2VGZh3owFM8SO3EOo1Tt0a/Mt
lrnVyLNAMToLkrPJ1tsHrdmuApg5LZWEyIwT4s3qFlVUEYzusAZHXkepmE7gd4dGzLeATFp6iDe4
whwkeZsNIufLfJTwnLfombhzFaz6haMEr0141XEPyII1IwDdunAvzYIEY5gQsdxtyL5yV9xEA7F6
O9tMex4v4Djj2DjsaxvRwThPefn/cotDLjBxm8H/mbRg+5Iou+ANWTFxPr05g8+JFFC95cKkpfL1
9pFFR7PevfHS4ADJzLvrJDfTD7P3lgnyAfZcDRi7/2Bxi9myVEjGj3hMo2eRQE6McROr5shiRVte
T8BLdwrbHUHC2IfYRB5fiOhpvbo7cPJIJCrsml/zzQagOqmlB26Gl8BjGqIXFm7/HA56x+EctMFJ
Cwvg8A97X1xuyiIat/4lQtMePSGq8vCQAmxnH7pJTKcShC0slZAwp1sWB5au/YP5mjZHZGrWznM9
Xqn1Ut4RtdLaLf6cNk9xgJoY6Yknse+4m9f5zA/sFnKtlCiHR1VnlZhgohk1PSqnE5MsgtcJg7c0
jSrIWBmccDbe9L/Pb7RkZPUA0/ZMet6qBGK+voMnf2ioU5JozXge6Si6jZ86F/moRs5wqTPpmyD0
trK/m8pDwhXEG7asDYAwOdACJ+iPLJGZ8E+4eoVs/Rl1ME6gP0/+DZlfKfxlQzC8iP11ls2dUKYU
4EODtW/2NRxq+OBUsljeDQa23RVxiRjgBsZtr/bEp08ZsVqnfBZfllsx7o9neVpQxQYdLNoPqe8f
Xl5lXhBIZSd6RrUpHIBrDw/vK2QejkcvkOMddNJl11f9HQJyc4MlxgLZ/npgMmbNHhZ+W3NajBiw
c5GE3AahJjgRHAWPjFOIHp65h6mfrHNrl3xnnBLrW4BOOJbHPtRSAYFlRHdiqpwh57s+tcDpKZ3W
SOnYQaiaF2bu2lKhziUN02PT1gvxGOdD/9UeQQtmySP1KCEiHnpX249jB1SDvMQmGolXJj4maIiM
/oHJYp8WKfj1fzaFBXBKQqnXXV6GOQ5obM1O9e11rRqlBVKd6QAGSum1DlW4xYW09YbdWpMjHM8D
usQvtUFVZfIC9++g1UH6uIgTclxThHsXVZ4Mt6Umt+tGjbDR8Tu2r9yiAGC506QEzQkoFG3bimOj
CXAbmjhOjUYWpAUWlWP8oG8mLQlHCj0P1hIdmt9MnGj3LPtJSq9lh6LPdleN6wGKBrz/gQ/ToqCF
gGhcdl2tPtwXBy+isjwyzOttXiVHvvGlAGkkrzVra3mdwkTBQHlhyfR/G6U0YiTBBO5ZYLpsLb0f
N67caj2zaYlR4a9Y7BcXrRq15I+pY6g1oxdaBbtZa3jy1WwvMxON9m6n0JGUplkUAYeWO02fmVu5
VmiJ05t+Qv7eQUQbZs4Q6uBU7zWJR7MmIvvjmwUiEERQna3mZ1U+OqaWxztptAWAG2NI3CZrk/BJ
QmeBd7d++XvBiCbPZ8+lgv8EuKLhNjtuY0X/opyCDpd39rG8lYUF+jjaC2DDvlypgT+Ijfxz6QAy
nd8+OH+YrEH7LxR6qb8gj9yerQODPQh4KWj5k+NIJTUO/7ilbRa6t3qvWAciiaFQLapXf221uM5m
AWolI70jFNQBfdh3kVdVbYWYZdHwb2AcdfZemS+QT2okafo0nEJPEb+d8kc4a49x1TIIrwApoLF9
lrw8RXgUYawHRP5McXq2ZJ958NU2I2gJYnfqj8J6ui0bhCInxVSWnJjiITsKsACB4huzuPyZQ0Qk
EYlm/Z1nO+J/Ow/zlegOtxG5W85+Qxby6edXunOpE8V67Yrx2DHFpEBogp+MgFz99DPhnBIEcYjV
pC2d/6v7ugbQgaDHANK9at1I79GPfB1KYPahR27dgRGN/IjIhlyzmYaAGYPMGRbezzgUN79w7Gi0
uKrdmw361+w68lb6nQV6R/e1r55IQF3KKtRjLXW4D/n0JuE5L77zfieGe1WrcQmIDfM0s4l+8Poa
zHRZQ5JBIQudhwb+cuIAcdzXgdEaU/xz9ejUbSRG+80YYPoG3EwyZp2ZxmRpr3W2WFEzj0/05fEt
85PLIYDLxYqot+pc9CT7yPlOnoIOGqWdU0XzEnaoh2WzT1MHVZz59psxOTmdTj5P2B58Sbl4OS61
ilaPOaknV/fKzDkN49HGaDi00VQz07NPPj9tfj+UPNHuxMZVBSvtYzZYn25J+jzWnnnDA8u45pqx
XtPTkVbGT+u7wUZlMjWOEdgzRdDUko0mJxo78sF4KZ8gff9QR4T+iE55SmnRBomS1xercFpmtHv5
XumJcqG49KA7ta1MLyom8wALpRw6VeZCwWSB1sXAPzgVrECuKLgh0+/BJdK5vh7BZD5OJ8MOTSKi
Gn5zY7wsqWzg599dFR/Itrky/xbHRxovUJKEak7tqrRx2QBqq5Eg66VySzOZgNMEsZTTzfg2ejUl
nJl3Lu/ieTRx6u83JsCMLjlHpy8Mjxx13I8fd78HC65T4SreiwZYUrmlL7gQWfb+Rp3FrYxK4zbR
07y2lHD6N+tWyz7+j/VnC1oR9ABbB5Gkf2zaQdkOadaAUqwE22w+ssJRFf6aXRXuVjTmeWDsTeex
63NY2bQYx2avEOrovrTe36CWQjbn7aruMrIfWIkjby2qQxR0VrPnTUcDqX0b817td1EX38FXAklN
CWgjlqpmvq2xdmn81lUOhVdNPAzoPH2TtcxYB2OyrdNxErFbEqcYKLavdXSnO9NOrhJSM1wwEKNA
dZzkW8Ks16EBCQezs+ABvuLL6DxUJc9JcE0QE7PN0UMRJrekIE3ZUSEyMSokB5oLLRgUPE65GhEX
N1nmV8+Qt7ZfM67cuVN+H94XkSDhMKpqDrhKSuUG01q+mcgf/qs+CUVxBTUfvkffUWq3n/04VPgj
/MjaJ0nNrM1DwHMOifiGRuM5Y6jPJxUU8fcTO9HQA+f7NwDy0hl2RfXDHZL4BLFvQuFjUO+ZsQqR
U1jd65zNeNBqGfGawDN3+ZpC3ecNzEFyi1kqGLcTdwXrceMicj4M5fHnRXJFfXZYqpx8L/Yt+f9l
Qw7A/swSYSpjnhx6KkoOSBVOHgGBXESrgLqIDVL//rrsEKtDQ+IDd32pmfAwFt1rFF61b7hLFm4a
dVmVnPp4hee/sX0sOY6TCPFTf5rQlnyqKGQZyClLQdirCCKj7PSXwfJXKeQ1WE5vRB2odGBlK+He
BepTBTlQBOiIlt3+V+N0qaWCy2WzUXNjCTNsEJBp89dQsxm04/SkUHUMq/zG+1augoRsS6dK6Zdu
cSe6tSHjxOo4ZzkXxs1OxQyCDytpvaqlhXV6s1jzyfxZADV/Rh/hKuRkYcq2smGlyr3tHVAl5EeL
tVce9T2lPQuMYh8qtPGtW7Qiojv4w4vrwVkyvfmjU3gqOBXh6I9JeO2CyLmfZFbj5zfmaWURV8Rc
tR6M02NpkyZWonAhTofvl6UMej+AIxnUvmQskx5iycXt++N9WpOz9IAZo7ZUDdxFbhPVlMCY53Mp
/ofCFvmNtahxVgmKg5FUsbYa7BjplvT+Zi82BexE23xrmX3HhS7zpSV7ue6prJx4bDImI0HNgJcf
gxAKRgjKgGx6QkZxGG+a3e9vUqSQxGbecRW9W45vhugqjBTeNKnV/OaRgg9Br4PrHMsToj79M8Op
U47SCyTEdVg8tLwHRD+KZhhNkV8BTeN0cZoFJoNg/0WsziOSWY+KyDwRIt0XOJuyvQ4F74B+DJ1f
GuD3acT1UjS+dDASZ/6b+i4u++5biMHLDs2mGT68LjTU9JJO664WL6zabOwkzhc0q/Nw+Yw0c1MZ
CoMArwCZ7zb8CXJYo09/KWQPCInDsUy+4+SMrC/7stGIGUkNvOTZOoA1nXSDjBHrUOv8im3Dr4Z4
T6uIzPYEKEo4sCFP1nfhybq3T9kfkTe2lYf1Scjq14DNAitvG+72aYCyAiHJdcBzeUMWQf6SqK9L
o8CWVxLWQmA9NrkL9x7ttUqa29GYDsu2QsitTg90HrbN4FO1JJ/BHZtnBnsvRjAR8k/k3fyXGsvy
HDiBq47A6tL84+52+dCsi/ZqtY95MFuciz4vbeXJXAmRJDranNzuChNQa+70GlsCJxM7leqnaPrx
UU6gzZEoqonAxpj5rBPQM8rLljG2wN+MPO88h9OB4gYhe6Jy6zMs29tUITPjLO0EaNHcKqOEOdb4
AivSzsRCAQBJ9e61kVOjFgh/1TCSdv63TkIrRLFcr0tWAC95FCQ7SCJx5wmiv8yIVjchUhKCucpi
EZ+jcmeFuQiZzae1zNTnNT8Prdt//f/bO53uxSfNjdCvq2uJI9HtStjsHLTegR0841tbF5YHAxn1
2nY4ABpPDQZ5J2Kbj8N6tNh8FcjCPQXJl1iYsQSg4Zs9o2ht+vMh7/LMHQT8DsxdBqYuGLX8K74s
2OEGxZdt3EWOQEEKSlz/fAiM0LEyhH69gJto3veYXM0QtQF4Zq2MWPdYh1WnAW8z7rTI03X6xi62
NBLZH/vNNJ1eXZjdIvX/xO7m8usm+3I3Akwz+nNppJgZIpwXC+iqN1YmeRP1Rl7oPAlk6HIvYioO
u+PSiHylUMUyKhDRJDepKyrtOx44fsxit/SApSZkBmoXFt9O1yptvJl/GIw+9hEc0msfBwaxwm+q
wmTH84JUKyIpoYj5LWdqxbsSURS88IkIVhkKu6GYGXOQKLjluf+6L6fTOzrEhzaLxAy0JofLuKlV
QTIrZJz95cQfP4HOJc+hVNNWpLKp65Hsns/EMYUhaWf5uj7D8HOheBl+kmJHKMGXeFCNb+k6iBRG
LH4G+1EaBkgWvb3qxwOC3riHvxapyQd0eQlxbekQ++td+QPHvic5L6W4W+F1ee255ZVkqA8sG3pB
cgcHqhAUcIH7jIHhTiRUcxbLJNtsxDuOb8t/qKvZ+gcJdiiGtKyEL8sWCnZJo3CK/xkdQdPErBUN
e87pIUtZEK7ihpCu+NBiNfm/LkNbNeEIKHLOHOkxkLCjUnCuJmgJH9oG4OYbE+v/h2ZzSq5UEd9m
qU16psr3/yBYUf4BtIRCgPvOkl6tIwY1iIfx0foShjsKFicDyYTQaYi0hRkgDwB7T9trAK0DN5jl
KVJ1+gW0bem4ChKK63wTLQTjzJMIwxXbj5d1vQzjQKlccCNRxp1XOgkkGTb93xmgdgts9t3z1Nh8
gW9/NgVcgvYsdmVQoVsb2N2CEKP7G8QaUrpfs42jRXp2rNHVi9BFyx0CJqpWzpA38PBh3aA9ixzk
7LLT1NKMXdxxRwLCutu9a/9U0A3YakyoJz3b9/WciJo8zITjowD6rBsTHBogVH3svvEuXtIEb5ZI
1IrfVQk4YJkS2+Nf4TazRqd95/U/CYLSxVzN22sRTa3Pjhrbeqdt2mCsLJwmL3IW5GBQuWbCILLk
nJlgrLQcajyL9gtidh+F7DpzQZ9Aq8lUgJMJJN9M7DtXCjb3D6LVIb7/FM2sSmENj2BoF19/XrjT
OV3ZG2PSH+zQSXAUds/kqMNFXivGg9yq5kcQKDgfd9Ou02TvglN7lBA9osQKSZXuu/uy7KNPdnKF
ByyUGoq7DGMqRbj0FGMlCcnUpwb+L7byZyKgcZ0zcMrSd97D5NblZLowte/0Ff0AIh87CkCl7rDo
4oIUIIoA3/H573VGYQAM9mljV0tN9n7leOhsBQzRX7/xXbeqZfVNaJ198rHannsnzeQKgPKI5Ilj
4TFL1H/BD+PptlEOgdiQfEJJNqGATG1VZ5BYG8UwOoQlLdNmemz0pupniYRuSQmtOKq4GofhkYp2
ou4cq0HzE6M366zgTddCpSnU08tOHzOkPNietzmIZ8XXz4LKzOSeKpTFNk7mH8UZyjPLmF5Nwh+a
p6oRdRsD08rX56DVzktsmGjy25aa3mV/yQ0IL66vr76mL9qQtdEnY1nzLLCWmwld3rolwkqc8EO+
9Y1woVD+R3eeIUi7/iLbR05r79M0nog/GYX4TYaYl9HCGRUa3JB8kK/ng0QRmQx7baK/8y5NP49U
TYc16eb7hYMPCvesKMAF/ZogUizp1ves7RJ+ihO1HmZ1Xz4M7RK56UYf5x/+auRk4LNrP7nLnIXC
5+dsLebbAz1W37Hq4CqxnWgLijkQvpBtEKA4tCu8ioGF4QSWBX3rN0az4whPXEUfaXmV+D4EFUkS
vwA/nAjV4scDeyKqIJR1+pXWsAEJi58LUJq/qWrZRp6g6YTX6R+wcOOpNEPr4oBGYvKAoHZqzVN6
6idLk85YGd+VqOewRrE/eR5PkqzEKTA2rWNE+rWVS0/mtXrOI0k991S2PDMAzBSM3CCmFbdrb+Gv
OB8A63I/LRkdH2CrMCTg7l/c45Zax/n+bftkYrcXWyKOW2vQvhw2q1Ez01qkBPflv1hb9xVeApzl
PjdrWbns8F4YOkfeSnPAox6IVuv0f6rJkunm+p73zTlajHnT8aNCfsLiLxQwum5l78qFStK9hfeX
FqENnsmEVc1CM9Bk8RHdSHc6eg7T3jsu8gRflfnpMZJ/BMGvfzTALcxiQw+6aLCa8IqXSf2c/gO3
UjUZBG0KHphJ4GH56gTtJZJGkVEjAYCnxm/z+vaL5s3wwEuwW0MSLPXDZXW6cH7/kRQJf827nldC
6CLTbHUzLn2D0hzkqXT+rtPmPyWY/jNTeLqDaQ4c5xkuric9PwJA8BXGyU02SubJvAOYSb9Igg/9
byGwPWvPpyvehAXM5ykpXW8kleSjpqTcyjdBBpYBndO0icpo7PRsfZ1Sew8pBfZz+Txv1/Kd045I
Ik3k6eDrF/ZgMLjX8nBcpeu7UjadhgtrP4E+wQ53ErqqPhFr/71yofGmYy9kXnGcREgyqulegfyR
Tq5bANcO2gkgfZhZCTng+ww9RzDehu8zSHLMY+v27dlNbE9AvkQHA6AXqNoMEgbzgdJtZn1TzA3Q
hfN+/hJ+UNKgtAWu01V43cn1+mSlswMP+trGMilYFLMdmTFh7lWFijzvqqlqW51VwsU+T5d2KHn5
l/GodOfxgQOJM4DOGtjitl+Qsmwz7zkhzbjlHSMUL1Bd5KpnzqI354ZsH9aZEBUcJosqM/kO/h5s
003j07wO9O9Jniv9PBp0iLWMenCNxM6BoOr5nfNiRqr1YpiCMfqELQJ79U4VCokiwV2caXEzozqz
vGX2Jmrqa7sbaWL44ZJnXHmDNRaKgr8k7HyeZ9a1TL/z+x4WWO9FgneVKTNMgPxmBBkQyDhE5kUx
54M+PbDbTe3VdZRMS9jl5jxTLt4Z03V34hJzk78gPYEelMSSB7zooaCXXxJlzWrenEeOkH3Ugycp
rQxJpyLOHmrnR32os5wYRsl9bSoAOrZb5qnkIJjclo362crS8nWQcgd7r+DmxA9y5Yi49G5jBwGm
6TGXiKKdiHIKro3MD60KrkUu0FmbIJZl2titIQqPu/a+1PAjfzN//mC6aWvqVNKcQAzTJGCuCoJ0
FX2fQLrs1g+9GXfCqbOGLtuE8V7QjwO+2qXPzy9CfggJSdkWhk+Nq0PHdXdqWAcChsA350rxE1Fc
pj9vgDHs5mrMRTYhKGlNXQ5TAbnLrpQwx0Ybg0z39qsUGsyAJbiwW2YNItxbmotQ61rl2d9p2mP3
rNpQLeGe/50I0GJKkwF2GDaGCTGPMEhFQ5W7ztrr/jErU6wMCS0R94ZxI2RtXaQoOirDPAblSZpl
oNeW/texS3pKbo7uTcxiqRBjNOGCCSTchH1LAjkvvw3bO+nA5ZfclGFdhDRuEdTfcEYJ2mlVTpnu
vG2bvnkIsV2yL5yeA+B+JMfrzL1qDYd6WDuA4K4TrP2ibeb8d6v9Lk3DdRyfKUl4QW+aJxgM1UdP
YPh8bIIv3tUOhw0ux9E9Tt9SLKHzCVGySOscjsIXma4w8aItO+FhzIZd3662EHytEp4ciYgOdCuZ
4fVsEVPI3NknnyE/5a7Ka2b4OyYKqfWu4laOTJwUWGLSUmZuPbvNyIErAA2TeA/bVjmhfEoFcuOs
Z8F5XuaI/efim311SoaEzU5ejvbr2V4N2eI8Ll0jNyByHQ3sUJYTlBn54omMasKJCNtUgCVaLeMo
yab4zB1IRPINntmgS6oJgB3SnVdkr0JmcSpXPcHXwPMmR54dZxRIHHnQQxtUUPVih1Ex2VucX87T
LQW+oIEfjZ+nNnxY/dM+m24Fuf50cVsjOkGvzz0bnYdhIkxx6gplqiOqSru8sdhcDyjNZbKZwz5F
KA68kS36hyOLZxQ9SvL5/uPneQmkamYRyc5WeYpQEQFnGOZFlaLDG+mF4XZIsyjMk11aN5GNYhsx
sD/PL7mTq0Hp0OpDZOexHPxU8KlcHwvGFyw2VDOoDm1cc1NWMiTQFuHJhFvfYhgJ1i2V2CMFGClx
XlorBHtLZQ0I6/TtBGoWyz252X4Gj/3iWF+9wPz79m6kHIoo3gzL3KOtMqpH7AUv3rLTazGgQuZO
Q2BRCUkVv3QC23jMr4gtkLRW0l90F3MVTsS8TjBzTYkPfOUxiN+otprQiP4A1hG/Wa5Ww3yjLmay
4Vcf4VMTuINJY8YYh9X8YwjUlZX7VEJV6EkqqHhVl8v3D1GPKMjmAdXk17War7s39wmokny1pBi2
1uSg98X7s7PB3K02TyxtEYLGcp8mTVLPVS6qENrHW6F7xreQFCV2AQ+c+7mQhsz+yeGvs5BkZKYu
/mXD+B79DPoh2hxYruXYE0a8c2fInCHLexfnJyiGOgomKHTVcQLc6UKLbVSf1HDfWlGJoLKRETUR
pO94/+DS3vIUgofJllo+nFrFWQDdj5yDxeagQ+pvIDHzQdi5lnLdrJdKRLctxfXTD+M0E9k67aWa
skOB4fEBZMX3oQRoDDpgYK5zGqtl+0J6Ro0Z7/Mi5FIiykd/6SRvvGdYSYuimhuR0chiRx8FCWFB
tlzSQLBwepg0yQWfWSg7YWBCzkWNCtpHU2dPe7+RbNoE6PgVJmbrZqHLtFeRjuHPi0SatuP7AlrD
g3jcOe0LLeUB+Vv+vFnFj/FDrj8Vrtl3fZTkpV+WAyY30DD2AYUq/7iKbr+JSWJRlRsR/vNAlMCo
UpSMRUUS0aJQ7qbsF/6QOen+f0ve9MMyBcX3CUgpj8Cpl0Pn0nyHBnQLpm2kcpKzKyqmvHlChQD1
n93B68UlSUyu5bsEaWK8KB44IRMEmS2Oj6gUZUvaKjFRAxDpPzyEeRIZj3vNM9GFRkknf0qf/m/Q
0UUcXaJ0KbsxwOMSc6kWHdECQQocEZSSTPYdN5uJhbjVr/VPZbYoczStpDaZsjyqsh17r2FEU9Xj
rdQyRytkENcqVohmJcO30bW9BZti0C0smvtBU8tVR1SqSYJtZBpVpAH3qDvgEryTCBmJCG+S8yQO
7g5QCG6ihL0C7K96KKSWt4ncX5sspPQqTBUcEtWZ/1hlJS6iLYfk3jVPUr11Wq0E6Hk3OgPkQyWm
AGTQd+ambQycZ2Y/29YSuTJl0k/DSC0lgk7TtwkzJHL7jCX0oxcVf0kXn8JNKFblnQB9QaLGCzyK
t7fTZrn/X0Z63r7B97fqDMqbU94N9eWqa8L7x7zjhydY+Wla0dchMDK1Sf996dxyjFFta9hqdPLQ
BDOw7ySO42FnfL17B4IT88GoiC6oB2dOcSOqKEMx4grHL7lmG00lLv3ZyNzH0kLiQWi5ZXq1h0xb
SDYvzlkgCjcVu5dRO8l/WVigz57ujlW+vPoaxoZTG1/M+qfFhjlFldMJq+jNwOm5vblSewALNfhf
wnDlbOGHDSCfMHCK9m6cINvY5OJsxXwTG2jEYXhhQiSWMa+SAFupQvNmE7rSr9M2s3ytCciHGVFO
TNFAZ7aIV67K47j7VsRvReGyoeFZEQAec4ouxMatN2z1TecaXziRvPJhv9Zs8uHHL5y/eHF5Biyu
Ic9xIwguXZkUTBr8jcY5TaVfitWUxcduFOCT+FVRzka95VdWQteUXJ7x9X/YxtpD2lygZDXl2wTk
1cZZy+Q4kaJeTvAOAeglnfkqwDHT6HOdGuZN+gZqjGJENAnIaM5YpuozBgyRoK0lacM+EzLisjpT
gNuEfdGNzqQv8VKE/g3Vdms1Uq6IqjhyjDQVKp1bKD9WWKKhGi5S8D/7kRVJvXCkBIu1dkPrRKlG
Ldxq2uhhoDKHUxEUjPsfnjHsjb1Tr31NjJ6hmRX5Dlak8A6WrotRxv3ccTj1IhCxMUU9gU2Br2MP
0/QqudeKCgL4fDQJUa/obrBzIzkuF84OGddg1wihULbMKgSyK+m/Z8xzBqWWGeIVExqMODrxXv5Z
XKY/lTT3duCEJ8h+wnVYNKCZ7186JCkTHiod4T4ZnFUrSeIxYS7Xzp7zlRnK8h9xkN7LLBbLgtGg
ZTDvSEvxNlWbQeQS9GyyhX1/fjD+gVD1+Mz0XjWoTuCQwHxUbX7F4QB0ZNvuJWk5ZLw478Kgapjg
lx/rVQESIXHdp42jF1hdN4h9xuv0qLxyihZKKdlDpOhaL7uU6lLKUgQZ0kZOaQqD/HoujttEnGM4
FsI67ozoLbz9wCfWQz2t8UQb2AgX5zezf+VgPuDAmXjhiU3b7D7oC5Dx71DYUKPsqbgY4WIjjJtP
lMHZ4GiIK9/vKUNVr9Nn+WodfDKxpZYvjjBsLfTxGVs46gt0FFETWiUHQerHzkX47QKMtt1KMJIa
/8y08gWisHO3qL+eHYih/37MLH7rIU+tEaWYDHH3lBuDOPFULIK3WSUTB0svuiGch95OwjMPBkh1
l9/pR0rDTjaR4e8Nyy60dRIQ2f5ORPbYBkPN5sSn7vsGTO65eBWYPJM4xBz7+jt166k/SkGhuTfE
llfl+aYWO+KlyLx9daE0DkyoPeJFC6DtlpuDkCJXrlxl3+A9uUNqY8rFrtL6pU9SmRLUGC9E+cAo
HfloQ/gKH44xGaSIexE8LKGUoy2e4UcYWFwLHaYa3NE7pORcx1MggAzv1c1O6xFJ9BC5ADIg6Mdl
BjUCIhwXY2pLOuanmmFWTeyCeaHQKGNubAsfOCsO9ogdNs1a97OBmsir7PDEo3B7vhgPfk3wTmlf
LTJPQgo1SNfXmkBtuRKd5g0ww/sXoGb0LV3aEjsCvVUCj+BRntLtl80Pz8CQVcZI24ZX9kw3HEmr
8bJUN+JuvTbXfLt07QpHMp+gQX8s1S1+r2Cxyo6zv67ldg1vDItce46Qy6uIvECPwe6S6IHxiAl3
jEq9JXDGUgA9+GzGhrFmyeWZMUvAe1adyU4tLYPlRTfLPMNlKyNoDxcmivTBw7CnPBx+Jq1wc6pO
d416yrrAwFhpBt4qaU0JYOnrJOQ8KoYKMqA48Du9BKoQt7ytJNH9RkZyc+0EDY35vs9yEx9jeCnN
vVkkh+j/WVADRwXV7KTnf0GU6y2TzLWJe/AVuw6O6ABl2nFkc44pLyS1XD6Ade59GIS+GRqhKrTc
hchjbBmsIWwXsZB+d2msGdv+C+4zOHM94MAgs/NSfYHZxo9OLfRbL/RVkqDZnBfGGl2oPuNiphyT
WZe5FYQreKzKK+EqTqnOyk6fZvO5TaHAHPoOXnB3cgUEJic2m9tSrkNytxAtAdvnGnzgDfPsuUK8
HPPctntAeDNJhAuN96LJ07XP2bw/mA4PMvFPN8cFKJvxTrGh+aQYW1sgCYpXEr5U7ktAPNOznrYM
7qu+Tdje3tmFFW+3z1/7Ay5qPxf4lPxfN5ZGpB3Dt57yWmd97nIJgWbhyjJJLZ6iIK7VwaA3x2kt
vs1efbTYZCxyERb3uGcu0Lb7efG+Aey8anb+EM10Eu1vWzEaSCi+5gx6NIxOrUyIDinOTdYnqcPq
XoTVZMBTYHuc7904CkofvJD3apVupSduoN6wb86NQ6O4kFEPcCcLm3MI3AB1d3dnYqih2qNRBv7E
OPFf8QtVSkhhFtTnnlY+D98nL4U9tvXGePAfGOof4UKmmGVK+99gipZJ1jm/mHGOhBqPwFQqgqGO
9EJtt+HPKmrJZ5pBt8Jwgj9jMk15rBNk3TjR33Y+n1z08Mc+pV1GpS0+uZpdZ54ZyPmWkhmxVvD4
5V7hHK9AGnzQdo15hRo+JbU9cD3PvIEoyDCXm3xjCd0u4t2iqsty4hT17IodjlTC3s9Chyr/l4CO
XWRI/zrZ0B/4Zu4tWTVA7ZuSkvz0VHmwERArVcF3O8tbiBbp5oufRoqMF6YgOF2zf3IkNcsqiydg
Zi7m7nnKBp2DmFycvx0wxNTx8X8K0gx7EimEMqFq8UlM4y6WZpKKWRPh3ipRqZ8/+rr89b6atF/y
9k3Z1pzbvvIxIYpLHWnmbhQmjL/1z7gAtSd2laDHPLdPjmhd2ix+PJ+zxCM1UGJToMMYL75hwImY
/V1QIfIH/6AwzCW20YtjKBDEVMLTDXjz+/oWoacjkvjVFLaZYitlCnYmrQ+cK9NrUQ1UPij9cCfK
PmU2oS0FUcmuOy+3I5y9j5m3sksBG5UxstANro3Fc+k53gOz/xf4j/kC+hjUoHQC92oLCzpcMgIj
FHXfbvEppFXizpJY1WoMf32K/HJH0gLC1j0wzcJ9f+Obz0pu9zRIXwk+lptUTMetRXlVpeZCTvA+
4cEEMdMi+oaOezf5dUeC6kdpTfvxeoD0CI2P1Alt5Rgx0mxLIDh9z/qb278EdLeMFA9CuFSaUP7e
6k28WhBYSRivBMUopAaNzDRmWiiPjBey8b81RZebrfMFrpI1PD2AWBI3CjrVj5zNymaeucWdK7P1
VNMWx1SMHp7bTkQKlYdhHhBqiaW3gMxvwGFxVglmBXUUsxJVHNKhOZ01dEF5wZA0YzlzAdWfkl+X
dHA9R1Ph5uGKUMDpv+d5kkSG0emYVlWt4lQ+rEQI9aAbHwumIPE6/KY/cFTOwVg9NtQm30YcozzV
wIQ5GChYcNXk8CoCww1F4+qodiVO6T8MYBearYWT41B4E349tgXAWE9BndLtz/01HP0rHFcrGSXr
K95bRcwu6tgNADAls2FaWZZXfdjigxvgh44C2X1T0lPntpjTYc95PoqZjbX86Bgoy2prZTFtNI7W
EifjLsKiUGUovRWzZ7TnW8QlhCtHjWdGO/4AjK66hADlzM3RhFVBJ9Ef+h8BMwx8va70m0gFNcjR
QqfGyFjKG97XC2tGNHHcsrQEwV1d4SBrB9saci7hlpS6nC8Si97dou0pqBFn/n/S4XPaSrY7CAvZ
urOH/H7UxMnUNE0CsgVZ01HrrccOP312eejh6+8Q0JalkKe0V6D6yiSL3d1AdfTLM8ar6dv0yWDC
aQJedmxEaZ85nkG/ZIRh3776PMh7I9u56aWtMaM38ndo8ukIsP04df7oK0g9O8kiwq9tohjXj5r2
WUpilL5OnU017kuutHd2Zjaa9/f+4bbo3ETrjwCrA81GlvxoEdcX3+Z+/KBmQZYhiE4QbW9smUjP
ecHYizoe3h472x6yeTcXVEg9L4NbQsglOjAZD08HEuudk2XXI0R2cQtV8OpQ8BweQHdoo0PBUppF
YgmJOewbU0AvXfw9jgQS0xcaXyvWISCW3MXyTDbqP44tePLxvdRehCIxxlL/wNt/gRWop9ivOsf2
UjruWzTwyXsay8zY0JckZJ9PtierQ+wnuDoAaYFmEOecInWaP4uzFxnE+Uc5YM3fR0RmApmdjP5I
i7aofUaOfsqlX+mpiYhXqpBQ0OdI2qUbVJhOTLJxjaD//JgMYlRmA5TOD1t9Qtl9Mr9DNH5Tc8zm
O1d+S/bpcuisQNt1WVlZFdl9Idxaq/41ln/oEjH5/WULMnyx77g25zjOHA9cefSTmhHye+od6/ie
yvo83/WCt9Mc2Oh5w0d9u4RAuaCRo7Hkeyt5kRRGPkPla3ziJBnxrfXT5xdO7xNAKMQuSMhg53Rb
c/PtrVT4c0kBWntOeMdGa0Jz42MUtj2yNpXsFx1byhr16R3WV1KdJgkJu/nILT2DsX8GoJCislx3
Q32hYwxVARLw7juNIQe5k1X7gOAEkA2Ee8Dq49WikVhYMeN9N6fChGBJWqztBXC+s87iONIrsTSQ
mFnuSEOxxTNd1Rc5zD7KS+nq5nPiBwftRDjJK1p0r5ciOmjvae4iSEFv94m37Djgm2EV9OuSCjhk
J3A8qexu2v7+JgFjOIGa2oXN8v9nmrrSY2EmHE5bqBbDcm0BYfCLX6ToaESHgBOcHIlAyf5OkUjZ
AdQ+48gfslLdtwz3wzdDqNnUdKqJ7IyS0akltr81VabbYt/8Boc7UYzmXnvBO9l5XvLalidILQxb
AbDqGnPwIac9Gd4fx2XHOu6I9UT+JTxG0oWo1uYjATZby4bx38l0WuH4XuP4a9+KeOLC1qnMA63W
0GUeL8Zs8cFBJo0oLE+p+ilUNo9JZguvwK0hYWAniytrWIRTUMgmlqCDwWP3Abp12uV1rqgy4jQD
9zxqRtG4tg7I29w1d52s2543d7jfc1VGB5O/oVfBVS5YarI738TJgUNcMxJvXc7tdMOJXNSD3nop
lsgQ5hz25gK3mESg9S2d4mUhFQkJGGG/gQZj0bZ+CszFLoEhVPBdwk9YXrr1F0GWTngkYNsZkfw2
vNd373ko18tB5WpqRuJAXnBUTDKRWaG7ObsJxLOhNJaVsPUK97UPC1rMQh0b/a8aGEUXjyC8hY24
l9ki+S16bd3dJbj54VszZh2kokNUzolWmJNHTtubaGGcW42BEo257H9psCs6X13ITIS15h9XHWa9
KFknh1MiIKEY9zRJCz3AXjnQG+6potZYLMdCbgI0x/OYrzoe8x0yJ+SvXu1x3UgTotQnX28DalUI
lva74AlXZsSCaCM8OPKqA9R91h9JT2NyW3W+P1XGiMitCKP5u3BPcxsKuEEFLJ2eNsE0IVLBpOjZ
L8FiEbtOy7va/Qj6MexCXoDLVeAyaCvg88gzA6pPgonmaGADeIqwv7ytLWsOEpg8emy/EGJ67wRb
NfmcsX1HgYDijl7hCm4KH0mLDGVaZhw7V15FQghMw9a3PkdDXv58PvtnQH8Z8HhRo5WLsXOjU0a/
NG9CtFQwGsygTeCxI9uuGEp9AxGv289lN8m0GgAdsiB6BQ5RsqKDJgNGlRa26ai1OD0lZEfaArpp
Tw/25zyAOt+BqochjSTjPL6cjT6VGzJeriUOKJqbrD1ohgKVrVjhcXrV/G7XOW0O6VKzmiDRwNuK
2rDgyl66X5BSrqUi0N9XjD/nt9acIaWG8NG0MPDo+ib2nKUEfazT6OHu80BTnpOvLoUsIpyjAlFV
9Q7UOqjGyTAORE1gCGP3dgXHYjcp/NoUURqy0gxYY7u5fNq2JlW0xAMPaa3pN7vrqibbB2bPHl4g
FzTytBS/jZboFqT6vb2uWjCVrTVzKwG8TpmbBEo5H1/6fvSmEkvYQtbKp+pG2vrN3Q7fjq7jzak+
Eved3TGUb0WKaSy7hz1hhGcxMRYlbstVrOfZTs1L4YEkJGVDgfCx0QDWC6CQ5kS/Zuimbp/lcEIA
pL9ZOcUDpAnHJyHxS++tseLT1zErFI+NrObilv8rbSVyhzf/4/W1YCgn7obGwXu/TZ0yS1pz23f+
3AGvJyer3WKw+pY+2fr/B5l915hvFTuW9QH4bbpWH5UrZPVN1GDUqR/q2mBTUw7Fhgo2gCVAblU8
+HYycddaTZQaCCygoXXBKi38k5f8piB9VJgLH2LEver4OC+DN2r/ILpNFHZyF8AF6l6bWZGO3y+h
DjuUeBxNTMn0T8vra9rkIKzo1ZFGALhQ+vahJbp7UStkuo6lzNHfMoHtNyBL6L2zFVYgEb2UE1/C
1qmZXfsdcg/tvkXFhKhUsbEhy0ZJRDoJ6pS8wDgHGpjFOjIZWCcEyvTH6ZO0BRIfTAAW9TRtt9JO
WsZkoUuVq4vZc3lV5M69J5ctJn8bpQ4f5HI92CEHWW3O/DBqHU4YUS+i7I5AW4/kccdZvAQStYZA
LahGKgzYjxVKVueLpQksTaTMQdn7AARqOG8S//1FYMuAigCmA60vcRXIhnSTc4gOVOeI9Hq8dE0d
W8upQEzXSQhcyGFEiB5nLhrfbBnEPFnduE0aOVqlPUwh8WSGtqairjfF+e62gnYcDcgk4jjUxJec
r9QOpI8Ly3YpiWY1PvVA2R4wjvBuKpyAfv4y2+/21gOwjq8b2O4f9E2X1pvPGN02KD1po2hryVwt
k9f6Pe08BtpBwyow0MZsJmJJqLOv3kVBD55tfdXjHlF8FZjM7y7enaKQUVCxNiIwDiaWMO6DIlxv
QtE4ZxrupaBYuH+YNR3XZCsYlgX7hX24Fl/MBhXUwjnS5C1DiDQKxX9uTp6PE1eVKArBPlppjyZJ
NlIuJdH8dzq2TuYBUqhbpmMfzGBd7hfaFssDJG40pkneH7EyA8sq0S7hcutj+uwfOMYqJjimTIQE
imdg8V9oytaHTNDpykbycLGRBj1vlmofbOr1OS+MYCeSt2PxuamZoNrKmduiifeZRNfY6aprW+qc
aGzoYG5NkLcPXH/x8yMdA65ATRRHWJjl7JuyfgmHW0YsBhhgR1rprL7sqKGw34pv3+3HXsSU58n+
K83W2PKqo0MODBSD9+1+X8+h01JiAev6A6NJN93tU8suA7+D1hpvMpPouFEbcjgeKRqobvisuflO
gwc2+dFqsaGllBPOGr5oEh4ae4AVdKsjl+mXFyuPO5OC66vHCprRhBiNes+jjiAFfYkuFoWv3qyD
9+hfKBSK2a69DF/jMhnWoqPekN5qRrK8ItUJRAnb5z3WcyrD/sHcFFegjWOH4OwZmU1WEuJSA3Z9
BnjUOtBiiip1YuoRdJAWX8v6u2tdj0rXRAblRrjyfS+OV9iuH2xqmDCDyyiOKFzxXdBlvBd26NqH
azfmVrI3Hi0OOsPFjS5crrB6iF3bz3y+JllC3DulsCcdvc9obBrWcyBKQy4KjBrMKvT3fejLHXWr
y3aIYBVNVOToBrjpkCt4o1MRHUapjnuZsjVXCii4tLKk0RNHa5SqsNeEAoWHaqP2FlL38pTaVG1B
HD+O/0oiLp7SAp0CDNgvp2ZbTS7fAwDyK20aQA3U1ELhQaTTzWhIvhMmFz6XV/4m3GTZX3h9r273
lB/H3FpcwvLqJ1nL9qQaBmhR03s4ZO8jbpHu8Wmu/ogVqXsCjECu4aYBdva5XmgcZ1zAQBGjSC5W
93Oes5/ZzQFQq0NAHHghsX3x4t/M9ORt5uS3uBKewkvhlItZF8M8lHvZL8TgQN82tZFEc+WrALF2
v0Ce2zr+VsonDf841G11FSlcxhFjBXDxro4+AFnOpG3GByTQS/aCfDiJ5WPZttiJhfoTCzztUYGB
Urux0fIRbzYWVJOlAWGWfdALsLlFbGhCP6bH1hUlmPdq5PDqqle/IpDJ7Bsj7sEwXIqwMPtWYYIy
ctDJ8Ehe+fyoXIUSPPbJTY3JRqaWldE7rJKZl0cTFKDwNikkFOMHzk01caLtgX97S2PkEl+xKmib
eiRZCveADKS96aV+Gl+ouRIvOIHId0K+Iv4Cr4ilTboNU2Iyd1GryNWTzGZsVkrUCuqZq5QJSXHk
5kbumvPi31NPoR77C4lBxA5HXmxfEBQZGEnr6Bx4g7hmFZzn9j5QJ18/yUb+OJ1skfkThtkRt5yE
8OHyln6+0mARkuNwB8KD5w1iIP6redp8hqTMEYSvmklBKiVVL06YF/IbrLYxC/W89Vv8i1knbAyR
lzGIGqihnkiRCqUfB38lyH+XekQHmEsYq7FwT2SSal02t9OOzoHBBRpI2ddhcr8HRCqG7KvFD319
VRk8kdsQrDSEFV96O2HqkSWjcY7l7M5/gKrTDwPo0CGv4faxPhueA1kM/Rt36U/gNCDBxpkHV7mF
raI6a8y5TX9jPvK64r07kKh9FRae5mycQKvv62iV6o6D2UUmon5zKk0sfccAJiqWkhxntm+BJ6iC
D1Eag+S2K6YhLGmv5tPulHn4FKb+r+Jco/Xy8gc4/ygpQsjTjZ4Kbm47EAULKdv5FZO941wGd0ko
UAP7UosL1a11APY/P4F7MbZoe5vrIIuWoFWNXS0uHu/NejGv7jPOo6ZUnG1W6w5eMVPgke46LKDb
NEGzs7MkHxza0oapcfXQP9h5Afh4P1qkHa5LqX/1/fpRPg2BcNH7rXNLeshadirIm8MJOmlvzgsF
HVCWd3ZcZl7VVpH/wMfPLu1vJoAGtogzyniq81WVQ+gnbUM6fCwj8eeacVlSkDcYmp5+JPHMGZ0U
PHVKoXhk+aKLwdARxhPJFbCMc0f0burnPuSTJHrXd68pN+yLd/9ffhQU9FdLidiQzvH1/4TW0CQZ
GSPfvU+XpNmv4Ag5kOq3T5CVKEeMWrFmzA8gJXzSUzYWY19XUBWGz9ewqddbSpNv6vmsafFONOfB
pxX2MuWadUfpXJBu4v78TM5QCdc3UFJjAAKCZVqClR6FaImKR9vEt0ABW6stxQg8/VBdgQT1JP9c
ug+7rVZjd9K8tHihMWUY0l/0zXGJoKeHyC1/waCjW6y8T53bci4KgnAlk8OAWgBwFiWmnzn0uK1w
NbqNzt5Zlc97TB3XJ0h38k0uz3/eoLxHWcK6yMYFx3njz3fdzd93ttI+jiK2WtP1iRBFbh9DAVW7
eB/F+n+aDED0WULVsuUaRDdfCTza3fEK4+c3DcJNzBdJV5v8+jRvzND8xtd5DbOWZ5FlM16ZuxZz
YIvKnHEEru7Ti82+wv0KVZKM4ioTOWTTD/PXE93AHOdDpq+fgKtO6zvzHFM8lHTvMRoM4uOgVk6/
ipudG3YJLSRKQ87KEbsGCJMuC+03Ewved2T1FqAWIZ8sFoWU+l6fAWEKQpux+LLJE5lKU6ODd53M
GZfrx+LIF8bEZzrzRw17oW5MwAAVeWSDjblr14zm4kXvhJWeF0bJPGQeu/vXicfGHQ675Z8SwSp8
z0C7hhQ8yHzssupIbGlI1Itam2oFe0gbl0NefQvojNie0sHQjc+qmJChTVjz3xdX7dzRB9BffgIm
Xif8WLcjLTYXzIT+GvdGkBvgmKrKl2TuTC2F72os9BUjY4tK/HNeg33x4UOQULMlbuwz1vZ9WvN2
Qh+m93AfB7Ogn0s8Gp9YLZ94dzrVypD6vL1ucEe6yS+la5UYYMCY7ymp2OvL9IzIt68cL32YuZpU
VYzsjn6d2CgkrR1xVx4oUwJ+p4qkV660VDsKpBmEeopeUsXUNmBv7kZ+VHcF9JaNy2mFb0IwIADu
5TY9kKJOZT9jUtILFlWOtpX0o6EwvJYjvY5lr/uKcLqqOm4rt0ejuaeOlnJjWPSa44Q6fpqxeyBu
lyv3aGOklEiueO36e0+5KxyouNOgRefh6v36NVzhM5aTjU/UK6HTDCvq9zCLYC38jzoEC9kk9Tuk
C7IAv/sUykMHRFT/5W/yy8PRfUhRi1FaIvZW5oe+EtoBzAzTk/c+AJw0lBzjmtkDlzAYv+t/IIwI
FdcE9VS+3aFAMxS5TY8929wB+dVTReFjWV0FO0SRNbEjjayq9UuG2msOW/CVWcV9/sEmXZXhtWcH
Lp8iPMxJZV35fJj0MBG/m8Pxj033eb7kceEYibMFfJz+0fQJpWHNlcXxcc0fxtqS66xb5EpXSxaU
7mfDeu/Y2kWDIDxxOoXVEI6F//zn053lV0ohiEwchjicQj9Eq9YtLS5UmA/FtdgbzhcOlgSnXzql
wMGEBuQit65yhB+7jFgKV7Av+SL2Sm5pU9T+I24eQ79k6onvYaztFqOxXLs+5CRn+sqdF2x1nG4W
nTSIHBWUYwSULXA43T50RxC39ro6bmIXu0YdPjD7oeckdNYZZLkA3k1zuwCPtarNbQ79RrM7bcCw
otygbVHNR5jI0LgVOukuzXqg4yc/J46yEc23/jHiM6EseZBMqbAX/9+7xzd4wDvAcIOS/CU8siUA
sKsF+cIdZwBAvnnUU0rwhUeebvxN03ZWl+2KMqjgQrue2Dqb2q7BmauHtIXW4apo8DeFN8TrLRBs
/ZO7+TtPnZlJYWj7uV3d6ZTpVWpB0R63x6xvw/fxgq2w5zLaNuhpKqk3KkoDVhivM0Fu7sOiBIkx
gS/kamkPXeG1Ovr5um8E8QdujwogjoYzRTslYIxgtiUSZITj43EY9v7E0ofytIoV7ub22J7MduVF
a5WCylBLj3oQEcobzaqCl1mAdkeQ7N8Ubd7suZpgAqBP4A8MWrhb5WzU4sg18ove4Hc/xgv52E3v
5oUt1k0txdZCKnVVI0LuVABj7HcnAtzlQvAUx75NbH50pvGI4czIV7EovSwIEfRnvAQk7Yoc0lNY
qvOqfTXOWQxJ542cG2j+DQpvnrhblnhI4VDw4Q01YrHNoW9mCPh7Fw6PSSWnnhu2bWb58BlLc1ay
9txtMPAbukrMp812rDWdGf53THng1bUgiJKiR1f7V71IYVb3M/tpe/qAlf9LBR/cmwz7feiJdInu
eFtoZAMnmMlhasJqBdNRdB+XBx17sUlUEH9/zsm9jHOSIl+scYowZ5QjrYLNy/G7iW9gjqAoKvpw
cvTEZEnavrSHDYeraOqBh8rRWJYeIUWiwyyWP5WKxeMOzeEDANocR6I9XEcRUFBPXD9D4DWIiQhW
bOuQCVwE6m+aOppem1IRKsEKuNtQLXth29VAb/sYb5CQrEuzgox7++k/4qQ4Fl8egZMlxRFvFrFs
Xi8qbq4ncuqyWA7dmKSh9eyWIhbv6jhHpxq9itSoY+Ivn+Jpdbteut3hPhVTQk9FvZNdqwKiEids
phvZB2vZQpZdGrQlS0Fqf/9ZqqHbBCd8aeMWO4Ys266UU3P7ffLrmDpHTpGgLVowCKsThOflJGYA
IcsWU/NEm7O4t60ABRXqjmBSJg+i62LK4jc2GC6wufbMkRqi+Ylam8zEyHXYiR7asUsyp7KWFbuh
rxoiHeFsvoxtINyj4SkGmARc4C0WHXSsRugJfgP3euVIylqqJY3wfzsatHj/gwGFK5wfsbxTxJWT
r8BzGz7DtUuD7mxqdMB3W0n/vC8fLci4LApo7z/UECVGJ8jAIu2p3ewdDhNlYfTmQmeYWETwaKS6
iCvJbAnAvqY7ZtgWDP8BIEb8INYdG371LJgfABToAfRZaGx+2kFkXPcKnnXKb0kxkSL8w2iPgAsZ
2U4nK/2fgcR2EVxn4oByY1f3K72mBJ0PE2iIiAmVI6VCBVnbdcGPC+Hlz+KKjkpI+EjeY4k7Jx3i
NkomsfLMx0FHfVKRXw3W6iyJ8JyTsmFKgbxz1+AKhbzt6AmUF4I71FjzxTrje7WQReeBFLbJcalP
GuFaDYK+Vdc8afQXCkhGSs/j0YSEL0BVOyACMdOZNO6Wmdcf6V8UfZoouOfLP2VssvT0RCz9Crql
Fl8JqDR/lwtJ1KEX4KBNfGg0xq2BFSXPUgScqpeNECvab0mNmXzm4UPt7E3Cvy9njb5k0M7Grout
rFDDNNAQJg1W5MFpUIYnHuKE2lUpyBWzxyAxp+InhTjfKVpS8D882xjFtyd/mx9sqYkDojXEBocr
J8uivkhxlIjIATKNAOHmhlJAenMnJUq5qtRGUx01lvvZw0d+WjOcoETmH8yKW2PMNjppxrDnsuWV
D1JHkQvQmilEQH1MPgN0zhN3ZNsLeb9rjIEcQsZWqqEJs04pkeebTT5KoXN652faIb4nw9Pr6A/W
kQzlFhS9aTHSX1hex5+4iSnCb79gAZEXwJaolHTnCV+6aL1sWS254+h562pjkyaOitAktssduKvY
Yk0pFHxyAfOq3k2w+oEr/E7THZHvcTnM35hh7hs8pQNedYpv7XI5q9ly1go+JV/c2XtAHsuNY7yz
FjBXW8lXy3bHlxLL5R8aTRy5G6HPAyYn31h8ARmzbWFdSmDZEamF70NLkn6yIOrcYUQQGbM/Iv7L
wt2TizG5jMZjqM2HtP92Dz7w38qtgT+WPPiqI6QVhZZtNp6W3ZTCGLzne9tj+SqGH7lT/ClsVF4z
uZpJyktMv58DPSIAMkiXRDldQb8TQRQejOXGJyg21UdMLS2L1YXJslDq8kbSj2HsBLoBhdZz2gIx
2BvDYLZrLFHUh0Y7ArzHiaX4+WqljxASNSvane3znVokfpjmjkTp5prfP4CjcR2r4eL1vLyPpDUY
1NcMz3F0NNuP4x9wV7sPIjHCyE2jI8ryYyLgGX9ijq4bCsNrOzXyNjNqfivTbCVnCeK418XdPLFR
tfCHXT9ex2BC+pHHuN13kFQ9wyyENtis/8293kucF1vxC0+wu/EzNCxbQ0XMw91sv5XCDhHDbPWy
4Wi2YIzNwRmdU2z2smhz9J5rLOyqImUH3pXGbYOhXRhFYXUNPodezS+MhOF5A+B+4Yy/NOFqR59r
IpLuJw0PdfSrVEt0ILV8Sb/DZe9r1/lUnQlH7JmeWK4a78ba+2UEXO9GrTHJij6Jj7Jwv4mQQ91S
9MCCJZvX8S7hvP8h99CCzgouQJXZPDTc1yhL1fhnbgWWdI8qvWaDobmMDsYnkHkxNbHcTAliqp0E
x90ZdDh8BiL0uDd0ewK5vNnC/hxfbP2jHoXB6z2lj8RQu6K2XoqeCjwNGL8GHob5eA0GmnH8ZS2K
i5+TP+UEFIitLoxgvdJUNxj+rmzMQ+/SIa7m/nkB2wIsoHj2rp2Y+88aaTp/sINgrqd2NuX4lr4R
HpfDYq28ht3lyJiskMkm+MrhtuvBAGrv0ULFSf2V+/fkBgpfbAXL+gPCPPSla/z9rKCGIRYVsnlV
984GT+GgH8WCnjHNnBxqCvrEt8jfsp4hFqO5ApKMbSOqPzR5JFdLm0PnmRwTzGppzMXtFcEVPoNL
yr5OJGtRY5doqzkxOqn5nc1dfwgwQpWBYmNzrk/QCTI+BBOBUKNGx8Rf07WYFUHjM7iDnuPqjj0L
Ze6xaLsYp9qDcSKbJHoDsmPdCzAvRJ3Hiy7sRsial4ZmxUZfIdrMMCKnmuioUjatLYDBtbte0HNA
q47puKI8pNLlpglGQJ/gXnDx7TAB9Ct7UZXGNRaBQfj4Mi+EVdQ88vmMcY0UWt22qF0Synw8ptP1
o3PmYnkrPAUixgOq545JnNtB6OHC96/oLPe5uryl6LnyHVi4I97LXrHtrjqRCpZy8a2iTnUdpZGa
E4E+SA/mWytbQIb1sso9VQi3bafll2+KBoJyhOvSEth+KcYdnFl+TJTcOSX2Y+YTQ8u74IATK/sK
ba/AzBvOKx+ZIpgQCXyzj/EEuMIX/Kp357ZC8vh1thNxXOQwhPhjxPdxZePaHor8neBY3qAMcbP5
4VzAowFWIO+tI3SiQNHgZ88kcaRiBvnzLIOdH1vh7pBaAFPuK9uLGGjTzdJjVykP8/4TCQnuuHkF
anhWl2q2U7gg6PP7DwMm5lvPP9MJCwCjuilBBaL+5J57NVccCk+qba6zmov97QXIz67tyA/TD30J
SfRECM9U6Cf++L4nQPkqZdTAJaMbJsEdw35g5Hu2+T0gSlT8V4AxhcUzNSlm22AWjxQJAXEfO7cx
Eiuz12p8FXBpRWqbm6RLbzx44X7QUMbKOq0mEU5S35m1RViz4Z1ePN7tMJDAC0ZB8I4X87bmar+e
Om1MCMlvPItba5Xi/WivyZ2xsya4TRNG6RalVCCZ5Tc6P8dnoyb8djtvOt9Fkf+FRY5Kt0Pu+hL5
9M/zqXAGzZt1PFvzflAGBV/PkBn68kaNBeLxAOpiuMUcGo5OlJ8+IZiXwWljxZ04YIm7jiLFGprv
GGXKzdAz3YfZy2C+az4gWE1Orzaj5+W7qUC+aeBhLK5RAPHpYYJPgXHjcGTtEg8ZGAeSIcbPnlF9
KOfcx/NiKR1F4Bhr7KM0rBv1hiXhAHd3WlJdE5vR4BhQLCdS3/sXFb+DzdJEsvRf8j9DOMukJRyh
K+DQoTZNmT2Kg00OBrsXEgsxbOHvTB6tRblrjuPWRJ/B0EZf9RDuu0Zjc0CdYEx7Kc4c+PnL9iC1
Fvgf3h5xPFLHSlzAYrAnbs7UxyxtBKy3QaVMkes3ISfgtPnINb+0CQLXFIfJDHHO+dA5/10EIi7d
FiqScw+cDHUKilwDTv8Adf8waQ4h1Ceq4kMoyn5n3R7yNrLd6dMbfDOsbwQ7m4Q9F0uVU1dD7NsP
kiE4cV3K1j2tBBbaO5kU1AQllMqH9aFprMx8tv1OI9LjA9vpYibftuOXe8vY7D5DGIYvBeWuO1y3
ChDeNgKqQsnjWSTh2W0zXvxycTQTVnqE0wlrYJHYt+6a6rJ5bZtsWylRSJ1NhwmLjy6NEEaR44bm
8emxbfQxLyFOG8Pd/QymS6aKfj9Tu+G+eAtnY0IsoUDNfG2DyU6/ZoKrPSM/CBQuO5lIOh3UggLr
/DbxFAAS/tJ9dKiv9cnWuwwPE9C0M2aIpYc8Z1kyIu9lU+vX99JZ3UD/xeZEy92KbAH8fLAiz9a5
CzlIP2I0VMQRFIgMfOLG3pOAbMUe7v1QYWnoMuVGGeJdoZ6ZRDgp9xlYe3m8IQqx75PZm1YXvQgx
3gF3AE3YQRVwef7w1QFMSq9jSz6KSEr805sVvpYH9I1oM4tVpkweYUJwai51UaZKR9lLYC6DrvZv
mFHMnp/9hvtpoFVcgx00+oc6GpziRunVs+RYBJFISRpGpz6SKpYNUmESje4x+yyOWXsqLd7d/ItO
q44Iuvwttdtwtd/HfIVhBzZR33E4Fe6bqPvUVesZG4tkgLkfQ4PiDdD3UxU6qUUckjCf182D6m3L
Hi6AWMOHIk2IfmFP4EfuzwOBLGAQzDdNbQP3VyPhu2FpG98fDaq0CHCJmpfW+K2tqOYRo0NxjFRV
ohpwiJ7oh1SYOilyugAkmX/wxO1yp2WzZlH8skI+r1GvGqPVpYqR3VA/Zpu/GSPlq15dQt3ZhH2N
OY3ZSeCqWc63Kf5fB65WFor9lelK011oq1uKlIaIHXYac6saly5LAuMUTVIVYrseHCERpt3gCjF2
W5BM67SlZNJdUixhBPov9AFBPesYGWo2DpiE0s1Rx+9SFkRu0XYI4s8NmAzekpE7UrHv7PCEenO8
LME7CqOezkfUZ0xrolD61Z1RpQDsuNBYHsz+g7BjwfpePhpxrCPYicyAO0nYIYajyIeUxwNO7+U0
MsUbfLRyd0W3iRXU7kqzeZ0r2X338EWvZ7bW2RWELrOCxDzfxxDDB31IRYb3KpMMWMj0ywkyaqwn
pHIBdeDTl7Pza3TgujJ5BAwmM63SrdvKav/oVPP3PJM6nUmTizcO8jHXWOeKa7uPC0FMnIRDLRkg
4L+KYRBjUhkOMLXRaxxDTYc55fBfwV8lbtyBlKqKLZNWgRrt20zU8I8VITUfeZe8MRTrTVShPCQr
zYdUaT9FVh+NITRtl1dy6nhtBI0DOWxQGLDou23egQfT0n5/QcWK1p7KUSYbKaozV3rcXAH8Mk0r
9VSqWEYqKsIS1i8M4sty5ZFAPqf74iWwcYl4XqhliHd96HEKkcMLSY0Nbn+5CQeuqby/jmcN/NtE
RoKTcr1xF7P1UkWhvo3BhryO7O9vRRmZ2pQcuHcNOsfYeo5If2UjnCPQH/iCf/4/nZRkeQZ2leme
eIZ7wTfdIx/xQhwOs3smwmEhfdYfBnL1R4rulKCAcR1uQJYxBN3t7PiaTxZZd4rsbTns/oAornaQ
BBdwf2rZW8wdtvHS8SQNAQNUDNorKVDp28iAujIl0U6A//b01RI7Gp3qoA0bmNam11hqYHmw0ej8
2PKtt7YED2HjLu3KGPLgZixjhSwH3Yx8+fW9SY1gsoDF8BoxbP5jvipjgYCGZDGpmEMaYJQUM0g8
f3AQ0AFsGZWynGMh1qayDWfgTwOMgTJifv7jS+5qE+f2OPVHJdkdBL5iDHcSMESrN6kRc3XtNiGy
o9zbXqQ8uV3jzwXahR2CGorlv3gcLIpw5I3FeKVoeeoX6rcItBi0aJDZFuesa043c5zgA2hUe/c+
q2lMNunrcPo2MvarnBU3Q/lYVf5SIGmXKeq07eVlJ3Wk+Rjc4nuPhPzBJ72IyXTFNk3LQ3K5WczH
uSzLm9kQiFrDykttHIPonueOwcqq+ITnz4R/L3Goigc4/3AyQwAbH+7c9OuToVjUMj4oC1yttgFq
HICMAndO6ZRpTkVZEq54yTXMftJJA7bywBlQBt8lmfCRwRkBSGW4mWCeBcBwGglwo08cMh2Sq6AN
rchCb+txk0lO+Ng3axI+QErADANGDB0bo1MfeLO973pimrPJml+4OyuLS/VrFrvzzaVrwsq8kddt
24JTTDInTgcZmoPa62OzgHoqnz/6ZmYFZ4LVSe5I7VFrO8qXuLAE1ZuvU33lGSsGiP8qUa7vOnif
T4tar6WNVuSuKsflEu220QhVuAJMQcqwlcb2xtSVFDRvGqFksZqME56xyXhaXqoWXHZNgof2QcBO
h+0B5QskQGJp/sZjOhpHHLPQeUWJhNPNeoXh50Y3geZH1OmEGfVkPYCdnnBMyAtQ7Xa95fnFPi53
BE3k9pOUs962Ad5BAnP6A61xenSNeZD5/ig6fzautUs1kxcbaA9pRtD7RwNGgK4fDY31JMESHoiY
mnKjmL/T0y/jZ5HfhS96RpukDzKVhWj/FLZEbSOMSkSySrN3J13h/SMtpPoCX+PR1appBAd0IXX8
envcAVlKLwjAJ7ZbKUyXEbNDEdXcN06/SwJo5+KywCcYPPJekbotqRFhVnUuoy1PNVwfmLSvNvMM
DoS2zm4LDRl0R43MPsRvBZLWQr7BMLB4w6zHxUHfSAUWDkKR81noy/jsuXlNslsOZhX8crqD4Htj
cIySNQEPLA05ya4qdnRKpy48pI9Xl3gCbxT3UAc8CjjrTL7Y4ufwl0NVDX1FaRizMLP1w0IXgtnI
qap3ZNL06XoM9n/RaBCAy1Nj2LQr8qGi8Jwhsihgfl0wmLsx0zTOSHsTFhXIAgJ5InCaFAaUeV1H
OL0dV2kaGQj99wCep6JbUxA2qSTNSpE1TndMv3jlP/nqPbDYE4OtLJTOfdVet9e78iayJEHkSOJo
5IHiV7usdjDP4siaVX1yxvnYgzenWslYo1bCwyx2/ti0EwPVAxdAOF0SPhWZl+/9IWNXRzVkzlqK
FF7aDbibCNiNQ41Fw1qq+Yfzc5wWpu86+Cxy950TYJp3WWLRW1uPQtZx2qMjVh3TlM66oFDuEHxY
EMtqPfkGfAotKw5E79lXe53SzTb8uHHZ5oWPpMVCCl0s9dn1IjTYiizAa39fbot1KvRiZIAU+i1h
aQGNBCJNyxPMhg4Gg3rpOMRiD4SnV0d3GSLEFUg8l05fEktgMUsgQUlQKiL0dV8po6N1CZQ2138l
RuefSL1z5ZapETHbIOQ0WoAHxRKHXvJd5/KW0bjM6nT7UelbssAScnPBRoDzr1mCsJM3t6E5TI7p
nuTslX2OBKQ19yXjJvVQz4ItXEp6MHu8RdorB+UAUb2vAvX65ZM9gjE1sDh1EPpm6nGcMtm3uDiD
Jzp+cPIp4kVaTPh/cD4AzFfn0dTeTP1AZh8R5GHH2EvYpdrmpKeP1aTXmSfpHQMs3CF23J4C8+zE
96nDkBIKtq32KYicepTyMN8zQXcDWeqSgO+4vN/jct13qe5r3R4eDwONCGwJheQsRXEIJp0o2HWe
uRtx8DzpPC/ddqVPVIpZKVRjWY4HbpJYzlfiAYM+WGY/yEhaLCWiwAcJ5TDxemKKhqz/alzt3MaY
hXZCUz7O5/5wAN0GYt3ylxX5UTIj6geNQCljqbGBkZiKXdPa/2XgklwUgz9ggdOLO0DkvGtXF3Zp
LO/kUZisthLWLsI7XzywFOA98CaIPicdFwNK02lWJjlIWrlD4noO5G5eO2a6/3d9i31PnDsPZQV6
6zHeATLqQNi2tPZJzTUGamxS2SCjrfccJIeexPKANcBqpbCV4zWr0KmQeJGDpoh4RmGMuiaeTB/J
S0xEYkhPXJLCqfRpzF03h6iJBk10dDZCjaCru3Iis/YT/iDAYYOK2CNPlYbwVsTvchAVhT4iy/28
Y2joT9PSH3o34ka8yGZeWe6wTaGn67lp+Vwz0iJJ9FmSTJL1a+zy9QoGNJEESPdaOpPEEElO53SJ
ir2mGLscK0OTn5bkIdaWKkhh8Z7WEnR4QYTRJwIvw/5KkoKhjrqEyB20do7LuHUQwaDPKpi+BNAd
7i/CM2+xTNzN870eQnEuLveyJDPgiIVEUCsdysDbit48KM00JlNOSOhvtHHwPUl71NKO+1TQBC3N
tnVJXf3HKqkdorVJ3qdF/lj2bh6uV89H9zM/gmdyy3isGZsfA6lCSVWXvtl7RjzzE3wVJHHy8oLi
Dley9PbWuw5VhAQGNTiUJgAGVpAR6WtPmUUiBa3pz74Kpe59xY0Ywv1cPTAxXzsd2h3fGspiqBzR
wL6hWgd1SbbP0933Fn7ZjDStL+iAZQX6TficDt6nXhJ0+vZWuwuVdtjRf+ofkFcPoNrY/cVD+fzB
ScuFch6RQQtrlIRosrqFxb1GX/oApMlfGrawpVVwBL/dYbdeOGHEPEyLt6a09Epg/4Ha7AId6inV
0IK1yfo0Ztw5LjhXHJNlBghZLvNLf4w3+dLdorLWMr8NGg+SNyrj37RecVzB4DQNKhwDXducqytz
KgeigHFgxcrulDCMzK8Y0XJFZKlVY9VvEb3gFrB/w6moEufL7tlCGhbh7u0kBvWSDZ0FZeJ5tZVg
BSQqy9F3n1l/uqN6lBjcEza0xB/6+AuOSqFwsr8UCDkCI8wNP9rTSg/HVDYgDEcqp0x7NI/sr9P5
Bdgeogn8LaHZsbOVy6j4L64L8pEDO0cXIu+4+bRXzwBuUl1y0D4wVQD2XeDFjNRjCVIUZM2M7AAn
FQYlar7QykllvoSfsjlzHy926BZ00UAjfXDsrGafDHDDiQQE0fpVmC/ZEp1iGqOvYz3ZFqnhsQas
+myP0ayqcvNbeUIhFBU/vxJip4G5WfOd+cqe0oT/cAG85dF1b030r5nhK/bCJRV8yHTu8ZwqEQHs
+fJaezOiXdm7YUJgvOwgacn8dk7FtofdKhH36wREO8INNh138mg5lK+baTIxsMZ2cfQNrH4rZR77
vuvuNN27/FRn7GWOnSBjb3D4IDtFMZ6dwRnJ+lUzUNWzITe5z1bbsxz0httj2PsxxxfkAx8K9ZcL
WHPwbbaw5nTWUPUDh1EIL23F8wXtw+KWaXgZ6N7yPHUCETv6jwHn9gBtrWU+zh7WwDfPxap+1PGR
rwcw5S3tJspjLbleeXNL+4yWS54ip4Ix+tXKx8/e/HgCZDLXyRpZrenRE4FHZnAVzwLXVshwBXcW
O3F9OLfmQiCf1vXmz9zsMkvBAslkEsJRSeD1Apj2uLtXaDZ5RZ9GBygQ1s6cs/7yPrLQ2c6HTCC7
gweNNFk9b0LK0mLdyX5SC4ZL18xMEd1sIIe+Z1xLDUiSkkodCAM+5vbLlr2QpoJ5YTHEehx5z2wK
U3BP2K/RAn3qtytDymRYr9bh5bKDYE8lfwR6RGiR5mgMf4XZin2AXeC46q08Yap4uYCnI6Ed24Gd
e/68opCJwrOQ6roI4Nu1UnZ6kX48tLEAGPLaP3F20pJIC6xda+hErmU8ZADWGTCA5KqjnLyTc1Ld
GlSbSWTT6IJJUX5pEHzhdCDnHTEFdlYnCI5XB3UAveOlRXfNLhiIurvhqfaQZi48zOlEU3MmChme
ZnLql8m3sEyTkqHF7Kny68LCGjh6WQ3cvAWqVYgzf3wL/HlmAVtrOYGOIoBkUbBYADvS0qw/HNMF
ioOzONRkM2vpQS6Ph8KBkLG9Xlr1a9DMKXNU9rDc+PHCd8bT1ZvY+vxChrVWLBpzjVhHXFHRr4i6
b+EeJpTnWiyFkmP5XCrTCOiZftlYxnwA0KifZLbGw9Lqbp5oROjtAKFceUDXkxFxtnfR5ANRPsGl
+zgihcBnLhSV9m4ZCC8x9VQRpfo+BKyUTsi5B+IHD+jKCvVxmd9tTLuHDHjV+heIse+F78+Wg9uj
L7q65LTvOoCB16wrsheeWxqgeUiLFVPYRw9ccp2lohHM74/ZMbY1zrAs8U8jSBQCOt8m4AoxyiP2
GEQR4GGXxc39frMrGU2og2byCUGLOIvwmxH+nUaTm4+SYesezy+ZphO3cG+FHJ9Sjo4QRGnQqW95
8JsUhULFE10+altwyQmKo2fhC2fNYmdR7fJgKOQuv2yquWSBvjZ/gzia5B3TMVlB8jVumN4hnnL9
Dnvsd60/fnQ8HH4nQNIER28WGqPGGYhQCsURxA39pqhI+2j9OgjgFBUm+yuUpkxCJM8GoWiVgT4a
NdPIxeBL/e1shxBremXtGCNc9pg3B5CqgnJdt0BoGwHiVm7tFjxRi0abhg7evEDQiBK26LpXirHB
+vhz2eB7OjTQmFlIA/5BAdG0R6Vot1ku7Y+83lVVvX7NDHRUuBXuEQXbNRfCAH5ZdbRJ4slvENDB
bFxcmhk1ClK8CusE1EcLlNTPbo21Pz7g8WfJbxgDuBG/Vnf/fbLxcS/tfpBclCQbUcKp40035OLm
nnjB6TWwAWcjywtoiMQy81Z/++qgeoWaCGi6O2nXk0zORr5TR3pHb7LnqyiecGSyBhGw64Vi2DZR
IG2vu6901st0/Q24z8SE9IAf7I9v8WtcUuVUCMTDzlpv9/CkfKayaZLBbm07tEQEex560FVU9VpH
FFGobyfIGelmve1IazYVZa9CIaGPQbXg4gGbij/z+kJ/J1UOn51HDOV+xy176pKeL/LbrQKNygN3
B9nDvq/KQQvPQGweHteZjGo0qMftzaV1V0O2oVnL37L9wPv/uV1XNr7rIXlYSYQAFCTUjR0bQQI/
fmQldMegsD5JsvwGLWwH7m12m0d707ivgAGd04rJeK5HXVtdqE/qSfXrZSzB7gr7+lyF1t+xEI0p
ype8HEvmZb4cK/b3lyQssl7qCjbpAhn70QixRT8ydVeWb0A9XmFWOqqiZH+UZ3CMO/aAGNwNhxJ/
uPP53U2jaPXZAN0yHXk/MLCf1vIOzas1/VXdXDA1DgQ2gJV5OwT1oFXgzXtGxfq4ZVJyb54pT8x6
EqP6wF7RKCZTbeiKz10BswLfIL0zKqajsYA9jX9gyJdHBljkgKbnxTjaLyH0XETMiQTt4of8ji4D
aw7IkrHjr/Gpd7bvsyQKky+kOrejcexs69VZxvE4SeZFiH87zy4fE2gI76qnrH5ZsLAnLKUQM4pj
W7bKL3xA/3oQ0PULnBLfyew/NkaQRVU7jZyqEwpIutpscVPt7HTyG85aJ8Wt6G6YQJhF1Rncs3oG
NVKtvLiJHh8nwMb2LKo0oviCOLDuztRjWp97in4TOxh16ePu+ay4u4h1+cpN3Mkr3wxy8Vp2IWIW
AsSfQO/YyjDk318qNR2VmVDpAhYlHMrvc+HLtSZcXGs7xvJiEzkZbE8CpfJCN6mbEIntfr7Zv07h
0Y5Cx0jRrqRBdVNf5XSxQ0OCjcoxV8eTFVA5qKT/qOR+5AYkKNw6kNmm0S2GKmya+5GTbdqhMakW
xDQvu7HkMaCTd/Ap5svKZbuIWDfnRcnSy6yjqZYEslWpcZQPSnvLdQSf9aft1GMBIRJQ+9n7Cyt/
T9Fic8CZrmYCqeetACzlGh0EZssgagAJt6pZzyRlhNJEwUsECfQ/LBhSKs6i8eNE9emP10SRbk4c
vsJzYBsGjRXPc+pknDFZpH26LoE1jG8P58AgBp5bQR7GqE7PCv+mgL2l/JEO4umg3HhMtfTrtfDa
g6uIozAZscCJ7tSpL6Sedgt6LHmAA/Kgm407CNDvL3IL7E11E4oaCkH1OXTFo1yMxUclL9T4XR6g
liPSxasqGQYWfIMNf1q1/PKlqW1qruArlt74/euCSxZQOOV++dFm3POOD+TlQNaep2zs9pO1Kpg5
j6ownVCGxdpnEJxXC29snlNQKCM99RSK14/ErtR9+NFR7FsmQHjNftPysSOx3PvopsxlKvNAipNf
797i5RbQsLGOBz+GGCRWJWeIvSMAuaBBrzOsIXsnBC/PnY0T5ONVDE+tzVMLQmgBFcWSzm28lQ0W
KUtD6VBMjNojSL5TZRaA74+l3BwOs4SS7dDGrfsQbUJLNgvD1SGOXvEXMU4RF5OmLwJcty9A9qb9
bQwIrZ2mEhAe1A0GM/JqYg3W8m2blg8CWtryvSc5qx4BwMbPxtTD+h8yJiZ4KkxsU/6kQfFf0Kz9
96H9io2urb3wRymDRIcPodAD+Le5l8DURD09slFcpjeIVAjXxOkFD2yOnNWiO2SVFKcHJIARugKM
6BOd2e5B9ZgbQ0bV9Fmqel5RBdGQ3jOTjdAi/Egh9H0fPJ5qSeEEj1ZnPNj+xiDDeb97CuHkk4k2
QEwkE4QEpPW8vn1FPpKQDUokrTpXz5fKYxFLzYX1gHtEG4WiuuSRGwzlUVJCxBDMMULGGqH6M4vO
cM5bez8JTN6wwzy5Ml/dxpe1UvZ1pddKbuLsslR0suDch1ZLrNpoYKt+s8+u4WWz/L92VGRW6zXx
ieIcG5jMZh5xQKnrYBRgZ6r6iW29jS1xP/0mNCqbUgI9+yt1++Ur0sN9wig35vAJe6ObJwdcAuzo
wFTKf2VadC0uZvywTpSZKfHlx3O6dyKvjGaeDjxhngFmLjSKpxf0RNN8srvMJ4zKcLllU1QXYbFd
aT9bPBuLpQkmC2FaS62Mhetr7cZDr2ALCxAeoaLQIz3qgTifMl3WMGeLwAES9eVPjLrGmHUktpY9
jSIsIoYXTH2Mvo5bvdbhvZ/nMwgFrlah2MPQqIHRW+JCrHh9n+RUF5y/PQP7BINv5c93L3mTkIpF
GZNhtVGeGiGYojXJPlhfmYMcapIWtCcNlgOzYRVtH4LjyyISgwNyCiRLcuGMzYKRnZAm2cKMz3HV
FmZcrjQr2X1iWWaLD+mFEcoY+dN2NKtIv5ImAdf8f0bKzy8GyilllsChB8sUBcMDSr+/l4WJvAL2
IVIaTSE2P78ZteEhgL3rGDOPE/wxX6BeRQZIR/A0PqOPSOTiJUvSEWPft2yprvGF9aSjm3L9GUv0
fUEzzH5NjeS+pTJxs4qIcKxRDLaIYRcqLJVUnX57ni+uFaO+QK81YN2YnAiXUU2qMznqzootnXQV
8Y3F3FdqsgZ3UoYaK2glchFADH323fkj4E6DmzcZS73Cy+vv9RBVgPcQhmQNaTpC1aBxnSSxXtm2
F3hrlnS+i7NdXhWBtzCmk9Bvlk8nlIAeftKgNoqqOcwRJGplGs1x+aFvl6zJPUD7JPJ46bJJNApz
YSsx5j3SKFEhM+EferTjiEA884+mw304zk9esP2ABg5aHhLaYEFx66ISE+UyxmxbKBSf2FkmoWWb
QEe9UJWhbr2q6JbBfc3BwwLk7GI1WOegWScy/3+tHPuSc1Cifv62q7AiaEo0MXWenn5bgKtt5rf3
K7s1XES4J+c2aqUBOuFyVu8tQ8Fs70khfWLAAkFKmpsMsdXkfZ4OOhmzA1u4WQQqCkItqjDg+CqA
Je0PS0OXHC1Q9KA2ulEhq1sOjUwdv6pQYGezzVt7NArRHqvJFLqNMaSc0VBQA9W7uki+9CRfcfLv
sC7gZi3FEkhkl0hYgzghGuCBr+rq3Jy3urvpvkH5lXgGl5SVXYd6lz+UHvFI+VhJw7FYOJrt/6CZ
zHGhj99pcNbv9lvBo8Brmrh4qh4sQ4ZlLW9QxCsaZ//kZU27nBHBX94PHcCMh3C5aoevaJ+DA4gv
QhoS7VROPQawAfR278A0P6jDw8Q7BW6P4EQIeHX9udkWeqmCUcD4Qsw9Ny3vWPGtV41gww3+h9su
pkl+4bZmDut/qZwk20DBZ16fBNH8mWXFynxBjmQU9Sjarw7Eea2cTOoALOrBOaFvz0/03bMd/mnC
H7PXr6ffIGzR9j60Nr/liV5FolgCivTOJny+TaTEHk9rfnPibUXU1hSm3XZ+mRKAfXwO0akreRcT
S7XBV2N26n648w1Ze4bgn32FOLr2NyP45ep0yvo+UCyy3RHkCS0Vvk5CN/unx9m+9C5krct3464K
CppKYTzkmr1ZRN6uYwzy/u3xqK8DPSnnZFhASuaVP0gmAb/iJCiSBsSYHmnj6JiKskUqWGCLDD7m
siJrB3JODyVQ+mSDtk+B+Af5e+DnZUC7udOpYOo/wq/3LRp6eLYb1TG4QoEqibYqvwWZnPHffVz3
FR0f8ADl0jQbkHq+8qELpf5+hQajhuMUvxYI+EHx5RX87FObsVGB0s2lBaGWXS5tksfjzuCy5E63
f0XOOyBPD1MzscVUD/XyEACAj06k+S8Kf8t3QnjEGs/H1NJ18e6fGK7QipHTF6s/A/r3LCbI52m+
K4elMKszShVwlO1fEnVucXYyM7W2FnKnAgbfh5x10MpBOq/UjVe+EcNbUNi4ZsCxXgoVI/h7fzX0
g/YypRyZsIfF3IiodeDjUbMDBpsSncN+ipDfcU6ywZ+u+/k8wpcp515ZyzqFHX/k2K4iT1cQUmcM
3pJs1BxHeXrTgDWHqljMkiGIx2ftG2GQLuesH+o5l5ZbAuhaBZyP3BjzrY9EZ8V2BLekDFH1Pogo
JW15y3PUyqePbEEVp58GabGllUx2UZHkCEMNnb9AiS++UOke14D/h6OJ8jwpToARblTdoN+Qnt+K
sbBbuK/c97ACSeg7eelY9m5imgSUHjpML/A1ZFaf7VHpS+aZOgrxpz+qozqg1/Ee5PB4RoEgO3gP
QDQWbMhguROTYi5eted/Kylnn7rT1cUDNyLyQuiLwGa6/jBaEkZ1BLVOkumk0/JAYWpWsewIdE1g
zZ1ymnvrgj2vJ9L607m3NPWYaPMwfq6unpWSl58C01zUWn83iy2x84NAhkQNXJC8xYCj3/AfW8FM
RgrM0aQX8y4VgN3v5sE/KX0kYv6qcg4ZwKjxRmFyl5lkUIFGGoZIjH82Fw7gP8dPcm+lr5feYK6Q
zgQSKwZxXrSCr07f5R5calKNK5JXaKOcQn2lnwniWLYDxggopiHIZxh6qRT0YMAFlNIcSuA3m6tT
rBMR2n24ENqdX8GQOLZ3xjTmrXaIQgyHbpZRGjYHmQfIRvBMeqlnqctE04XHr0Cp+exI12JnsQ/p
xFrGPbENSwxNmjjcIFGfokq0GWCSh0OvcATsdps+z3NjN470lBB9ZqRplLRYFPJDwK5eJDT90uQS
RoBjHZb/GVpsjwYhDG0yg3TOxpgYaz/lWrrGbXZMMReJpHT0A85YIA61eYPkNIvVupdZqfN3Ocs9
s3ZnoZURPm3NppwGPciAAjXIu/sxYkQvkdH8u5NludQCzGwQWPGHM9A0zosi9gsxFKzrqSw83wBX
kdDbCS66pkWKha4codCM28iwI3P93A6JgTt2Rw4ABQHsgp+Mpa4IQqQqTt17pFq89Pfk21TXAk76
09yKhDjXXkS1T1Um6rHypvxhUkDFzyCiuDWw38IZ5L7Ap1VV9UtQGWBHiQIBG4iU/ZRmg1IkMpiZ
1hSEnd7W96in77cOwHOphyLoPLSKpVBBNlEr2fKbaNqXxMdOniSZ7NAnsL50keTbXrDwDIj48E/H
FvATPPTd6rsVM4+Qj3uldprUde1iYDywHss6llim+Kn/q6J816Ie41XOF+5cNlFtDHGv6EPZ8LgN
vacdKlFqQA6BwK1vhEihwlQUPejXgZX27Wy1ivT6ZtBEFOi/71xHoR0QJbF24qvjlkiSpqtDsFhA
QqjeXSQeHqZrAirAlfU+vvs9nR8VTy2IEHobCDg8fwCT+LkOHOyFj0YVRHhvkbrbqXFWqtzY3Tuy
HWbdmNwzCmyRis//FwtBo14WfO7IQWHu7r4ewf5Nd07bBCwvZwn6EkPF4Boi1X7HXXkitkxpanvq
r06YtnrkuVzmi5+VgyATnaQugaKOAn+Xq1iIcnWhU++iAQUjYBipYExljUsyK1wwygtHB1tDz3hk
THOP7M79pZHR0lM/wCH3nAumvz3i/fHB3Sa1KDnLu03ethxAXJacr7uQ0P/LnKpFfB7/V4dGEkdS
zZ9wtE2ZGH70Q7bvmU2g0xHqhF1tF6EcHa+TU5CjR2iHu5RFZCT6b+3nRCgUUEX2GjfVG1ycXpho
O6YXyRzVfY5CLoc3gs08ooNaYjm74YekXgx+miOnkEAc8OIJgDwKecK38IIuo3wbilkAziv+WvcY
fo/JNchaMNGIqkkaS4tLTPRnkorZ+EgSEfpcalxmYiTlskc4X9efZ9qn4SwQgPeNY41wK/F7b04o
rXXkM1GjiylAteYvAROGbsyyzgbEMJTuI3jv7CId7Tlmd0PwtVWfSIYHG9jN9kmxU9X1VYCnY0Eg
tM6uK80jDzwbI+1zoua8JO9jG8QTHzA1ENS6hixlKko5pXk21wU7W7N939w+Hyl1FIhBtXmCq+F6
PbM37++SpVzmjs9ygGOyuBufEkV/HDtNQX602WDg8SPf4l6nH1IDiZ9On/OM3bCgV6tmqcJuTj9z
pSCXxL5B1pK36Gs0D5dJ6jKoiZ5lYqb64/BQNT1G0QmX4rv41ihurUdib66AiQMEDBYd1kirpvHT
hn6y1+K3/1OLeGNjFsehYcpzSGvd4kNwnJqaxOAgLU9QLllYH+FWBzerJLYacGNbF4EWNjU08TjC
mGOIZVv6Gjc9SmOJ0xAI/WoKgWb0wqorZzYUfQKf9BSnwwQtgU6Wi1OaSK8frvx2+pElU9kbcM9k
JFEx6Fo7UqJRtWNdgk43vk6j62taVBMl2z96Szzq6KrcZ95jOI73w3p9DZ2aH+yKDfiVoggubWGh
DYiz4H3aLfv6WlEhHtu0haOW6uLiJ40GFWEcVCRQzUU+c5huYOMxlT3t8qIWhQA4RnYHZt9Rxl3g
9lOajrp3JlXrgIRQo4Lx/nNmiZ0XAMn3vNixEuUd8wYrFvf5e2erKyTAa+TwwyjWNmH9oHvSt7ri
A2RI40/7vAovdXuIw7Lgu3DALFVc1GtQjDEdFf/04gWC4vDB6HMYOr0laI0Y2goMEzCChvZ03W7Y
YZME0LvgMbMKlWYNWY04VRHx9tNlONQA050Talu7VtyEUtdGUgnUot8Qq9KjaLbj1ONYGatdsvgR
e0IOW4AjaapRDV9XZT53scMc9BSWSXZRUegnkNCdVfUpoEgNxNw0fjTAWZ3Bx2Ey+cbSxwMMOE2p
kvcqYjF1ZT2P5R6uYb3qrQEKXdUKGAOyYyBq/L7OZWvhfyKepLnRO/3jvO0x9qt6ptqDfIuFtNmw
wbb5orC3NtBdZWyi5lUiDvnOVR60cS34rrfUbMDOuLy4avSHE1Y/uxAYNolvRUtlQXfwEhmsx+y4
COsu6dwCLexUIicueztfVfcJBztFQcdYEnOkqbtrmoGl565vxdjMXtTAnKUBav7xixPSMO2mAnPu
B1RH3mdD1W2Bv3NYgg0x61h85YhZManiEYH9t2Y0hB4Z/cMshUR3eQvkJLQ0touyXVdI3Vd7Gz2K
wWIkgZxIboopiw6wdYfHMBw4OcYKxVZlGk2YQF01cezepj14SVRPxIYGbvqAci472TC4n6ybsc7I
lsOAeLJle5H8gOCBBSOSrXdGAaAutV9zUn6qGAG8zKXtqoVeA9IBsi/T2/AUdt0k3KsXNyWNQ+tS
14uKAe86IhEgZtYEZxIQ2RLB/n6Xdv8HlhoY6U1CJVMHUwPE4QdFkIF5Smq9sk3l/TMojwCZnA0X
PzUznM0mtpBALsbF3wXTy+diQqDWv7Fe96ai0OauwvwUOhF1rKy5UHmFPOjF/IWTAcVWOmCTDZrm
ZVcDWX3zYMMslOyNFJSru9rb/hdvFpEj4QGvNVkCdMlvXykWL+R+igGXkZsYIbSjMVEDpIvSbRvf
JrNGh4AxSfeRahLY9S6VrlnuR2/DqrzAaBkfGMVWq2ccY+dAyS9rMNxDhBV3VPtBEVwJxCS0NSS/
fl2joS2nlwx/SUxSnkcJ8SBbGkEEq0JE6feGK/4prkPSr/75ewxFDO7dSFm+ZOZ3SJEQvfJso5Il
3x/5gg2Hk+PDM6hZyCARzUpCnIi4CK53Kfr9b7aGN45frp40VqEH/p/IefGb0gyeWrBlNIaFZlyr
0JLg4ARzbJ6fHQofFU/hAGH+abdnSHibQT+wxdwo4mQbLVmR3iPtZWENkgMDCeeJaTI6B5kqMTMy
2qByS+D4Q7luwQSxOfJPbFvCHLYXRUxk0W/dPD/I6U5AToj2MOik5sPrFXRfqQyJT9K71NWrRO7b
OoPVvbIQpAXjpHra7ft2fZg96xAHR4poeHhc6O04g6N+ObZyaKz7qyRZhOvoKKTaQi1cb5/FyFqE
u3MVP3ZG8tdJHQvd9z69/OD5wiuuWhga8jp68yDc4uj85b8mziCHV8zz4v/Ba1corTelQgSrgUQ/
9woFE4ATzXQW8wQrBhqG/HiW+EKYGo9wh6TCrFDKzcPdsO8kdk1XUGzyuSGRHhtp+tPolaaPA+5O
Urlgxquq2NJD1PznVPpmtkut0Qw16La4OTasveFBzt+mPSUtStobBzVq9mtPq55QGWHhrTFboHmL
GBqMC5/rbbOmOI4gBs31xysgB7V+SehB7NFcq2+52pr85+qbpIcgmqZdqL7kHWtZEEUDfG55WSey
g+TWeFhuLCL1wB2PdedMkbKU60w+7nA+CUBq0Og/QlbX2c17iXoJno7EH6B3MpogMBw88fKmKqiY
ne7wrc2VFwEJ4aeyBZjjXhl27G+RY17Ey2viCCtlJVz2ixAlmQc3biGEIXUgBb3V3zYFsPXyOfZq
MbTSkPRUuorzRhzxzrJtexUBleufxvoKezRADt+BeeRzFf7GcHp7IKBHtc4gdUgMj7NdM+hZniHD
Y3tnDf9/+r5+rGRgUhSF3zylUKfw+S5iq3U/764dXdvfsy+U0YhSLxIWo0lITBtRVdGacN+m9mZD
mSdk1rttb2cmR8ELWHjJqTSZUkt1OuWlVwDL0OOMmMq4oORm1EYaNko3rwXxmAy9Co8YHaHuQtFB
LR0TY15GVhLTVnBaxh/gbyuJZn1haC3NrH9dNY9z2zzr8Mf9XNBNixoglGLp+u+AEwA9xdJfLcea
aIxuBtWBT46G/Y6cxJGWhk7EJWuJow4nbNolHrIOgKaov9Gnp9Rbqj2uhsgttm6t0tyoBoAQYJK3
ILas+4jX+BjXV+iAc+Lmzvfv1hVsDQBot4KH0pot5gDLsqdXXUCHyvjbjuucDMNe6FJvkBUeIMnf
S53PUCKPaZsncYUvhoPBxxGG2rY20LTb3uy9XfVqYOO/Yx3fLffWHepO4iL1m35qnbox8MjPTXYu
xsGX4yYc9VkcAqQJctmuq+TQYiKi69fPnYDc/TSLC3Cle2uYCYIGiOmsobEII9BmQI2QUyk+4+u1
1ft/9c1YCmp+TAM6rdNfTY6tv/jg/pOD0mPR7BlvXRs20wUE3ojF8RriuV/GjsnQ/RqpeWXDd/lX
/t73h9AX+JoKiJpNPiqcybFy5HgHrR/Ev4Qz4QLg9ZXhFbf34vkGN9tOs16lgulciCyuhvbJkqzR
GtV5nbR1OMwxYIgcDv+4S6XV3kozXmPotMfY249A/Ij+JPZ6OQFCk/UtRIy0T/3P81r4JXUV3Pta
lTBVBvGvdJ74R83Z88TnmDF9leDSjqbbiDWoVkUAOF/d++0N3FjVv8J5WJ5ThjftKG3SLhlmpFXS
q7hQL+G2ngUW7uaJPPe+ULDpkUMZYCfgNsYW+1e/fJpZStpjxOgqFOcyadARqvvT9Z8GD7Xj0+xP
ig2I+Bc8zWCDcp5mEmvJwiqisCMTHB5XKBm9gxW9mdsZ802sTzBjxvvHp245i2PGitDF9sBIz8KM
20TcGJm3RlJxRNu5k0sCyxfrOFXptnhnffnrTfLzXd8fnAFe60q2EjyM3Nigej0H1LEh23IdR8Dm
/J/+XFD5YVAS9MJux346/puuFvIOXb7e6dnUrRrIFwn7Z0VuUUiM4wBrWgwRRl38BsF3oETIc5dL
IRtYn9UeG0pzBIX1L4RR6EVLF0tkfgIF2keaGokRYWdJkenSJk6cJPTqxqgS+JSRHLHegph6M6ni
2lpNLasOEAscJ4/O7xXC7NPVlvMkzUxi0WoRM1olQSaxBeVKEbgiY1YamC7VUYF0IwkATskCeTlP
J+2XE+4znjqmtcC3RhPBvMUShh0Y+GZVkA1EkyBd3ZevKg3XwdihjOEquVmQ177/5O7F7jxgaQB6
GRvLOqAbcG5SzVaSrRv8C7zwWgAErLAHfaWPEoGcFPBHWhHCCnCrWWAu9CIvZfWCxQfemL4IBvep
kc9IPXaq+5HnM6QIUv7y5P4kbFDqAfYxk8lolKaRLngqO24+zZyCErwrHv9SucH3nQAYwzi7tLlY
zFGiV0VBOsS39WdQuty8/vjo0rmyv+WrtMp058nXFfTxeeG6BibvZW8m9DBQhXMd+IqwcnbVrSPp
q33S6Z2mHUR09jRdv535mqVtzWeTNL5cLPSTK//OjkB5vLWdVWPzgoiqqpP9QTqHfE1Dl9AWpJiM
V/fruQTMgWb67MSvgPct9f/9uZ93q2/nbHScl5GirRzGySM2vWHN4yXpvYQ5jkdNlh06RL7WzJ9v
N1EiApzSki9/WfO1DzQsyyonpY7wDJW7qsbb6aPM54e13ylh66cSDYQGJgbDdVpXMJBijnQL0SEh
GEWply6ANyoOOrJjs+aU4dhGmtK5e9cZI7kocIf1enQGgHPvmt6QWZXmrIA4wN/7zshS3ab4Wixf
Eh3CCdG7mNzJAiZCY6lyaLrBdMcrtEwrUq0CR+PrlqwRaFGR1E4Wc2briRiM+62veSzots5qFj8m
JDis2osGpozyDxSRhhmW7NP+EYhhQbiYgHKASnNXLUi9dQQrqO6Zt67D2T6fMlquu8TGryNW8cgl
cgE12EaEJ9Vwg/qMQJaAuPMdFuENintpt/Nr54yJ+XTS2Inz5ppoaTMl4pcsBIpRdPexWJz/Mxs6
ZY6v07dwiOFID/J9gWb8pMbiOkdzRAvm/c7PNz/d9h2mSHUYVTjK3plDdRE4JBAMPf5P4GXGrIZv
pdu13dIuSsH1SxgZhZTz+fGAJ9wTzNyC/5Cwagr2nMXtF1/N0cfhpREys6/5m27wkWcP8PJx+fNU
M02cl8M7D1iFdMRe3kJJrcLWk8jCs8ksUvz3yTQS7sGUIBrgkowSrDIbST1Xa6vi7+dRiU68udmI
a6Ww4fte+UTyIhsMZRMTfs2zTSweSQ/s1ydcKTqxZ9LfUmoQABKuJL/L7HZGgfppRdQ5ckdvuo2O
7nDsMj2IQ28ksPvNeoAadWN80yGAeSYTMf1/K6kbXoAfdOXOlEt3shn9mwSbwJ+RElgbyUqGepMx
LCmUEorJ3vj+xfsPARH93HAgLAP5z+4XedlX8A/TVbehGtezStXbBWFv9QGOjbIPx4Y+Q2/qRYQi
+jGVNCfgKQGcx6VGrJtYGMqIMAp1oCXdwVn6hDYlZePt185aZZN/DXzQQ7kAOrmJzFrLFK6WQTnC
gRjoUI37KyD1tT7LOfFw+vWzygIfaAFRTpWV9CillOLNgwPPGYreNfxqa+Z9DdwlgVbWIgeSww2F
pbEngUwrCBN3TPnQJywGa8Ojn7ci1+8MBjGyoErc78UteAtpUmGa/eauEz9+Z+cTbUGm6ErI8MMp
kcGOZWj5trSIkD4cHSMt/HQGvrC4ZywxfVZRt92meRzS7bMlvKFslNgbZt1KEhj8Cy4uPjt6bl9s
8kc0st5Ev0WEUFe+va2nO9n3zqEzTnV69qiijUp6JGWjLNFIBneGcipPHZW2rVwtbDHPGWdDxxoE
gnCszkS1Egw+Rw5qu7aaRG3Xrwpe+cD4vl7/zvLYd1wgFH8U4Ao1aGQmCDLctb9zUnw5gS4q/T1S
Jdjlo9i5TUeS1lYdPhJCx3VQ1aoXMdkedfZRwUqlHn8vInP2ITGCtPS01ry47DRrV+fo8PUSwn04
vFiDCkQd2NCFDp+ISM7OmoKUhWIH7U4haVGlXuPAtUT1vYVfXqvdNi9FqDP/T0l85tceLSu13unL
i7AXUPicZ/yjN6lV9mMfJS9/dBmMHreTVPo7EhekHTedbdB4xLfb+YTslYbWkALPZlsw1H2AmbQL
DZAk6gAPdVUjLEjax5NgI+1U5o1GLAU4saGZ2XzXMmhaFSfuIVf/fU8LzvjrJfLmNRJRNwzeu0/Y
e1HBcxW+yPBKp1ezjCXDmAIq9bS2NE/77neU/nKhEApi1v8x3/zgP5NCf/iv5C4iWWBOPt0pUG2E
nRK40pJMp7LK/bFBvK8r0JEQekRBTkFKj8DOCWHnCJoPMnGNWd/aOQEcwwRdS2/blRrv1t1ViWAd
YBmAXQg/kfNAcoJcOpcszFPjFG1rkIsn7iW96/ueZvnpHZcMMDbMjoontVOyvXHp+9yHDdOLiMOO
xTjY++TYvIqprCukHq8EKdT87v9pxvML6SQzJ5wKa/Y0GDcFubHgdtmEznmslddVqIDUXpOh3a+9
3d3Y66zcJTwDS6usuTjjWgnIDSqcWoXHlSRkIBd0XoUsZpdOJ39GX/L8D2V6ccWgLKrJ2d9AkiVW
Neud1Q/SYfIghxivTfV+APr4UA5Ah3KyP79Kqa0ts01i65/wlFmiDug1c733691aYPw5YU8WNOXI
OZWy3jbbBztjSKUCXm9d9d2X5GEndlY1xKpKMsJ69szDOP/E+v4vPQMxssjBo3N1NkHRUDbQfe/P
k8ueIsbYly19PS0WB3Mu6AW3nXG9rxiO3HOpa+x4rMa6q3Px4pSAE3qA7TUs5+92qDeLb0MfEbTC
nGct8J6R+g5ZqHY8KiKkOK/qJC5xxVYWGPA9ZWyTsocs5bbE6OXu6Ia/yNCn23rFMzMz2aOs4dhx
oPZlASDJl7JOpqnX7U+mLYCSRna8IhgkOzbtoNlEdSsEgSluqDemeyBgfizHNxgaqdvSm3WWtqfu
pWqGx/5d6nCjaVUNaYkgvqUf4CjHMLVrUJvhFEVpyWZrJcUfdIkwrPto94y5Oroi259wBOHN5veN
DPy1+7jV43hSeihRAwBITp6bdDAiKQGAk2fJVN7UZubLmKrjm+CBrPGDKlWOSZMSTj2O6F9sXc4C
XQFbcopjW78DrT+xUP59HOxBJghnmd8ukfkrkTvgvjv9MN/pgD3lAyiZq/46vCxnQ67gEBgsoZuw
nElPxQDKDvfrSWJrUHnPOwFG0cngRF9PxnElo7JG1NbR+bYfSKF/gXsf9mk5aICeuX5JgkVLD5tB
2cq4JQhv7JDuXbLE4pryhsIjP5OglMk8e28TOJTRJ454GPlQqVM5Zd9uw/bC4cZc7INyCngzuf8G
Zmt3weDtZpAqMHuMGQ91Yrsy9obF+zU7c1j+TKWqZT4AkKeTtS1Q/YBvrjRO5GYVyPvWmiZEzI4o
NgwpbgwM3EZcSbkR2K7gzzg2v9S4w80YGihJHOqip5E/7HxH8mJJqxIMJDJ/IE/bnRthz38tLokk
MaN9uiULrAQ8DWHek0xh2ZRT6De54twHR5TVtVc8dW6BuGAs35f4ghDhdjnT7q2Kr6+Ya6fFYy7K
T2BZnYHWBKKYBJjZehURu0EyzoF73dkcRfFUA5MrUaYEETr/MssfH7AYfKTpV8EqwyiMvNNP/kk+
pP9ngYTtdjDVAfgn10LCQ4rkgk4uptgdmhymtt/hLzh1RIwD2IB36WbBx0SPRNzUTyld1u/GpavP
HjxDMI9xNCXrehCbC1nZqhvi4+LIiCpcDhZljDcuOfAolRLrVv7tjsYtxBvqpYIzWhTd+hRNj5+v
3XZURPzvWJnMq22/FPJMv9DG2FrbfNb6xg1bsfK+9W9WpSKpVEkdxw+7EBCo7NPluZm+pO0eHW/3
rJ3qjEa2G57DNBZLJ8BxlrnoHPgRflz/rMQsD2KKWUCallue/IXECxVLFeDQ0Vpnz/y/CLKEM6Jy
4Ahv2j2gb0La18M0BE7KnI23lhmnl47QljBZ31JNA5YlcuzKMPYwwcyJSqT4lDHB0vxw3M82OhpR
ocCRUTGiJSTS62RnAVDXEQ2faSvkSRTFUGfNZfLdlnMvsvsfYYolgEXHf8pK+alaYH8nL+jZuNi8
gNPSIHX1iuDm4KWrZh9QTI/P2DhCMs5HUNaLBeL7hJRp1cEVHgYcqFtI1aYhyZ7QF5zKFDf0xGGR
eoT/xd8CzZNHc/GeDgs5qyP5XasgDy/Idg8c0CUy310n+4+nb9xaCBIb3PEhtTDED2QzImc5jf8x
rn6cDAk+cvqaDdasA+XL+HmBGpvmqYZBQoKbMHRzOg4emWZJcyicqQYMKpyyI/jf2sT3yaXizC23
JaW7k9IwecVe1RQwFqlhsi7fvtSB1a/oaqCh+nRG+pWGisdCDygYteLM08AfrkEa3XiU7j6O8ntc
Kd/DhuM62qVmmGqsKDgIOOvXlIBlAJW3QFV0Xi7V2n5bQvuuXuZkobmPSzacLPyEiKWGCHAeLlQ4
4b3UBJS7+HJCHawt5IKA4klPo8eaSAXhPXqEbDV+bgzRqAHxfkepQkpSsfC4p194YI2wrsxJkZQG
un7DT0B0tHO3pROIQXHyrPMPwNQJjU+tnjmggBDbu2chFt+W3o+zygKmMaqXNA+DgWqBAVhZpqOW
sbr2Xskl+V6fXPc2/kkiz3w8BSTE846FrSVN8jdqizLqADHxmJLFJ/4umwFtma3pzqaQeZbzravx
QKDRNYi9HsStEuR9ByZh96I3hMmYq4sCLTuhFyjrQeyXLvI/4cMxTwZ90JuMJk6nkKPYsEAPB2zd
+NnIF9UBlFyiRflzLzIK2Yph4WK40wW1CyyJXAGnwGAapFr0uV/96f1bgkiuEaipjZZo0KaXqJFZ
UMNCH00y8x2tB97CVPTWkB6LrKC6BPut0s4EBkZLGKeQ7J+PqanHhRMoOXz7JVtiGbyGUUtCTIhh
+q8m/I1Qh0VvMurEf6xv1SD1kjwTP3hP18ClXRyrUUdldXGCKXQpcqlWwSwQSgss+rO7A1egozSm
IgzwLtzoOfOkabyibR7b65TmZU3tWuQnqowFFV418lbvlIJSKNvDGRG1MUfhxiJxc4GXtrbTfgJM
a2rgqMJFUfF5UrI1bXf7bu/MGEPKSopwOWqHf4X9Yi1279FbFhscj7TJHcwpGbESzGfbpr/yPhwJ
CHEs+0oNDes4xaOkXokXmSOTM2Tj/lPvv4YJFDWFtYG2pjQ5BD6T1gBTi8ZON3wJezPtMO/NnIgI
RvDvvY5Kg+TPWqU0iFj44ayM38Gzo5rC/54nhlh1HUOdfMJbXw6je+S1uDVR4FIDCGwg1GB/E4kF
RNlyWWd75YJAcKr8xyHq12+9rZcuhBp/pYYcSM+ztt84bn8sKrOYxpGXSSv4kzYACy+EcZJYB1xM
E1ArlqMAV9VZbV6iizvgf+Fg6ecDSH51nyDCeh6ySKrrnRQVbLNsDU37+vVUR9VSNUW0Z5GEvtwm
myIGjUxTy4Ex7CB0Xh3tI0h61+au1VkfUR63L/uQhoqnfYxM7EVndiKfOLwaVfP+5BDHV0MSUjNW
fcKcoTYeKVyqTCCMgX9ItaoAlujxbXab23tHL5TWVChHpOf2kFqMZUjr8jKW0nIkyUpAOc+CTw5o
c4iVnyLJyYTAqeExOEx+qBJp1woOhsVlSyNLzVL2j6T4FKsPGTgxzu1uvsO5ImPSLmJXkZWLI3mk
A1d+lplQSviSuYMaZHvBHYYzzHra+35rQh0gAFscMcBrn6N4y5hSuhy+QHxcL52y5tvg83kPu/tR
FNByx77gQVbGFi3d89Vz+29LQfGgPWJ8Y+SPW6LTwW0wr71zQtYN9iZPFLhjqF0QfbsLSX0ej5+w
wENg2ib3+v518YU3Aj/ARa43pffod3P2A7S1DBvmFQxUzGbnwTySyjzEL5YrJ49tyFCR7pGwTQjN
ly65DckTUiOLjJN3F5aOIQmPq/bWVT2QiWT6e3N3POCkAgD7HfcW4Rq2WkJC+hmQ5sby6jGAuYcU
FsZoL6KoAOFxUK8QWObzKhZsWn+qf2T3CyFNj0mPn42XnUjcnTZbm5c1xHqLtn8/UN1KmP7f5xZG
h0i3d5FgQA8uFYka5bjafrOMXmIQRNlu/xD84k7bMWvvKbzWCyrj4IW2rWyqPg1Wf4+Q9BJ9GrmY
Etc0NhvB8d4LBazNdf+3L74ENd4lcOFE32DCQ2mFYvVIQ3tVjpFuszJlHMRU/VvRZvuy6SxtV+x8
wl1qJzHkQd5R3epsbQXihoH24tMQM4f2IGcB08nQ1ePTmDOzRemZWdQigf2Iczhyibg7HnrIXzsJ
YxIvCKRb++oW6j7f6N2SPiCsIUQm4PcDuqEgdnrAHFjTYbQFRven8H4XKq5SBJAY8X05K3Cajuce
yn6Ds3McWZB7XjqZRymt9oSkHPrjEWWIPMCEO3QMoAwIyDJ1wJbF0qFmpldGuQDukpx8cxNMxLPX
cvNUo/C4aWsq66bQ4BO+Sv9kiMNlFCKBNQEYBKAhwlzvOlv54GmlIitlCE0EWiPxww9Twfy6G1wA
CS86Urr7l/Wq9XcDlLBbNGq6c1L/fIfWpTR3MpWF3V2m6HdDFmj40y9pIFHWb6EtIJx/LVXAPEDL
Wqqm+Uy5BikKuEaNpcJ/3wNnJpTxeTVn8tpZBzxuxXw3u4VbcudHq79wBhbsZziRQPP0tzmZh2PY
4vKO2HjSNDwulPHDYhD7OWufcsL6rW4sA6GUXyZI+wHKg+6xbFbXFq/DhHcgddJXKF2LWY09C1q1
kxMBugf+8WP/P9wcgas2+gQBzAHdEhtwCVLGavrtTB2lUKzgjq+jTyKoFP0vTRLptqmzPXi1lFro
szz4UEieSq7Z1EJCsScsTgtML7XDkYniwZAtHuefrVLwkRNua+r34dcd2WveX4ROSm1lKJeG6tTM
zwtWIkNAkGi7K66scdBcXJuQkkYgJQxh6j/CQvsEtiR6kDjdqq8TdB8gbi5HEST93BWz7hySFZKA
mPznS2rqRqEcw2qHiH3AN49vun5PYycdYsk233HEaz/cGSrUIWHADCs6Wipri5QEZUyhhs9qjCBn
GIEvwHnEatWg0iZjkTxJmD9sOIPiqLo9Sy8OFEp76Pqv+FncQY6Bs8u5by8F2ldXRXmwOj+9J6Fo
GZ53K0+TpVIOHWAvp599HzV/1C3Jv4+UyHNVvRoWI6R6J/Sn3BYTnUOi00HA5N6MVQ2k/xKyqp47
fmeAkO46ZqdXIzjkYghvT7Cuubm0687de7siC2JFp52LkWGCRMkC0fIoQ0C4/v6gQ8r4K2aQut0I
awV7hvE9noM8bHBm2Ns0bDE9TI8UCqT8Mq9ZlUc+E42h1ojkT6H6M3J0ZBpwWL3SwHqVyvPeb5gM
qrwTjl4cKVSOkiEDiOnlVTwfQ8PcYUf5s8JdmEqWXfz0m1f0W9BIOhQCceomiXpXL+QcZ8Ug9KBE
waDUUKEatJIGnvKh6llPzlerVNem/2qezEUfgfMEm9Bx+eScFby+0984upM7clXgQ7LQBUZDfrpM
uGr3rqLrksjR18Xf4Oz/ahOt8ot2VSU77v2EtkeMLKTxUkfjA/PnUb/UkvK0Jk+UiIHixQeLh5FL
O9KEs9z48o/GJwRSRrPGjtcjHW14EG0F5lMZMzhrqQajX72Dcta37M7stFg7O+oCGKH7lHSz0M3J
SuojzKCjSWNfLUGxzMdX6zCsf+k1xcSSZNr7DI9DKT65jxirurEUeA0nfmC6sjJRak91mSKdDC9d
g7/U5oVWL+a1QghHjMypVG85pnS/7+Jb1CVvsvjoMmaAjtHYmBpY7Odt7rBJF2tsPbxSclRK4/q8
Riz4cjoDQoSrl9VPMYhLEGtSPMCWDBhryvvOOHmgbC1xVjuiyKcxLM58sv7gzqfMruHQ/+ju2wJ8
aOIKb2QGZfJZhFh1G5dzXUYFpPWTcLClt0LL5xirLJ0xs+gZehJsEYAJE3+6+eE3JUdgtoPe+kEC
M49308YAOG2RM7Aa/HYk1R/xKtmzYXotDz9ocDJahzmIaJjF4qXVnyuD50zxgXDNxVAW/sldzheT
ylVGSmi9iI7NNJBa3P0yDT7Q1Ee6URY+55olMJdRwhxwinYqJTm5JVhJO6ANJOHXYtDQ9fB8ahDT
6lHjeWLCv8MPh+PJq30vEf0eJbf7ntUoEsY7e1vacIWwFNOCqztGM9cZVpsKNpVw2noD8cl2cnV5
2HRH6r17H7sprgwtkyGvve/TljoGxekHC6Nr+nPW+etTwOFvWV6JpTRK4W2hVQLqgZZRNlHGuuRc
ZM7HS1f5SbhoRTw2EmLJQ5J63phSdRejUKIjUtGlCRRm+U0ERHL5gAfzCmL8p8xjynfaPZYsoMum
zws3+mTCcOq+tTozBIiz0QpwbZKBJ8yp5G4Ri3/ZiL3oeRaX92AZGLzaTYZGkrRmwpgmWjG+ZWgN
FS199DlyX272fXI4HaPOXkSBea5uBRK8nQUQtRrYmslEYSkqy+pNdTGvHS12g/wXzAdbUY/8T9m6
XActMtpx6yEOAt+y/HwhPi+jmL6lAXhnIlpXhx/WcQn75vBXozveqzOjY+kgEr5ITECrMllpYSIJ
5S1YLKceoMFcir9Nb8nPh81QKL3dblsGaYLYG6YIGq+7DFHAWfVgYL48ADdnWGn62HeoDeUVyopd
igWei9eMHobGihy3+MbKFiVjNZo+Fp0kqwRGQBqtuGQBi3+kQ9e1x6Rp7A9vhyO5uvFjruNAN5iP
aR8bcDl6v3FFdd71l0ZCwrPaNmjoq21Gn0a5dbkwIYfelvpz4JbUMaiGy3IYIO2aRkRl5Nou6vre
Ltr9K+KiAl35M6fKgYY6xmavUTDYs/59olWK3556ElXymUkvC+396VJ36SKlxmPcxnFP+KWA7F/6
PyylLkXyRlwpEWr69+gm6JHw1OiETgv53Cop15iGSf/jKZwhzQlUTud234l/nQauZVC3w9N7by3F
r6Kfi98MisgVxMKwblyssFrHE6BCm/k3MhQZvo6vd7o9LWYkX18Gyi/ALiXz08piKmiVQRLZBcFY
Ac4DpkUOKcbfKxtUm4uy42ksbM2P2vjCaf0mWfDpTm1i2TlVMacv6JUefVRWN8mbdEd2I2fEERYY
ybPU/yoEiu9SkVSp/EI0QrOFrNCLbB2kGc1vUEDwrFFbvlsDk9WHK1BhtXqP/WnB7EqA43kVua2q
RHLWp2yst92SS6NPojl7UfejTCm3s8pKkxAAzRDh8kjlkYxv5MscPrUR8criwZp5KlzK7aS1k7bx
AJgPjXKwhuKPXrp5+9Zg2iZq3znhyez4wVecPnKGbalN+Smra/5FkrVceQIwJsGCLPGnQmszFDUW
bGdaKvJfgP7QGYlKgmn5a9k8+1E8bmaeNYEKUoquBR2l3V0AeH++BibCPeloJU5zksz33ER+ESxW
0DumjSfgBWlQrLw5ZB53ZegiIswB2krOU0G/nKYG9bhVRkOa/aPjgw4P3v+GLRCv7c1pz5soYmrX
DrIYLCw656RCU1B3gosWzzdqUVGi5oJbZSP18FK68QI2cfoCFzMDEnQgJM6BtAefyEEJ56PkHxUP
HcF+ezFrJUUWSmt3rUCCx7JIICMrx6cNBJURGEU/KXqTGPwfS34BmIqTxolmtrFrM3rTQnwqs40f
X39b0RrOk89KpJUZ8kgMqUW6ePyIviUzIGQPsgfdYSfYFigxFBezYuAa8Vy5NTqE70ZKGVyVxWSq
L6dGJya4IX5vIEIrQbwO9nnS1eSvCRGyZPs+nEpQTr/H4GjIa0Y8gTa05uKNvsjuiM1kyg5GPYgq
Voyf/EiC9IMzDTKKlr1sSyADQHIRB9BUp7YGyqRv4PFgW/xMKNyv3E7VcQkK7QU4/mJv8s1NhQx4
dz0kUgJfVAZRTXChsX2NrtdNtqvD0vLqclsUWCvFrpAGIzlV9YEM1RTiGHcUriO4XpNO+13YQuFl
0e2EJWdMMsaiA/oCasp586S19vpmprOWSXWndB5c6MQJWkX/plm2S3IqJuoXxJaNu9Mf0g1Z36gE
lQhnqqKY24d688XAFgYKazjcGEbzwHsdqePcvM4J1tN+q+teEmq+zcqY9wta7Nlq1fhyWnJDyby2
THww/G/4O3q0wvUxpNpZTRyXBD1GiIwAk2qT2rnf1shiy4ekwPc8ZM81SSmS/eEA+Yuu/lvYq8cX
ps4wFQGEw2bJPezNU+r6AyyfpOfK6IhYRCPSP4bz8ovq7f8SUVxEn80FPHWYw85BQINvb7WmJcvz
qbuqgQxeT78n++v3kE8tb/edqtxOd8Z/Piab/9gNVMHd+nRYGG/WjYGcqqssnCEwaA4lvr5hW4Lh
idYyiYtVSwkokxjt9KO2sDb5lnmk8siiEkL8nNn8H2DjRD8PFPWZS9gvgd09ew3xOO9yUH2MJuSn
JzWaQaVmTgUfY3sHhhB2QRxbKUpQTz8l40PkPefkEwGvI5iMz0j7AVr/iUsdWk6TLc5ZzOPrB+oL
bujwAaBoZvzrwoK6OsFj/oMId/GXGwXkbZfnAa+lFdrUhsZGiFLPaiP1ZGLcnVKA93UHTrSFqU2W
dAzHOFRwovgCJvDJS7EGPQV3xE0KfNuiMijgAPlzSkoK9fqWoAcYvqSgCMxTjBeJtOEbyJDsRJhZ
rppPvxJqMejQdYSRJONDhuXOvYB6q7rjCVu3GgjjwHXa2ej7yPgv/qHFg/fHJPq7yhwbym7ObfY6
5iLe8vM5vzPNrh0bBlil51FjJUOn3SUrOiV+/BSoTGLCpGxM4+TFXG2fZ3FpUVQd9cXLIApStfEZ
NbcZSW28nTGOt4WPGaMFO9mQPeYMhqUTw3NDdZEDcfEheBn+Zw7ezEXU+CjiRpQTCAGE/NvKD73m
KgzaXX9Ho8NLw1i2EGjDnFUZxJYGjVI4vvoG1/LyfCTSADbLnAlvU2Is7y4vMU/L/s+4sMPlxuYS
c4Ai/fdNj9UENl3UxIbSWiSiL9tjIaJB+KpZ5L3iH2SyFii3H1MbMNlJLjD6fXLLq34TZhVwCU9E
WumBz9DtQbUrQ6xp1Qcd7WB+kdsuWdy//yp/gWMPMNTxT1ErE5msnN3PlxuwGaIpQ5m1DKG62zXB
NEVYhDXcYrnd1a4jeK15hbILOS5Edk8EzIfwHVzUu4COPLnWF+57l8oRotnpW9XiqsBI3pddKN+O
BwIrBDDqV5xoOE+cK1RpJvTUTBK7AzTOuNhzKUMuZayfKpZPe88RTrRWH/bA8hmQl0WiuZ/SNBHG
ThyaZzpigZOOILStncc590u48QFDPh14GivoMcKSWG0bPm7zcTtun6o72MzNp6pGIYA1g4eqpKcH
4muYr1HbD6KH20fZQZknJwFMCKbEKBMDieFs8/9pqks8pLrWk9C3XptSmu1ePTmGZnjXs5Rz0jNW
MIuI4EyWdiEoNQIup7L2PEsaetqPOfhN6eJoLeurCz7U7ftckCMYiuSdbVOA0HOWOPJlhTxESON+
JQwT/nOu17HsHF0gI53FzfbqZdMV5iGkz/IDQLk6IZY9rngVu94QIyx1PjlFNUxP4Qq8dx1h0Neh
mtj/Zcn/uXlzidLNgEaX9kCpIfS+jUo7yyxP9+qiE07huDTv0xt+ZLfva6iMyL5U40JFLnslMeA8
e98qcyOlboQaDKMC9whEwJY4RXsblYPU/qjGaNPUdYNOl/9Vkwws2OL66/fv85h0pYeMGJHmojAw
0SLEFvwTCKnr2lvkCA0nt+qgnFxVYSgVZinzG3m5ZL3KR21N0ksmz0fOYNZ4agUCSmoo+zPtVfT5
5o2LINfxEbixOT3SA2MYxs+Ugi32ed6g4TJMayGgAtnH5f3kNHHP1kD3y7rNxY5bBg1i4zfcplVo
wtdhUVdzacrSLx8pCyCrLIdzbTHWLSvVaO/ib75CBEm1+Bf47ar9acKqa8f5OsTGKU4rmLNtNEM+
r/exuigEjYOcSW8XQuX0J8Q8Sr5hfdZBsgnKUx/Lx3lDA2LWGPOXAWwqhB+YMSYWVF8bYoN9itwH
42Gof4FI1DnHGjGhDQ3DiMsaox1/ZBGYJHqDUH6tzaBbyGC+ZAHoWwP068Y4+c6BQNL7wmKgSRDi
bwn23BQmY3edYLKkF2u7ya/7SkHRbBlpJyW+ewRodLDOnweJux+8V5WbRUdMFRvsMnazCdZPUU6+
Mikwk24I2M9EDCYIW3izP1T/wUKGoAVFS7YPTFfb9ETPAuTFcrhElD+rJKjzt9pA8yNDzu9PwK+a
nt1lQ8EnGzEo74ZrS+UkRGivfpUYLEze72zjHgVwmXv5PBHL4RmpZdotB6mpm2tImB/hh02KzS/7
WArHSBo41wt2dBLVxV+zlgCN67oRHGdEiSxa5ZFgRz+vE9mJcQlQSoylycrZQP39VCJu3t/BgZu/
wCEje5bTwd/YeaDqHn6JyxFbj8UEgARfYOg5vk2TRkAgOp6Hvq7hTIyDKIJ+cPRN+YtA6CbLoEBX
gNSIMV6tnW9yNZK7zbizaBFWArWiILp/njbYBcLV3ggOmyibxKU5kVXFD2drCiD6SFiizWDqkauc
owpRCq2jrwwWwixYxybmRJ5YnV+EF08KqhL4/Glkk59YWY04I7353QkAiTP+s7VlgICFe1u4fnPz
UbJQ89GHmD5FyNcoZiCBL5nJXSGf8B7QJFO8tSI1iEPTSWPswn6k3m+0W1vzisCcPZEybVJqaFzu
qbkEvPpONdE65OaHraMluoiTmKsELs71mJvDYaCHojWei+hOnp64wKbfkCH0n70D5ZMfc7TDj3J4
7N27hS+Vy61BWFJVpbIcK6FzWf/fE/uhFyUuM6jNmC64RJFseI9murSuBXigPH6UxawlQaBDJI2i
g9zoPZHQdH5BL9Ag/SUotfvhM0q8vuYJgeoGN2yDwKlV3ElaskvWFrVDJ2NR5opUIO1i9gUmdM2U
F9GJSWiD23eLVzT2COEzquO7lt/QVKpGPC4O7YMcl9RbRQPkOHa+eV5JAf7SBdDlZSl7jlWZh73i
s5eg0bvUXiLroWCaFiGaKn5FFbCbEE1JWoex5VqVXa8ArokmaflZLD+WEMP0w1Oks3/5QQjEiwsy
6ttnZ7I/OY9w3ekKsvBMYi8bHrE+YEgTHhEXhTLVuREo3Csrphcs5+Y/Vtq4AmyPJB3NBrHZQN65
frZZpw5e9F1wCKbzOQASTs6YzqnTezWNibSGhORfm7UUNs212M5AySUczDavxDLhVUZ45w6uNH9o
g6ogDqmptqgTLj7Nsjf6BgM4Wf82Cpb74IeQixl2ez6XZLBauUDpZ7wXQVgkAN+VjilA/s4etmq3
Grlm08PoZeNHr017uyXP9LMoP9QENmFa84BZyUATJsD2zbNh4l9D3M6OHkX4CvNNNB7Rdfpn2pOl
X2QFw6W9510OkiOzxDxQCab/9MdOl2HzM1YVL80JUwY1ufpVrRRihUT3/RdYSELfvw4ItKyckIfD
43tIIBiDIAtQaBSY5tn9l5mheueJZ3lSGMo1Kc6B44rGCaD2zGomYPaoIN3KsLs2bMML5mJMGQit
dQjAA8qy2MjEu2CY4n9qzWwYGceiezRUl9vZYSZQQalxrbU99ibralPwROQVk+nargA7Mnebc3++
mCyRoWtQaDgkyDjwnNNwPqruiKeMh9GkiKSzyl6pQ6Kfx8YnRqhUL4ld6vlPZZQ2iYJnnxomHAJb
sQsnx4kalDy4DvXlkv7+C4Jb+8NLyVpl9GX90Jp13AuqmeoehNjL/Hho17JNAxmzT5BSV10vRHot
BPe4NYK8ywwE5W8/TqAcdILFsnuiqn9PQqbiK92SQYtbI9TXJyS4QB8PJZBy82nWCDPOgtl8slXo
BGwZ7/ku6smffu7BEc8tWuLLuG1fyG217zNFFTa62yTJ7CoYxr8Xmc6EYhh+qp5JCQtYBm3jGb16
T2EkQxqJuz5U6ORJI+bf1UgavSzzK+l/IProoy6KkjoPVNOTSUL8T1Whpk3Xje8EMQjvPQJAOJxJ
x+etxfVySrgBcevFKIBozGB4EcclowSphKlZfGUuCXeCTGqDBk4otmpPo6NGO0n9gv/uDOevVVXi
b4t57zqoo0WIFjDkUAUJ2WQzynuXC5SRKXowgoi1Idx1KWDASTvcrTs8HcQpoNMFZmqqlLFgZkDD
2zFchVhVedJEB0gi1JPAh2jB8J+Ip3OnOkwpcVVSJrQiCad1PGT2ExBZTBLsmIi0foAMvC9EiB6o
ZCIFnV6mbeBj0U5eG6n75WDCSYHxIyqnP7FcX0A3hiP90aQaueZdYqmvCDTNjHTy9IaU3oPCUb0N
4DS+JJ/4WM8z+KXkoP0VEaqOjQBeyNgFhoPE/N1F4c7ahQgXG5dKXahBE7fJ7aLDm8eAE/NB30iX
HC41O2qz+kJZk5lx22ZuJLbNVSJNEZ3ips0qPj87QpGVOGxQOzxWlHy53fY8p6decV+E8lXk+7OX
oTad7PBGRj3r50Jmnl8LEUh86VelMepo69w9C5h2v+n0f5skWv19fZ/vYfQCEhIkPGn2EaCQ2sj5
qSE3TZrW9HxJModyltbudsxTeQztzBPvRY2uhwXWYIuRrcXOfjZL9xLVCcYxv8/u+PFwB67KJSI0
k7WmKg88G17M/XrHlndUWlG9VclxjnqRKL590BFUKF9zgrDONgEOFoIdpjArru0kP0ZfC1EM8ATu
HY9tldKfrDVXceXBWLwjLHhz4nFy3IE05Svjq2ZRJIo7EVNhuHLFJ9nDKNaczIhw/FeoyVXb8XM9
911Qc/RtW2brx9QHp5WZKhAuMfcebp89gryEXjIEgTPif32PCUVs0QbaxpmPHmK4wSKoDv++TP1I
JaKmEX7rIU7k5096xQnxTTNq1yju2KLsxjzlj80qiXeI4p0XBm3UuQR/xn0DwyL0zk9MCIpv2Wy9
UbyZw/VFF9vsielHBIdZ7BjnWU7jy4eNBnzTYxyXVMqO4zJoxdCzHYlzSYlew3Mz0kb8kri1+Gp6
nJ/gg2Ysw1Tcc11e3NMWrsN4Pogs9c/tikiyPwRBof8k9gM/dNqW3F6XyArFdhgMuOS9YU/uaeft
ipVyUVuI78hQh1YXO/AyuknWfrwzgpDTpvX3UZLnuJW3VXRDs5T9O05+06UhMxcHAKdymelGecZ1
EnIkFpXls8F5hkNMtJVHzXwucLmdKhRBKYlc4Iw/Dv7SKTmd/dA6/6CSGUL27n70fui7LqdPJILb
avJ4KW3v95ypVsVng9fn9fgl2saDYVxDOnjbcgIuzh23de15UztEoM2OiOuYcHwhW3tX/8YVjKiY
2eWeNPSmM056Rf9mayCBcrxiSsaIRqPSjmRyLxwDAHlCNUmlLkiJCG9si2R70pYnLuYERlKHJg5Y
MNkSEVuEYaMaMThfGMuwfwJEuYnnaKmNVcx5TPDNa1Q6M1OQDHCEvPT+I5jkEUK2LwvxypSIxsk6
Mp+ISiFYu+FgGRYTAbdYsX77E6lQft0ftUE4xvanWWBAEdApjWbtbQicG3gmKU+UvXVodAZm1Slk
LO6ZERSWJcOPP/WpmuL0jabC21qCFYNXK5dBRc9PC//QlmyL1fiQ5d3VlNaFyBJr11Ur7MO0In0J
uyTV6iVxoh3R7mkbEQHqtTUk2wxON4Oqf3E7qkeOCDXBJcs5QqjPkDac1jYXTUlCS6EqaBOMAXot
4/78PWvqlrf2WIf67bvEjMDYi4YSqDaiBeUw2XPZ82xAMISX0d3IZF6j0RgiSzuW6SU8mXRLySdh
f4Dd0gtT+F2Ain5IX0DvtpC+JKhWOwVJw1MDszZidpvgm7jPdb6ic1A+bcwYGsuDIEOL2daQuxPe
a93M4VbbyGSPbo7roUlkpOFmQ2I2ctxBp9kFdCw7bza2LilS8zPLAsEQT3pAQEAE6pIsltNDDvc0
a1/Cpkji5NGa/HtpGUwZdb1YRKEXewLBwIvWUqrGj5jEak9+VGwVDJ4n/E61pXkVRB4N/0Sn4ktt
EtEFJZkYr1fyXGkgq+R+cV3hg8sb9vQK6D97gLj13nPbKSq6MzNgH5ektGP67wJasOsnXif37w5q
RbP2/ePa7Dn3gFdIFYjCDL+mYgkTKaFRLKAhsiKNfnTNuY+gWxD+b4lkk70Z2c1XOzpkjwIQZsCP
dCRpt6qqkHfv0z6KLgL51w+4iLUrJ30C+4mooW/bSWrQgtf3hUYXlhAvYWYowSU3m7NPuENyQCm9
wNSeCOqJUdM581IJ1PthqlgRteyfX6xE9N9x2G30vdWrheDAzIKj80rqAhNFJe/udr5m7Zf3mnVD
PsOhkS8geCFtuhf/87e5fDqeojjDhFlsRhV/F63uq036JAvU++Qp7wvLkG+57IFBzJOxm0BrEoPt
h/BHpFzjzA0TX4/eIA9l4juDIabazKd+hta26Kp7AJt6tvsMGHH5xIlUFP+dR+IZr6U87LhSoDhI
6hoFEYwnmOy4ARI18oe7VyUYOKr/VcMDOIDXQjpv0t5AlrLvlsQYERdK+5ifXWVo5L++6gl/NbzH
Z3QvwsjCdi3t8nQzsdYBu3NPGLJF9Yncafkn0UGTOwzR5Dxb82IifTEHLrjn8CLMyEC7P4VyIvQ8
4vpqGhhAlc+uwEOwlvSVap2bG0MGKADi2MmKCH/n6Nw1bdIsFnrHZZGFcIaVaEuBJ8VQNtO0UV7B
3Ug02T9iJbMrxSFtUEAc/BiDBq/BrR5XJcBJAQ3iVfZV3+Xtu6rU6kHFN+/jZx7yUMRDaf8KYWRV
PBsUXJ3kDcVHu+LvYeJlnt/8H+fB8OUdR4Kz4kbwbY8rO5XzHHl/vtZkTfBA0d4K0P6vMjOnhfs9
nEGSecdifyqbokcc/3PYWX2lU/PuMOYCQNj8JYiq9RwB8yyMC4iWfAYkaH4jsZxu71za6vBicrAe
RcshiPbXVpX1G4HX/z9YVwHtOVy8aun+XlygoEsmHGBehQRnC9/Kb2sBjTT+pPWTttCCU5iv0XF2
xTROZuGEpEgPumaImYAAx1sUUfpSGCTGBtiqCLKfEV7SKUosN6POEs45NhfMdNT53/J7ktbaFDFQ
k5RQkeek5cSDJSgdJUBegXxEPj/ZvTppzx2vJJvBmr1D26Oj9oWJ9vt7+ge2OLCBaKMOVDxFPQMV
/CFAK3zq7sth1e8ac1AmdxvOAmeRq1Aou9tEfA3FOid0x+T55dTv9iDhc0XeGSOAgAbmVCDW+yOo
APBsoHQjvWlOFWzdQL3O8aGJ+zoyTtn3+JYSuwn5HTLm5bBobim9R+e71RcZc78xzqYSbDHwlt2L
AKOXYBAfSvLYob6b5qVVb5bU5v/CcL5NxFnU4whhQf198eGt86v+PudwsaC9deHFjMCm3YhAzfwo
DHvKh628WHLOlD4IPY/bU8DGruy4PvWh7atsthMEMW8SOTrrCJUDDGh83eSFJLXtYKcsW5qfLcwm
jKlOQATmvcT8yBEwJ+feGI+BbIm+qs+SG5WdN4jDVwbW90uoKhe3wjb6ychDx7S8pIJxVElQVodp
VEk9iye+IzAcTJBUGWVGic8+G6g1KMUHt/P3zpgtib36lO9R18V5onFV7Ly1rN1lWk4Xq/ObhV0t
YGs+0KDyDu+3gasPQvKTDpbpkOyRL5s3752D5aeur3LranvsobC3oFeJigHWsc6MIKtYJu402o5B
4wX+j4yPB2FY/lWVPY1eHxB6oRZVLiLFLsOdXHXh+RiU6ZK+S2DTUPcOK5yIRveu7WfdxBDh8Wfa
qe+GAUn5Fbr1ay/xnnQVTNhttEJfvaPJBBHA4fJceARUCIg08hlGA9CK/xN940GpcONHvkkA3Zjd
uhL+b4Eca+FfIGJi4DiCp/SCJnCbr3tshkHTSZ9BAGOxAaZb6njnh9igppl3UrxIAmV2RkWCgk9N
zd624RSOFWXFogUICrOAMMWy0itc0jT8D3UKXjIkB4Y7NkIxH5dW21ZbJRMbf0yCwdVTZu4aWx5x
5mRV0ZMHUHsy1KsuXwAqLPA1FiOYa8rZOL/oAPLZarXKxhJXMya77RaDWdcBw3YZ3XxdiMA7AH3M
+/uTzJ0mNs4K9QraBnoFTNXybtD3lJbdYHmcZnHP1dIihNXEcWdQCL7lfn2ZA62tJnq6setQ5hCm
7BJ3qeH62j2E51fRex+yoqSNohX+k25L+oV7u2sA2qgFsCglDy/6cLQL5DL2hBztG7O2YXFsb520
yUjqy2dFL4mNK2adZgPdIGYYk0b+EyiXfBvchsW2+FD3qgVBY+7Sgy/KYLEJMI/lLOzqaIPJkqyO
lN4mwPVxgtQEbKnq/a6YnWIqsSstn5HkaBr7vq0wPEobiXv1MrI2VKfbBZWXiY39rPJFp4YFcNBh
VLCsPrUXxm6WjXLP9uGR8aFJVOAwkGmibvvFobP1p/L5APyVPoSPZycO0Q2LOrlAJ7UrGWYGzSFb
Gkz1XPdMFH2Tv8RTLw8W3y2wB2w6TKrpwDMeVty10QEafPMNEfZU1D1FQgutNwl2D7PrTFNBhbxV
ZmWHsrc4KVz0pv4DsbUcML5ubOp+d9NbRWU98WCZE+JbTSQhmBKqHhxnu0JlW2UNNZgQKfiX8jkF
sG2JYvxmJhVUHZyi6k/O13ALCDjJtfbwKJAEM+TdDq8e8Me5F20Wy0ybeWrOEGBXw0vqrvBvSzB9
XW1YI+Gcr8+LbZ4uSeAxdSMTe2ZXxnSFs+SWegXDyC04ImCtWnRViN7DpopcSyA8vo0Mc1baoNeq
YcWQim5yDu5hweV+qSPFAqZH50s1PW9GBzp4D5tjClPJVkiQPrkePrVx4I3GduIVvmRnxUx1Ijqs
WIFtfeJ7vIT7ZoESpbNgowI1AcdcyojmuVmE/6CCot5McqVqm1/1ORUBR3kGSJC5gfPSS+czV1EJ
1/9op6CDlj9h+NcZ/ES1ssau3IuQXGnBNJb1Qk/sP9lt268gkye2T9fYqr5g/JiaEVzGsG8Au/p9
v6xBxv7ydq9fM1E0MzVzFlJa7EbhFnNdFfk5wyfKTVvYEGAztLyL6+F+724q8ETHOWeH1aFyWhSe
vjI1UnCeuKs85GOtFjhgNQpywad9jcQboOXWYAgTZsSmtJ4TuXFbB2q66uDhvhv9S7SVetneU8+l
loRmwM3EEAaxv9xj0mJB2IP/nkHcxeDpTeeRyQmFC6apJdCkTDxwg1KoXdMNwN2a66FAaURD5oia
02FocvVkxRpLDeI66prhkEEmG4uPdvt+fhPXfdr/SfKwsIPT9YDK5jCFxormWOlPeHz4hmphm2h1
QlSENjvmaK8Ehz2F+m7+Yzl+aZqOE+wN2sA6LS7SDYnBVdioO2bW6bhAHG3IKkfRHXruXDTrXiLS
2TDEpVTzmtSXneEW8Xf0SYXiPaVxAd8s20GES4AGCAo6l2zNm1rDQrItAwb8Y2TXG+p9QJSjMbeA
Gy+XNPkiPVoa94obS9JNCxM6pfXMzm5DthmPCqNmXqN6ehlwf5YUPf4ISzh0hs7X/F7v6Mt7Qmls
aySnFPKAj0UT0USwGVLKh+zsKJW2tOLVxirpy5RVfOjFlyD3+H8gX/CTaofgXjVtMhFzX3a6HF8q
o1WJL1DDB2rrqUaknZuF9CyzPviOUsOgD8AWKgx7ZjHZ4NxziRK01yDC3fAYcLEO+HXRCbcFdchw
F+ydY65UA0Ta1rhi+S8ygU6IiCsbRUVQcAS/EDh/v3r0aNoFUAtF4N228KsUkwoYSRMktZSiZGeT
LTlfr8BgwaRTgE1aaU5PiwQKPnNfIh2sMvjx2G86jZYOoDBE0mYJA3BIG6XdXDV2RTA3IC5Fs0vt
Zg2R1TAP5Okep5Crgbji8hg7ZGSdaC+ESyDTnRlv8m5juqkaONnrAa3LWPpQ44224qXB3UIg6Bj6
sXMT+Rg8sBdAJDtO7VvmBWpZWpOw4gqtIvIs/8QMNh7xnfursQOm0gEhTZhaekIV2nJUtSefDPe0
biQUkthC4HKYZuJpRolm+Pi3nJ9xr57ZXTLL2/TxnGQNmp7vzODJFqP4KgKpMCCTBh6njP2nJK53
GBBTQ9aN3eHrjkABPs62j+voUBRMRDdn/vF/n31yDEZ11DraxCffj189f1eVdvp3EGAvEYEIQ9c1
X6WmTcmDHnEpITRX5KAiks2m/cneo24H8MyjYgmXW480FP8ND9oxFFZF5tMv7qUpgEIVTl7Cu7uw
gI+dp5D6EBVLk2XggwQlKzMw3LTdSJwo9eEWvbdXUKV5Sy0+/crVKg9eudOiypIB4APYdp4iEUSI
+VDeHplDeMT36kAKS+Md2SVxyWeaR1tHLocuw/ZDSVXeSQ6g7NYyyaCAKtNK8q21k9Umrw6nRFrZ
BjYv6Szmm0XKK1k77H8JC25VR0qPOvuUutlLN2nSxUhQpPFMRXZK0rwjhCjiLnHryDfF+aDM4oaL
JQGzN7NX1JpmZC9WB5D54afABdwS81KR8vqTAAaOqbL962Of10kX8o8WW7nKpYH+ykKD7fRt7egr
VPG89ZAwc1wPxGx9uxAbr4L9sBtbmBJTTUeFqKRk8blZLsaud82sli4JlUJXN0gEELvVko9+GUGq
x4wkABpdRDM8m0NStQQHP33pvSZ0GYOjVYu9ZYLAOztZ51bQwDkHxbWJpLyD1F+ZyJ660i+6PrbW
3uS/7y1mBw/pezYksd7cJwG9EgeyRdMV9b1mupweb01bcHEhmQ7hWtndtyMPiWfZDGyvMPxy/PQd
gWpSJwwc7rbUsU9O1NyNK5p3VAbjMDIPh3jeXQJMzBm/nCD82Etf28HcV70PJZ162pPXu+Eojd1R
3Il5Ool7fe5fza6gu/Rx2qqEmK8FZ6ip9QcRsuc+STKjFpEefXangfH5kY+YR13iiCKcbWmqoggw
RV/T5HvqVP/pdXXe1ajtKTMs9z5/a04+uDtPUpX+FpKXm4GomnPvyKlhT/UICFocq6D3sOGPw3hw
h2pY3hK+Kbc0uFTV8Gt0Ew9R8L1BjzNoiOeHJLkI91/48rsI8qhg3nVhUHXdE/prOLwRvFa0hqyA
na9CZp2YNS06ov8DpDU9wm/QBu8D2TuLRnB7bfB5G4JWdtsH/MJtYy9BSi1MbiSIuw1oybDMOz+o
YF1auKXiLH/q69ejvJZIbPjSfjlfFng9eaD2xrbWsEQyXylR/hJW8A9Zs+Vqu1KN7tMJNvqLL/Jc
7RY4ETfOOELqRNBZYSvUKqJrq39KHdtVTrgXmLHrIbf65YEngP2Do1qYcyORvhnJEPMDKQWbe8PM
nulLn/gq+ygR4mOLiOghNPC+QcaJ2ixEiBvtKLjvNB5MvTeMNUVjq2qvfP9X/hZfw7BH7LYUYJDa
e7P7vzOclqWZ9Mwa6ZfGzmzoLLtyMHDRv1Qs+C92lLOMH1JbLSPQmYf7bPi3aOIpKRiJoaiVBX+L
+zA4BQlBBSL65TDrScZ4FdsDgRsbBNhbJ9aOT61nGLwhaK/Uuz6mRgQa01cMUfndDopqS8l1VvwJ
PPLG1/ad8Txozsg+I6OUT+5cWErOKWBUurxHHtNLy9b2I1fdTckuvI831TM7TyvAORVrWPXH9D+1
5yRYbLLG/7RKla2OrbPcXO7xhnfIqykM/1/dpBI3fGKAspX3xa1VWLMAxdPXKSTs9F9csArcFqIe
1eiPNrbXMb1W59x0V850zW8WYGFqHHzsAymr7NLlkosOWNBoKz+Ylau34HBreCTRAnuUDbqaclwz
akHo2AarZ7MecW5nD95RZu/+eMm4ZwBdM2Yi3/djGV6Ezs2gZgjYOPRziOTaHqWOqqtFXaXEibbR
UV6NYGZuLhNOdkxtLuTPoursXzQRNFCybDndZm7bnTUHetzTcm3JnBfkK5W4ZLwMRHqCgRlZVRPH
UsNZ8Odq15R2iIiihoR1PpY1MC0nFSgDXTodO3Ln9bmf8IRHlwB8x1KI0XzOhaScFdIk8MrO++78
a6/PQFN6/35RCstSCHjimtQwaPahjgY89+86hLfS+97TYRYWZOn8MhcTSHGpIbZ1wH1KGbOyVuO5
+Bd3xR+YRydGqcAYvfHjGHygX/+JeGaeQ3o7TGc9RBLpLnsXHhOOjVC0tM6VGB/r5qrplVw2W2+U
YAMQ7UqFwLQuTemuXm05rqsNK1E1594T2Z3h6YEcZ1p9MReYYuG/NSBCONEwWWTylblD6yLVQ/mK
3lrcp0f33iOYOCeahmYMQmzxANMzcGc9xwmGDToIhQWbW93q6GgPlOASR6FxFfORZX1efh+4t3Re
WauYb726ZO0PtsCXRPWnxl9ZrXQTIyt227dIUxSAPKmiUalYu0IK0Yki8nm3sM46KiQjwvAAStDL
MzuBMAs02jhNxqduKmlJcT6N5lpe+a6wZQKVPYwVHhDMH1Z0hg2NRKMir4xGLu7CNMhk0xLBRApi
mgQUmIgYzEEXK5h17MoUSAQtVnr5ZtjxQD+s6iryZbvAOucZTGOmytqpKK5/zO/Y9xZIc3yY8oWP
Tb+FOuiZhjMCRDM305zD8NuvKRnVspHljnkFkRiO6WqQOAETlVPUmLTXCiKQfCLGLl52To0RNABN
4TItLe4/pbkf53qUgkJ4KcdFD+uGQu/mnhrIe3ZTuVQsPKDEFZDMLXSBdBHfgWOIFb/pTOkYmUah
A1bVtqPbyDHK6lYb4LbZRT5jgsLGjAPPhHmG46pXDuhh8outYqbwg+xH0sYJSLVCuimGYs6ZXv0R
Z98IIWWLIzhsyYPvW3KSJ6G6haDsZ+UaWFhOdA/tzSRfMxRdubFcp/R9uep7Od9Fo/IOKjjPfc3Q
gcRdmfbcEAnLwH+pe3rjZFl83rd5bqPYbBmFMINbWwAVGr6Oof/BPRBGv9pivnA57GsNM9ffSVcS
yXQOfkgf5uUWogFo1xOeXY7CzS3mPiRtLgV+UJ+EzBm9VztVJWwV0LnCZ8jX/up6W5rSbncEIRu8
YHctllPXdJ63+BS4UGbcD4Ngb75Ee4Yg8+qxRlpyZjGPp8DJ9k/0jCn3HVZO45UyKglzxt9rc9EC
JNobnRi+eMAmnnihaMGvfJuOIA/tGnu50E8pp1/zz/IzFW0hLGx4BSAItdg+sfmrNSDUUSyvJb5S
tjF7V13ydt8rQECcHAdOT5V+abmxr9PuP1PeSgVIaxyiaVtp7+DywEVowiDKfqTvPmy+mKiK6thT
nI7qLHLdD/BfEW2AOH0lKVLwvonNVCBH4e/i2cuaSUiFbyKWWQZ6eHSq9/n6tPSisHN7QhHPPFSx
Dg4AKtDI7YHNeiL+/jgwcTh7A5hOHNtUSi3MJNJUT/qfCzlo0jJJsLxCAbGhMbxDQzTCNwa1aipJ
gHXGsAtLAVvLiv5YCD/TkfeIcJHllq4NpjXX8BECWxEPwOrEJjuufGAWubfXa3bNLhNCMp2R6cdo
gBND1dUvTvtIR7oS0LU7HXBPmA6MlCytWOh/nHXo8EuPMY+84sbIj+zN8puMnOp2fb77PAmQF/I0
Q8L42cUgoZLJpsNUAxOcm47Vc+Wspbk/Ys48xIvuCbx/wrUpZSVNsM4ay1y1ZgPxTxs5z6uXcl9a
X3qUL7TxFZaDTSr4VFxcY1Z9qRPY8z1FluGwWuclu0Jo5Xrz+QH9iGPPwcM/hU/lbZT93ZKFKNrX
eN9MjISAZ6ImZI/RM5lYSSHctRnor/lISmrVh1Lhcugz+cLICJrsxv/L/tlh05o5yIGyYjuMpS3D
zYmyDm0tQPrwpa173P6ULBzKWi1Oevvx4Fp+ZvGjbXjqUMA7ik0mSsjuGYqePFu9jHL3i3Fna7Rn
ScvLDxZDGfZaZtCICBSKqzWz0phhRQrhBmHa5kS9gj/r1bYfu4rTchhKaocPMcY84i9Vr3/YGbxr
IFKzvqHtWJzMIpVVniO4SRlfpqKtHwLkVMX/V1ifNPKvUOns/ZV6+VVQq+/LKCvnl/tzLCoDRlhJ
leXl5xcCthHXtoTQD82AgAQSHlUV4lzFKBvQiMuSA6MI00fjfUK9wcC8HeHyvXDlpDeoRIKLmlzW
JqffGRxN3LfEr22CqdKVeNgu/C7id/kutyKluW2gyqKHczJB9pQpd9xFb24Kv7C3Y5Bz9yrfjGcJ
dIopFXgERi1+PQrBMqwcGw49AkRJck+BpbLpy8raGZ4nLAvCm7x43dJryzH9D9Ei64z4Yx8uX0jC
OLTqOU1afWcMHzVYzJBhsiFEfgV2vQvIe56RB2CMNtEA2nEzJwkDLXocue8C34zwxVlZdkaYjh2o
5vG8YRxl6oTC1PvgDlf5T2lTvAIhAdJL7kIiFMw1EIqmwvudBfyes4vFps5CrrCnd15uC6JS7zxw
/ftQy8bwyavIuN1EVpRx8iAKYYFo0xT+FSMJi3EkjoaEIksuf10Elz2/1kG6A+o2nEXlWWVBH+TD
eFXZUlOqsRFaF0XFQtsn4hbb97NQIdtjZBHNY12qjL8nWi2EJLl/cMe1JbfL1YATJsDP4H6WUAdR
EYb7PR9BubouMg5EVioDdqyqE/ae55yzKj+2t0AmmIYAI7bsFU7V1dWBC/X7jBsWMQ6PQtIUSZhy
eXr0+mkCNoc6B3N3RdkGzhIoVEBhO2pxJJC/gEF+KuPc6EJttRtlA8RXkd3V5dGJahrb+iBIy8kR
xKI9FRG5t6ZDn4O4jpa7vDw2yOtRfGfcOxf0pULSr1BYUeBJ6+0V1BolAOzCMzU/Ltv2xPZQ4yOn
rKlpq2q7fBY2N5sYFeip+4gzc+Kd4OulSn31/s/HqHzoCzoVSv1j+NUNBLqw0qZwqA9eig8xC6u9
LNPqa5ul7W3g5YBh4KPXbKpvZlbtgn3SOwPMCKD7Zzx2hIM2EOIUcfHWUtR9Dr5JiMf7jSBy7trF
hjGhHNI/064978NHcySqNwlkTv+8KEVVx9PV56l7U13jCZNWkl+C3ni3pD605Itnwv+K28D5H8RR
RLOaybTNQfAnwqeVLWzr5tAirAeu8rvsJdcUuFiMOoPCTJNYKx6DE/KqsODTXCVVHfkPdp3qwvHM
UPUokUubgduMjeVxCkn7KV4j/ASaC/0zu3TNiXou1KldQCDoO/S0Zn/AlZ6tahK+aiouo9CVDajS
Lqvbn7Z4rBDTem1oH3sWgyicSMbZCEuWqg9bjy0srwEBsWJL3hPlAdDMVasPaYgwbuP28HJ0jYxn
eC5Q5mTUiYx0CTTTq0s/GnHgC1RcJcQamuE8koHS/C2gZ8G8jXxc5nhcFm37O2sK6S0BhwBVHJme
FEkfImAqUWsBWwUarV1W1Pli2Kieht9PfzfBmEN258jQ37bT7GyBrNxWlIDjhbIXnaSzOPp+q1zj
4KQHsSe9VbUp7G5+e5ZcD81+FSxxVutpcplYWx3b8DCBRHnfPC4tv/2djcORKFjPKTDrLW0zCaZl
Bi2JCVzY/KJSzjOwV+y1NxfAoikAZwTWKfrByQELbteGiIcfvKUvyGrL23Iluev4Q7LxM4W56TYc
fGY5yXX7uJYLDp8K4KST6HMvmXSw11RHljaTONEUEWUhz/V/6ge1HR+Cc/2ESdhm9JqszKZ4BIF6
JPyn6ijHk9fZfYTjWj/XJvVjP/4kwDBk87LM2AxSg+pA8Zx4ECcfcikBLzIFjrfoQtVvhwY2qGmj
C9fB/5b9xT7iDp5nkMDJQIZgEJ4R8zbklS18crAObvLNzXidGLOPMxsGTD0yL86as9fOmEPiHz67
3k9d1FHa4J8BUegkXsB51+nqVeZ4cZy67e0uKByD6xBDhE0tft7VAet33mhHH1PMQhwLRk7KseuO
Nu3nQi0ZJLimarkfSgpOBc/8yhnRt0inLNTbNdak0JG9nB1olEZvdwmsVz67igP8NP9AqjLPkYsE
7Hep7Axwj7JJicrOa1r2U5MuKRAThwVHwnwF4qSRBYf9YqFzeQBzeRwZeEt/XBGSIeqwgbVwRble
B58PDgRcNDHAgiSBNMAekrxUixeVU5uNdVR4fIzi5Ybo1PI9437RD4rpmFUy3roFV0Iygj5TqXsl
7IKAcr4LkIQOQhRPIAYFL7DytZTCWb4gOEShlZKea981rlW4R7p8+wduS4XBTdHXcU+8I0T7ZuGg
MqsFwctNMoVexcmltHE4kTvy8ncA3GyjuIegSsrs8U2DWYDSN18sbejENT5gzK2an0o4J6OvftXA
1EpKZia7FLKOAdPxxnGt23w2DgQ9Wl/1xiShbQpVM+B7S0APcvEtyrQTVrzp3JcMuGZ3ISa4o+WP
BOE0T281Ox1vHX3en3DvGMJE5+Gm0uDLRBUw3o65Pkf73EYQNC/128yFNEcowJu5CfObgpkfkMJ5
AP0fcqKLG6zIAJOW25DZDieYVytieEQsobSbVrNtlJyTddfgHuQyL6hkmqMEKnCWRccwik+H3RB2
eCZ9u3noIc1gbQ7SIx0adBluioccmMCYvZQZcVYOMM/h3sRtdlFJ1dMXw069JmkxF+zl1ymYvSyu
OjWE7u6k6VNWWKvn8INQZH1iU8VLA3D8f3OD2VLUBho0r7fKiGcI9/Flk+KBgPEgd1KJsruWN0pn
rkXSjp+7oljaRa789E4AkhItyn10zK1ipdu29Cp7B/k8Ji1SgDqJAcSL9s9cslY5SFDYgZhhsV56
az8/Jd/CXVr6m28b4U5O3XV1cVpEVGU8Yj7Byp5NU5/ETdw2NWzLnvWedyE7VXikayqZkQU+zqCB
3Lxnbe2hGCX8c1F7+eJvuu2gbl2Phl7NZhaEY3rIVpAL2px5geVqe1mgdjKIUqDVw0SiTeoG4r9M
/jLHKJkyMYimIdPR1J+GLJUJVFtN10Nh22ZcYH8OHoX34/w9BdE8UuFFHY1cNkncFby1xufnUMye
ss53m6Jgq93jcIbTH5c+K1OrKWdDlDtS2M3m5XbbUgB/I8BeedV3V/aoWAOvxyS9kjDiRJqmnFAw
q/ILd2rHsTyefDs2oOFmg2PH/VvrdxriEoSiwmE5t92D9VU6jSX6Y4qByAOcdCGgvP9O5rWhdOsh
Bx2644qTCjAON+b1SGGhle5bcQG2H8iuS6C2kNWMHgdUZzyydSgwPeiJVbLFKcBmOKdUKoNJP9R8
EU0x3xvCEOwA15BIl0QgkW0/pIhdpSkBGa40OD3mnmUM5ZYPOloazRwjnv89+Mbb4T6NEpJEiKty
m90u3XZQrMeLG0PhZ+6pWZNvxuoFF9wIfqVNmVofC0FTO7Lq0F41tRZ3yfe18rtCekmtMhHOxJ30
ZryOSBaklW4nTF6oPowCaKciLeejMRCbvBfd9H0hnl+gpDM/gTHVqC2evgRsrN+8i+ySvP/a85ZX
Nli1ilJuwZi/NU1uuEdOutOJ0vxlINN/yXHBUQxz1nMBYBYaAlF+vrrB1y83TrzlrsuFe9jxuoIx
jMLVcQ5iaZ9F6esIs9V4NUOfC0svpinq4kCMxezQ0quDlr/koEcdxeSaJFn/2TwmY5sMw+lM/MZr
a6JqR9pnvtTcI43SCrD9UdplEuHNg+JgY0xfDintAmMy6FTx5x55hzTeGnV/iKnLvuEPcyopBh7c
fHpDaQ+egTUjoBONxQjkacSKwEBJ2WMG+Win1pbh18PAUTKm0i9Hrpk1etaDNs+x7BYkpe4GvIN3
ObfawwGg5cySvH67mu/3nyJHDMwGuy30268Rck7moKmnobRRVYiJ7yOkjssHOmHzxsqAbSAUVll/
5h0DgfbZfVZdpZLDdTqpFsXxUgwDIzF5ycwCOgILf1JHXwKCIj1/eQ9FBIemLVhRE+mDzaErG3uf
LcbDrpn5+aWx0NdHzYk57n6ncNwnVkHNe5JsCVbeq7xeugP9WVDRlkv19D34GOANZbOuyELCEGpJ
4p/rz1oDCDjvraJrcl9NZKDj8NU1i5ETuCnIgJahlNleIS/SE/En2xUy+1ETL/gjTsL9WJbI3Fep
6lEYG7YlHvz/5kDCnx0CQpNJZ2862pvE0MxIdOh2uARDdZVJbH0yjhZvpoe1oEEXQJHcUMmky4ac
8gpWyXEI2PxxjnPMwbbjitVzeV7KxGBjR/viuqa8knJk4cTow1KjO/g7kqLoH5GY+/m7FQJMB3CD
gNW6mQKt7+tSJh8FUBUSluwTUSLRf5fbMDGGuJRVWU46KMyOw2tQvY++fP9Eoh8vpIuKE7dh5JZb
8cEuf67HH/SsR6qSmgBtq78oXm98Y5dPpiFrJmAivjQO+PyRoTLroP0F+fjsHTM7kHkvG529hrAm
20Mc4ks/3R+ntIumQn0bh7KCgJrqGppjcSGKmDXbFLEHy5TVR7Nt+KwAYCt5bcbE2TpLmpnVJ9wQ
soaFDaEbeQdjx2tO7s6wcaLACgvS/HByF47ssyFeW8ZpR8pRIBd+NbD+Kc3OLtn4/cvjqz1E4IVY
fRQC9W6okmuJGJmDZgTX12ZoJlMhPbmiJIv6iGu7n6g/i6HL62wgzDSLyuyl2CtvI3BfahirGca4
63Rtrm3sQeucQkMSaQ1H6VnW7e1E7mlv5jrSJP/HNtM51P/Yi6sJgvobT19fC75mroAw/noTpXef
AyuMkViEnveH7COlHqj8SBbiBsfMrclNUlIioa/pcJo5OZonUyET2pRX5CWlav9M4ytmjRbtQyS2
DVDK9AkBrcokwkOrpeN6nY4d1zwPrbsK2lY8u2nR+6rePCCkpASOAXH1JU1kV8rC1E9EsBpRBAxh
3hu8E/zN8ZEBhpGPwPMDKxIcGSjul4sE7ivR97ayyqQxZt6zrr8dS0QUwD6Avm6abYGUo+k5GaF5
7/NPxA1vB1jzBOqb+e8pDQqGrtjWNTqVUsuNylsf5C9pEwhx1umxbsR1ADX4VI3mPEqDZQAcidBK
DCMi/hhQlHYy+V/ibu6a8IzZdhSV7fS7beXwIA9d4JRBwdjaUrbLDWK4sJVGp9PQodJDb7cJDXQ+
6p9PnzsZeLXiusLXh4E94HMbuPwRSOtE7c4fQ/AQeAm62qjO7yhIgSiLY4mnt5gK9GteY5flrGhF
AG6xoalaR1ruqUm/sIBH4n/TXB+6v9H0R7Kau93H63VcJjUPA51+OoBCG3VgQeR6sMo5fb91TkyW
JHfA1JDyLBSICSvgERngkz6Zrbw+lqIMrbdj0qRyyFpvphyUgREVZuNqBO/SXmXAws/ErKwtT9Mx
L0QC+6oIbUxcM0dNx4AUT0wgvLCb1fGaetRlh7l6rvrP77BZDpZ1EUk7EqlacQ6oOMpBjMYnuqk9
qSQJVfl6mrCoHPR+REx9SLManMZqpXd6bi0oS6TLpWwyFS4BCB4r3o7F6TSzEnAnnlyYFAfNcUOY
LG5KQdi3BQRfCnBTp6S7lrMGjHIEgWjTzw9vaUjX9HwIL4rWnMcrYWadatEgBTbYlGL9w7DQTG9w
NP8+MpQFmpxPN3ZCZIHBG83Rg/45XiTmILYaa0o2FcxzJpsyivVRNerhXtNuOOdG0NbdioZreKi+
pjCd/juaJxUnP7QMZFKwRfZk4Wu3cL3ELH40DDiUoa9dfIT8fZmlU+NK/yOXuOMmcl5hK616NmqE
oM75ptoFuvTcJLGYt2W56lbGVkLyKK1kOL8Na6BpNN/NK/0ytsL0PlzSPiuriW2Q7WNWq6Nvquns
nFHdVVFIjqR65QdpajrpTcNfm4UjoGyaC82Mlq1vrgQXO5fHLHyAXqOHUGibJnAtrOSMgx7JhRZg
o3PSX1W4331pY267vShOMMMq2XpGi4IdylgVbNQsax2/nQlIcHr2pVVHvzstvbXhEft0fFbg0UiU
PFniCGplxuPJ6N4BnGpZWpsgzlJN3HheH5OfMJzzwDXWI7RKeUoXZ6GL5SOa3xPSVHTK0FdYav7D
Oz3CgH4jImAxAwjtIwBQQesR+kEHmLx65Xteh+6Pf9/wRc/QRNaoEgL+heKNGI1FM0iKKsjFu72y
tuaYFzGREYARhv0E2Kp0WPSnmrBG//Gjyo6TILCgzY6+T7+RgEXtiVnzmNH4fNILgIHjc5haSGw/
kEwPC4gk3tUaidMvnHUR4rlrl1dQZ9VVnOKu77gesWe/g51GRfCvCT+qDwv1btD5K/2LYvL+4i5M
Xf6g94K+D0AbWqIxIo0mF3tI2Mzxb3NhEGrUOTt4Gqhr/T6tGnCe2hPA9vpvlxsSsN8YSadjVRqf
0VxOQoYK7EucDGwEPc2n2p2Q9Yo2zfU/Ty4OxR4noKos2DQHw1gORSmRmPnzgYhpR5arNAxWLG2l
pYqlKO/Pdk2EAS8XDPTBS5+YtMhpa+ZLjV+CBWm/D2lSooHUzr0i2IuXnV1KnwxuO+RT6mbQd6ph
b57vI/iXgHx2/CuLbwVfNZTs7/MVvrgaUAK11zhVFCYN2+m5YPbrtbXgXDo73mBn3BnE+JEuPwBf
Ww1QFB8JpM66kNE5f9mF6nn+OX69luDOOnmNwaIDJNKuSLoqqf54vYxPi6vy+E4tF0SsHJk/dh60
0k/0QVLag4AILdPpwVYKbbcNyT2cLDhChC7zqdJ3C+QVrAKQ5hK/4rDifRO3+jmcuSWTaS2fx7nD
WRvTCcCfmHUTK+Mj76GDROPhO18oHBOQbQ1zL+JWfYEdobRjm5Q3eEWT1J2K4WHQx+/SHpdTnah3
NV+CVMvtJocP4uZEk4VB3+JDofDA/ou3j2AAWCgJH0rBYhs7wxSJlXmFALWKwCNuTsqBaTU1bzEw
KNmb82To4c7gPChJNyZdSCMjKIbek9+7/Myii5xR1JTcSLwnyr09P4S8xS9O39p1ea28cVqOL5SD
77Z1RRpJSaKU+A1Dj0Jp4hZYjtIm+n4xroxZFU7uTWXiBYBOumkYRzqLVU5TYo/0IFJGbAbV+jcs
vKk7QmZEaRInuLo3T4y/+iK4kTT7jAZCjrXWlv+GjzjrvOOSV9NQF/YmlNHsDl+PihbJgksdtJl7
dbx46sDLDL1WpBjnBqHAxUtFPAF8kZ67MAFA0Cns2oBR5ja/Ux1+azKzFQPjsXFybVVQPZgX0wCg
kcKn/vTANSCFAv6iJdaxoLB8rMIoyigF9EXVAoT3jSrvFlFBvLDXzS7faAxn3DuYHGvs0Kg6JHDs
PMJ0PCLrZehnaoTLXEuvmxgJ4ZHIhFR6Ug4hfUz1pPrxsSKRvcYaBHkybSHQTYdjbElOCPK+72wm
na37dvNW9B8+tovKxaaP5im5iZaZFCCF40kWq7ieZebU2jzcnrhZjBeL37vGpmAUtDnite5W3NYF
OnMLQsnZYMSx+0UaMk6EDzllJq7i/ezhu4QlPSqAGch71gJRGqGWCIBMvcHYuR3oGv68HSZTYEnF
M4+K9vNc/vYgnEA5c/DItXPClEtr93xSZZB7zhaCczloYQsFujFL/TrdKBSQsn3gut7nLQ7uFQQE
3Up05kdqFMjv3tiyT+1g0k8mL3LFN9DeE59PJsQn9VlRgwHJFe3U7iA1f0t2r0khjur3UOxmCsb8
9IEWYFz4JvvLiOcQ2v227suwBYN0+KaCMPopLkxgPFnf0GeiJw9zKbuWoeLnJthD4SauaHzRxSJ9
slBp+dRC1a+qMt1AHlE8E386f0WT8HPPP2/fPFmP2ZfBtjvln69jSziycWp/MD09vJnC1cq8Y7xq
DIxCUE/2nOPdSK+1Wdcs/nm+4a33/MO7SnmQUhcBhfKyj1URNyfFrTFDVIF3QNEec6H2+ctX2922
dmzWLd4vscZxNp2cekrwivpDV0Jwef108AQLwLY2jUIpgHtcb6lYlfCcL3415YhPcqDPnmxDUZGR
0i1fWvS2dEl2f3FkwMj7DUeXEMSlPZYQYjfH4HFulpYi1j+wN9KEam4dEpxMio/kTlCXvznqw8uP
TviCG5ouDnDAy4me9zRVNzHZ/GmjbcJjmH19wZeRjPf2zorRTrwFBWXsSXzBI7edcwXn2dwFYtDw
jZkzMWRNgaxPgVchpeRrIquPuEq8sPv1dC2+zuUQJCh6D1WArc8+Kf6bKSKCSgasGX5rO9dIFga4
v8wvSIxoMANgj9HyyrTdykF6PZY07deRXEtU6SEDLv8QFsPDxGkFigwtUHrIoH6drVo0EIN1WI8j
KeraBkm4QowGnCcASwwYporrPcSfWA1CewmLExs+1BJr2mGe4Ff3z87+dAHcWaoUhi4pdr/QmyV6
bD6Qvq0+6B//4T5gmrf769EW9+LHF4YxJkSB81428/nYENaVwoRhuIcXraUr4VQkH+FwRzXbm7K3
jCli1UgSztES00bTUUHYjOgioP6L0FG+Qs04xYyfBN6Ek5J1D0Aoz+DQmA/XmS4CT/PtfUwuPWBJ
mE09TWhU5XZEr1Xp8QtTAQRrqO1eVetPI5H1YF2dxvruHEajie79TVYJLS1CQTKxbb3PsMTAHEdK
jzOdrtc8i8roqsFYX3xHyfnXt8nNtx0bqvYIezlPN7u2aJ1SGIpzkDliaTwwoUq68p1BS0FLk5GV
o9XPIwE0qg3hTy2/lHQzzddLRQJEqWBJ/ApRMtHPCsvRgVDzYsmDvX7kgQmYpoiG6ftUcHgE82RC
B1ajrFAG+vj+CN4kUf8Kw237Q3OSnOebubh4458xu6l+RJy9X7baBp1rLwSX5C6nONHympiRwOKJ
5Jy50gJ1i40aR0idk5+azSubw9EfPZVK/5jHSBxDxFUO77pU2Nrc9IQC9SC4X98XShWuiHKwKvrn
jyzpgwGUmRUP8ALzwEEZ+gRUwijMRtyooo22DiapHWi3szu9yOQQck/M8cMrUqgmEdNZCJXLeEVY
+rydOx8mGQWX5ek/z2WWLDWPO5DA/Ni8BpGf1mpzYUuhHWebmmO3FWdNqf/ey9ajKGMkhPi3ykR+
lOM3D3Ull/a5EK4AlDsrGDAfqRaKqZPfc2u9AXTetAMgemGDGcMLj1Cxv+d85JBGYRGi91Oi9mJE
IXPBhm4rkIQnJPvd6Fqihp//YXcxkS9X8w7Z6ijN68RQ1dNEb57yxd0LqVWjvoDmM8bsI/GxCgw0
J/ohBg94s8u3ebOR6l7JDrMaA6a2dgw86N7z8W8XqhUG0tJwIi6gt1t6jh0wAgnf0v+qVElrFSnA
DSmU6NLvqHJhdWXDAsevCCDmbBo3XoePgEnJ9Ttzoc9pQedWxIqcZjQ7GtQzXpbPaNh7EgON8bVe
E8/MRsi4YRO/nb+b1PY6xWtRNkaQT+S2dM6O+bGGQC+4liSr28U2byQnjywsrWYekzyILkHHvqHD
0RGS1iCgJ37xxoIa+7qxluw4uUqdQd2FOadFGGqRXU6b/LyUuSOAcbHzr/uaDiFgxcF5ukvbibiC
tisExL2XHd1Kj+Y739w8cJ8XmxlGYg6nU4o7Q2aGG77luBaI6mzlNIplvaXzC6OEoISKlgNG9w+Y
xXY0WYvp2F5Mbj4jmoF0/qM1O+sVrlY/sNx96Wangh9QmjuqdK+9m4+DZpVeuHTKOsRG63TzCPCj
a8wCpWBOwByZAlrFZnnrq5v66oQdlBPpJ8f4ktBxtluNrwDMLa+ThxCFa7JDAP3qBCX/spHOBnPw
QHJacF7isx5Rs1VAUGj3aON5HJw99sYavhdOWb0u9xEyKqGcjQZaVCNN/0ildZFutOcP48l/vJs4
krMpmu9X9GPgtjE7I9Sjkuj/dMaJLQ1nowWVMI66DXmXe+3Hxc3pcD4XVCTVxzH+Z01yUBR/QQZh
4pSRl6oOl0ki5CAB9QzjzneVOSTxcufT9Bt/iWcbFqgEsfzZVXmVEIe4qGGBXSF83w86QJRnhRHF
NxKuxC9LE1teNPGwiQodBMxz6OX3XMp6cafnNMH4e6uwoF2JfkMTWIfMjyMo6xrwsWe6MqX+CMO2
tAuKcdnr10QiDJi62R+PWKF63FGu6o207q/wh8oM+l18ElyiYIjYHJgPzCBAo5Losn/u5U3nfpfM
ozL7Oi27P1BUHJP+JWl1Jjs6qkfZf0LLPl2r0KNDVkz8axvMkRPIS7XpQCmXu8xZpWyIaylGiNaU
UX8y6UDs3njob7YToMNVV4lfV9cdorghZjVS40+fD/1ZabFZGhw8aRthiSKZ5Tgau8NUeVieW8sN
sTvXcvE/FmXQCPlXIUAcDZ9Da/Y1qaiVOP/djHRhMSARiLGyLIqqaSoa7inXCQbifnjtPcxVyNUv
FMpjDCYPsihn3dRGK1r+87cvS6G9vmoB1Mwdj2f3jb02JGnmuKG0QGaoWUOhyzjxzIRsq5gntkdM
d4xglzenyb3+LuTFRv/VwgS9k89Q5bvbQncoCLp2oinDp3cLzmpgRl2gIdZWVdD+pof5pGgcxF8u
9vIfTI4+/ExhzzjfHJbEGdOhaRwNlIzbC31LZ2yMdzfmn9bNptDbn9jQxR7Ba9ijT81+tHst+LYg
qRcbueMpMA67owMeXPTZcXx8/i4qZ022vd7YLnGRC2sB0IgjtVUV6M7TikuVYsyClTYZ4R3F7hdZ
XFc1CnBq7HGq/1irlC7u00oHIJ16JkoCvratRx6tYcp7QNiVXpRHLfSv9+dcM6c6OTFSCY3u2Kj1
FTV4otcv9Zv2LPZ0SVnCyWV2vo2J48CBc9wzyuwynrOYPsJQIWhQJyFzE5vtGK5j7LBZ1SLieGNR
iv+op1mx7BKYljrUQjpItc3UUqRZAdMlXb8/phoD8WE/iU6CTMMxjtSjLf7JmEwi/+pcxrk5KL7g
hRcSWdNyoINV1rIUTqIkbWoDCtcya3oeopBZrRivIoPteC7Ne9tdWFRrpVKEBZFAeBv+Scgd2n/k
HBueTv8gjeb8F2BpQf99z1+hVDThfNA/2Hpv+xNvlxe0zuTTb78GWkIdW32jWDX8Wb0Fpe4djN3W
dxBRm9Nl6B4ENUlbvfkcVzUEKnUz8otv+EuxDV4bk3LghC/8IIMJL/DDEvykET9QoGKmHUGaCdWf
WL5BeyjQLF5PUrJ5PvRz1H9tb40JaF73oX6/eRAtLP27JzqjTmM8/h+0CE6P3sx3NQOoR2zrnSgw
MjFrhriahpa0xPFydG8RhDgooRB4m9Uh4SFmU5LrSUty3DAG8FnOTM4ukSjww3TGBHfr50rVdTw6
2WzBliaLCcpVXc5dbFU6A2KuhdScUSiqeGK7EAHbnUs2G/QGTiKMf/Nk/tyWz+DF6nC9fb9HBCeG
vye4MGAnqzJxhcEFnlIuM8PgZLhCfIq6OjXaSzBiS/gZmwf7TtjzWMsbbGcu7v4Vswy0hVGdT1Bw
fyjHI1TopsOk1d4CTYOjhkAGhEyb34WZJ1PF0dpSuQbttKKyzCnZ9Qt1Bx9Yst82IAe3Kz7Oyzf5
RHqcsqAizdFi2hOmPauwq75Vi9ElOkCapGTB/ju8QqSqSy5uGVahkqLVJ5x3dU0q8FKJIhoWyJHN
6VBomE+yYtAFD3YyYT0uq6SHpmdOZ0ydB4JXj5TAL2OdqrWl7DBLXE9Eg6eFR6kWwgaYYvxWfdhc
F7COqkwaB0iWdh2K6i+4BOTB13j/6gWMitXp1Iqhayje51w0gKzKs9orImAcXlfIPeqFaZrF0BFu
fN/94GxjAfrnookyWlhujmgSCtxyFje6OjZa6WVO6st4+qq6RmhVDQrZigGLAnLpQzGM/UlFbxal
UBYdyFA0smILA1O0tHVRhSG9aAd3HqCEIdqD7bnVp0/iUiHYzisQrLw4e7OO9VSEOREQUvj1tsCn
xV4NKg4HG+WoX3+awxCFT0QOkxoFMZKMOeQrmxoESB265OLPRwkguxsnpv/Odwep+ham41TwG/r7
wUUSTKzCcEm5VQvoGJfR3az5HHbW7iRylOf5c0iHuHg/RUNg92lD/Io3exBvIj6q4bHUE2jQSIYQ
8jcZuwWEfiVd38GODCqvkoqJSV8bU6oHq5VMn5ECay8B8oBQFhsIT62wSH3QyyekynNzKfmwSlmD
Cezyv+9ds+UuCoZPaOi3AcZMMlL3q1fnveap5BF1sdv39OHsRptVCFmiqqbb/z515zJdHO3J/MxN
Bc/StL5yAY0ovMVFL9Bpbwu1fhCRPansl2QvmWTT7pIQfJ7kehLVfU+vLUNfwUgwU0u1bp/bB6Rl
qzSKMudhWHW9psBIHuLEbS+GpKhnCsBli47sxfzVaRIllDQLIuJqp6PcHdoIqbLgm3d4NF4dykP0
bUluybf16nITRc0kpGTrIn3Ov9yP6jMEbWv5sn5VuVPuo3tTG5//i/adopkF/r9f8Go96ZG0FtF9
z/Fuz1m/hLjLHqIsnhTN9WwruxAvMbnjsJei4xCHxlqGEpml/PlsiS+C1uxxQ2cNwTBf3WYxLfaU
wKqMqJpUi2tD0/CP9CxNaiWS5bs0FW/JonP3QuBF6P/o90iEhtui5t5fj3jEtcfDYWEy9dfhUlSD
iPyxA+6fegY5Z326yaLgB8NYDX8g6nLvb6etapCyTHXkKBVQt2AAxDfpPMA7dYf4T/cBYvgSRLWu
p7sNIeeAks+e/Dy7QDBkVUcLiBcaFRonQsgGdQYL96OMFTyS9Ea482vM2w96KZnS5qHfEBth2lUU
aWYOINvTjhur55NdP8/xkv3MqZqpoVlCxRCiakP37uBXVu5ScZpZixx4qhJU6W1jsnkuLIA2ILsQ
Kf/kZVSPYa9Gz3qns2PPM7R5PJ20c1M5hFC5JqBMwp/TPnxb9wkuPVPqi3crw4vwHSKcSRGZDXmj
g94W3hcGdfv/d5oOMiIm0PBqab6Uep6pyL99StMKBVgOHEKOy3qARL8ZpCvjWpn+Hal4vVikDZ7f
NbFNG0Jr8iLI+9GCWA1IbjcnWNSkCu1N1b1f3XNmoL4XWjbzIDpydF46zwnMpaz/sat8kHQ2JfQX
CpxnG1r86cJcs2T8lwCauiACrYt+61cNhd2q1/9TQaxLb5KyxnpgnWEUnEwQppDoCClIRnZYE88q
98gvPdslk02KibzPM7OkkGDxiMqch0WNMy3h0QTCWwEfmaxEpe9rAln6mbkBqsYZeMlaKITp2DxP
Q1M5Sz0k6xfbiLSNnlssoeNykDAs3iZ6WCIGT7UNVHFQA+YzMCkcAOJuq37oI3ZO1bZfOjHA0znR
qCKI5XhuXujEBsktYWqgGdtwE0CFlF7zDpdgNqzT7bdkJ90ufZBIAKN9dZDSdD7wmzN4+GB/60Wc
tzkdpYDfi+ssj9HVY8KDUW934rGc6kLoc3x88oUp1OdmYlIsb6Z5swSOZUnQBjItHr0Sl2ukKiWT
a3U/g+xFXeErQdHzbhiZxTOYr4kBLZl31x229TJDEIb4UWpOB9UsZvRNtmkc4C2H6/HXJ7nt1F/y
ysIKfO1Tf8JljwHBYUAFF14lzH/3Fq1Cfqxqr3ejSHGX5EHtvqkGgVVwdhfAwHNjOcq+DRBpQ971
+kAJ2b4AqYzo/dQ3yriRFU0E/hYtufexwcIcUTbOWfvci40LRLzHkR68DTia7evPNwMQQJ/jWtsn
qN+4Fa5fmmPFZEO9XLzGgROJKBnJn7a7ZHr40uFtTCF3JosdS21qNaoo/6SIHQbDhQyu+/bDcTEJ
49AUS0b+IMsUcaqa0dReH2r/FbMj5j72vQ6INgVSidEmNSajdasm+jF60N/8QUB2pZnML0e8dpfV
VoMBbqm96aV9KRVrswsAcODUP6vH8HEx4zo0/d8ihjEyGHqFkT45I3j6qVWWysijVtU3IjXxJ0Ve
PMhpcmGEw9vZF64LlL55H21PRxR/6hDOi9IkKjeT5vOyaXoLqskadQOvqRAMQ5jAoq/O18rbhhcT
P0In6b2h5/lssOdJL14FJ6/1iGfCqxx0cTH5gZ4oAT531qCEMeK5TQBav4JaWZrP/F5sFqkK80YY
CTHjE0OTJhSQH3FJaxneMhmBqZFU3EaE+2eEe/efIAi0j0K7NVTf8cHT57juf71fiW84foPc2MyK
vMMcVYCW4mcXqIPRldulw18lz71rpEmiq+c3MZJW1LpcIhHr5pwQeUxJZpsxyWj4kejtTLddudo0
/BeUbxuFnJ1E0soAxRp+kHrMTtnPZXxi3wchq4ZdInWMsJuVjyzecQ/KjQA3wNXWjTeCDw4okelm
j4WoCtjiq4NZUxKjlMsFGHeoOXP64bRuiw2nX2j9Fwa2BFknYlWShrI3YLZH5Eer1PyAw4sY/Qtg
sEKBM4xNqeuSwmuLDGG32xfwAVuZJcIj9tsqI5pPQ74CuCUYKpYmB5aX5tdXmEfu1dbxw30I6UF7
D9gzzEibRde/y++BVt7XHa3UBg6HowDYWepb7OYpg1Sprm/wCheURPH8b8M4IAbHOA+5vfPAY9ZX
oiJMpcR8+6dU2cnLVNTcXHttLJN6a+IKKAbfOQoTmM7IhdXXCl9CgWxxLMfBn1TktY6De6rxSPzV
xccbE1o0EcDpTsH8JCiVajhLXEB1KDJKVU+IZ2hk6cA91cPKHpMzJbQLQTmcuZuxZ/EgMr/hplk+
Leh6gZt11m8d+IU9PlHdkC/FVFmoBlbUJxBDnxDyqFnI5DeLZZFkCaA8JcgJnWgiv5Av1gSkfDMN
YQp4BbULTMiJkUgjtOcfwlu8iJOPdejJX1izV5Y21iBODDpp+Du+qRPAVOWZDcWuHUfEXqMKxhFd
O1o9M8pK7rAKcPweGpI+kaZWAe/0ZieaVDuhmflSslN9DuKWBKZZNTEXmACfYRWZ/K5yLBXtuD0Y
91iTa2Teyd51M1gLZMebmZX3zj6vzAwqj17/KMCaj8RL9+hfGFTA3rtxmVzdZwNSxH5qGKieeMsa
wI2l9sj+iFbWGhY7ZCHNj1T8++UdmV5k/ioiy075LN0+4wyagVX55xmHTMf2t8c1aFeUxxFJuSPb
7VIlI6Vby7ANzS/jLH+2n59FQz4b+X9O18f+DhOWSnRJP1PeA6JrH5kns27AvhmG/cjBSiApUblr
vArCc6BHX0yT9kv2CHUOgCI6V0pKrllUHYWpAkZpZrNu8W0+NklcaANT5ucduKNrt9laSW5/yKdO
JurWG8siJ4iN9+EzuPh7nJ5OUZ4uwEjN1EPh+evJX7QZn+WSg4CdSf3D+piKYxoaB+OUnlBolCtE
KqDWEJeCRbhA9//p1csmeNlznLO6zJKP8Cb4w0hX3QM0gx6Fsiip6mKH8gGtlg38xX1ztm4gYJK9
dndiGCwpAjh4JA/aAZ87Zt3nc8CvQ6UGaJlDFegRNJE5SMxsvPO3l2tMpbKNIHPUeEAKqwk3jU7k
GnuHfzy+lwH65DuhrDWMB/eyvt9IoyWwU6WQWFDqosylmm04omL/oZcc+C9uFVzOqiYc/jM9+9jm
CmHLbPycg/Vp53OhMNTDfJnxIkylE2Cezlk/4GJ9urLyMccOJuhvSAtYkmd5kBtnfywALKpXdcHd
LEPb4oHRjzUTNo95J7b2Y9evetUv+GzHsTaD3XFXszFC/kXXNbiIJDNHmnYoSabY1UgFn/stzIhW
aMFjrubztmZ9tFIlTSB5xoNB+UVoBTs2rrZ3v/R4G+SgZVsQglO1RKNoZHz55mFAUdWo73/aOzFg
iN335u9ln8JNb0fuWNI0vsHqV678QUlhptHDZ+Tk9L44aiTBXzkDAA9mmtg6cHQgp9EbUIW+TqLZ
LRCe600xtED/id2d/nxJN1jl2o/8zxMhWI9MKjC/oG7xSsGEtb9SHvNZIoPfn9ecOGNy8GQADHFD
hUAa5weUfR4JljXj8dKOAJWNAhqMdd9aYYE9RzUMCGREirJrGsFH7lfA1QFOl0qFr274IxrRSkvY
wep80mmXwToB7+zzqPzgMQYQ3J+AEWbm4n2RBwuBtITi26s/fVr/1EqBz4hBiq1EoxtrTl996APO
lgKze6KI+bOXBZ3P3fANDAZn9xVOCZrwV0XkScsxnw0gbe9Xo0OJGRJDAbXT9W+x4NeVr2ixcqAB
LW9g2clNvS/3TpRfaatukD6gaVokSY3gmgvfZneAmCQUHzz2kUXn4D3uXaDWaj/icWGPjjrJpihT
d1zcm0Jq2uGQecWZOqHkWPg3lAx5U0JZst3YopGBb/lPQ1Z8S8oFtUjepkOHvPUUzGwyD8+GFsep
/ZFNw1NO9b6oGaKBY8fC7C7Ct/MyM7MKqAN1q3fNSjM2iruEnxithJE385kgcI4Mpsynv6GWYcaU
a/iu8nu/42yTI3JDsiJf8iexNdBiW90JDl1vM84hF3mAfft0lnBCG8HfQBkVhJQxBqZzNVoD9awr
jCnkiUOX5xFpG4nlIRpj+YNXu5vsK3by88YL+Y6eGdzP5C1O85Mu8SORcSPuH1Fy2jiJIpKJNvZ0
8+sPlx8uyFk3qYWk3oU2PS8hK90l7ehoqkOzQfSHj31I6mHe/YOu7YR4uN6P/aDKebl3GAkM0us7
fyYewVieMHlUenaoOCNZ2SWw/7E51bHi9WLedvFxhmr7I3PPeH29eq773lgSXU2et6ZDHTkuNb4n
bqHkaM6ko5HtTfsClQ7eoa0NLkV07rOd9WjeUPW5CDPSURpHEHvo+Sp/jPFHD9SuEgCRtV8Pba8T
zSVB24/PO5Ybg7fsBkwyvdgesyR6v3ph4uZvAsNnjyo4f/XHj3xMEs00PZpEdqWCF9IJJ6BMd4JL
fAG0gBPshtR1hHtl41nUSjzvul0I+rcV9TGk/vuzwZK5gVZf8EEG34je7dGJz1c9tCA/5ZUjoWt8
7sHKugAY0wdDAamlVlNQF3JjF2kmI4+H1xLSVAPInAN75iO0KbILHelloNiblFAD3u242BmOhHNU
ehFflL1tllwf7T51uc+MefEtCyzlY6HDl8IEnHbf3R3atkrOhFC7NiUoN8RpSb+eW2ptWENtyyGu
DLrbdzO/U5I9u0bT3fXQ3ZeJX+LQielW3d2OJoDBUDSZ1hSxP0T0tHdg6k6S4xsRx5fpOGkLXc51
CxGtQgd35/TtJ2ifDZ9nPyUaTgScfxj3K+lLaWs/x5S8qOSIq76jh6uSkuX8+x1jjM/lyjZ4hYL1
eef1qYsrBXVAm1pXV/pjPHhL3681C2kli+cYLFGzKRXMkukLRFH/lP4mqUZahlq6uUPgNlf02Swh
WxNmwLCruTmXt57+nmkh0i3YIBig4eJ2p128WIDbubsAAvhu5vk+quEdw2lGiQ4/mLMsaWH/Vh63
zsQFFIGYbzriAf62AsQfFo2RxKV7c5NYLTyE0VTEYK2vRnfAxbig6K4VSP9BhuhzuJeyVeMMrC4I
mn8vMicDwRBlCRsc7YcH90fOLYR0WiWNO0bhy5P+ZgBrqotnV5S3BClH1mlNtRUzAMwQHQNSSNVg
mnkcAQLhMx8XLQGxUO+oK37dtuotJpm5ov8RWmPmA27YHjZARmmvRDPOPoCmVw5IR0I0gevj1Ry/
gINkt6axiiPebqA7MccS4r/noWT/SFLSUKEruGGD8VFAxyMJMYbGBn+JbGfe7hNZq/p5GdFN0dfe
aACTfqjRQHQaRB7GDxsveciJQBq8JzIGbq28g8cTpWkKvpNQfYDcTfPadA4c36Q4bMSaZdvjRxfl
M5P7XT2GkClc5Si06RLLa1Aun10se9n3qJcSxZ57epQzLcZuEuD65UoC8qDCgvxV30v589NTj1Rp
R3EDxi8j9WK+iQt3109mDb8vOZQWu8ar+KDEWmJ1zGi1rB0fUxqsG4CWjVcLBBYCrJtHg7QXIjFl
+pDs2dggh5mQb/6VYmWS068qVN58un9SM7LXKpnnvozj8yYtcG7GgCMWj4jAtRBdA8TTOIbM+jkw
8/S7CejBo+mAtdEwJ9iFMLnbYzcAqSiBXQmk2KwhnYh+JoaxH5X29xgdovcaOn4aIAkFJVYeyphc
87LxjCbOygZXaydjT06LWQzmccLUPfkH3MTZIo+M/os6OauChGZwLXfc4WwcVJcNArGsOoTPTT+/
EAhcgHMU+YpRadlNWSA4sX9FmIR2EcoH6mBB4TGDHNEAXVTcQ8vvlRAjAY0ogp2tmbEdiSuyknLX
NqlBoKJF92MDx6b9QqaFEp9inV0KsIeK5Y5h1P/pjfGcAmBLQTkP0S6WYrY0UXBiweiLUITYb5pD
CiJRf9VJMwj0qMeC4hFQxmuV1Js3yKim/fs/+KbHvGEsXB3nokhvCatle1l86WF3wH8J+FRKr/9K
DiOi8L/vc5FarHEFTG+F0qQVRNbyLvhQgy+YBmYxDACIyG1Emh6OJHItSI/tkJeUTNvBsCMa6aWP
BQyQkycPthgeNw/OySFulXnJQPKRmBVTnoJLNZ1bo8kGkUZtNWwYAijl68UTk9fKXdzRNQj9pd4d
jrtkGEBRIPRNTaV1Xf0r4Dhjoa98PsBkq0jlB6QyvnDDL2trP/hp+CqcH251MILnmg4Y5H6VYmH3
Nxf7LEMiwoNUcm63ZKHqNdbnLK5DxFJuEkPqiA5rcdysEVSQ5fXTgkkxzyRkAL0DtzC5xp298jJP
xT2yqcDwyLB7Vx8cEqRmw/pO3MgHyoEsxUzzgTS8O/fTrq1s8gLBB2N20i6FGD8j1zWVkY5djhuS
kV+iKS13IkAjwiJAfyYTQIaM20WwKCnlXW+xJInxA/kNTtbIHIjuQx4J7q3gkb8gAL5M7f91MQuH
9OUnIoRhPyBijKk+xnTs1cBW/3Of+j7KxRGo56iPjajNew2ftKyAfxsCf1n9/Kzrg0qh0lnxuXUg
eTJ2ZJ61Ii0EnbxD2UN6KGSK/6jWvVlRsT0CUwibiBBqGnFfxJPCxqwEHkOT0y6lgxH8MC83NIUE
QLoH80ApwAl+8g9/OBogsIuw/QYcXXJnFL2ZZJ2sYGps8ltRkpgm2VBbRGsJEH54iogBYKYgv4MZ
Hy1XNy+hRmWXH+c6iSK43OcPVyUNjAn87cijfEnqAmo4SCbDp3D7VIHtgn4JPejwGRect/q/Lv+W
6RCJGTAC5Zoo4AmVvdwyAEGSLoB8BHigNfS5uPE2iYwnIwRIuRccICKqolBINK/OZUIbvpduMhPS
8KPUMrwUn3aDxqRKqUXwmu0e5uPSk1STQglaDu8L9dGfFdc24haxsTBlOmqtvFMqUtoBTn1KDUm4
7E8HgAahmQ9Ho3cJY1PSIlpZatwfCci6+Z0Pcay5Bud3IIoIERVRRWHRkkYqymGiWfoPYw2E+lYc
kwt2SXQaKZSXg6UvAl7rpMVTGqBzN3A7xL+Af9hbNBYjivXZLVUFVBTtRNsW2FSwPzq+HGAM/JSy
N9oo6a7z7Wz6MIRewmFKuo0fSM6wfiFULYwT1H9VaiR4DwjJE9jxl1Ei41QlFnDkDoqn+g0B6ylj
WrwnwfdBag/1BNvWc8i8sS808Xrtfj66r3ItgzFBUCB3IS0+1otUe04+LGqiIpL57stpB0IGsTQP
sIAAck32AgxRbWRIwt2elT+RBq6vgSX244wrKX9/P9dTUjkDGLL+wOKz6hq8h9PgNi0IxxMm84wT
qyqrbW3qxOkQQMjMUsYhIpL0frPNlokU80/jBjq5ki50u8DSPgM9rSi2Jg1gWf9l0M5db6PajYrU
diKXT3nN2fT11+AF+P+SfQfuI/OE8mW++6ImwGjH8fCSv5LUElzFaw4WFIO3u1/1E3/LEhQxMIeU
z6mlIhmIT+ftq2BTipxcj3wKI8Tx8qTm98HFgyD0jwDFhYISjO22OZwZRRnzdYFFFUX2cscLHXHo
lW2N7wMkKTpAS/kpSZA5jXstQmgGUL+EHcQyNyb0Khf1HF+tplqPM9trVsOoj1ugohvJwS1jNLmB
0uowHoOsQJevC6egtM3UD3E8TSn13pjwI/M2UVPPI8W7feQ7km5LTU5aUnr1cV6FSvxEiJG1KUk/
NsiRsPwsNpDPNRnzHQaGx395mKOu2V1h13xsHCFCKZac272T8+B4rc7h1eRuX5BDpwk0eY2k7VeE
HbEjhmxkKfnkqglpoGSPOU2dVquBiXzhObLFZwDBLIkzrNhJEJOUZaJhUcE09zRF27/JKvhmQfBb
3p67v/SjvksxAEagunH4KoALi/XQ06znsBnuyoy8mZ7ANfBHFID+dZYQK/89AQOtk6bpH7FhqkrW
ArbK9JZM/IfzTpLm0n8K70gKVzwO6KhGlcImH9zuT8T+TVk/q4RgJ1prpKL1dmVUx99kUg/0/+5G
VRhwn5NdEQpxMBQWktEcx0j5rfEbfCG3BqRxDx+uhfK2lmoYD6e1wAnBL/IL87dIAhS9INtT9X/y
LAZ5dAOVFNwzxZZI58pQeA/gXQWM+tn7rrYvKRc2wGoRU7E7m0JjVtWhG61fcEZIU64JMZ0lkNJ2
8yTXNbJgpFbm2LPscbo/KDvvhqGMmcRYcKP+qPqhm2s09FN6wBqS+n35hVUiSWbLA6CNUBXMzp3t
xBGlqD+m281PeFVFRL9G/1EUAgbqeCB22TKLhX690v+8djIKlGqrNGIPiJn8D+QpPLBC4NOxsaUc
ge/3AnHKcKvRW8Rt0pu88oAipLvjrCHQ47mFTvazpmFOpRkH7Xl7qisgmoLaXEWEvIJwm5tMuFKP
+MtyQ+olwwOw0nhCxlNaXarkjhm88PABQhacLBXNQm3sJMlFkThESjkEQYY4B3NV4fyLCql+TQa+
PyO9bEnoSeOTOCxbejQThpo2n6Vql8rjGaTeYdvqQBOpfaMUW9udHVx1U8lN3Uv4lzXlW0WqVIRR
9K2+AT3LUkunPEP9XfsOybij53yjPkpGlhomoV7/kbhybINIZXpfCDu7lp/yele1YldYkqdiJX/P
Tqe2ZheAyP5sj8kVfJhazJAePeDmR0TfbEBfyXuDU3nsnhjL/ElPtF5EIvXxj3tugKPkpCf5YCcm
aLQAdfhAVydrHm0Qz91Aib1jUrJBilGnzfJRgdCIkkaq62pSIWWBEeNdnNZJ3PxUTbfj00TTp/Kz
SsnhrK/espP+zrSvqtzmWBrp/6U21FvO5uxWTsSMvit223vJ5qyww26exnNhkwrARlfFgih3+7kT
BNLNuGDFLbruSdtfmArvZoUKtA2v3FlHDTTkZ+6EMmj9i0NAOzijp1nf47uCSKcie8EerBYNFFWl
ZlzLRI1eKGM8IK3aEozLK3iW3Uuf7xvXwBPnpanSQX4bsdPfdeG0qajaDrP9C0+eYw3RECGQoLJd
pVJCIy+2LA6KjWo3JRywQIZlaUXjTEcbEuCRTmvcwtXxlbZnrZKKMtNhZhoNDO7zfXAdf5rVMfEB
55mKfnRi+oVzP5e3ytaJs7FZiI/Ojpk9+iBIrsw8dHYca9bQSJwJph7Xwy94p7K46O7m+jOm8i+v
pmoJxKlCxY6MxwanJZPc+FS4coVytYQi67oIwfKF0TR5v28XNZVe74SeoClJSFDoZdcR0KTmywUO
iT6BoB7Qog5aaRMQuB3FKuj+r5Jsk8BaATVDFwPGrzdWH/k1gRwLaLqHE3VEefwB0zurrOtx6/ru
FYzEqU8w5VyGRE6jxZFSpp4cwUhckvkTaotxbb4yFXKFDjsrLqNbk9K19c6hPne8F547RZiCsVf+
V3Dfk+LeKnctb7sqoywVHMKjvByWhCGjYz4oufVek6vukGG9G+ObM4L94xvea3vxqy8OPTQXFEan
ICnpFVhLeh+AzrmpTlcQNxprFKD+ZA319BhIWv2rbh5kxYpYGxcVgqU9n4QQoGL1xOW9QRpi2m1Q
r08SgEd1x5SIROhKL5rA0+qdNHooqQMqjJg9Y+zecoJg4Gh3qgUm4CX7sTNkpqNSvD4LcBHiskpl
huSQDze4k5k578WyaaA0e6fYfeF3h+LubbH/LBXWZ93FXawbasHSVCDvnzEMvf1QVfVTM7eUHI3X
JhXOVM4MKAHVGLH76slFO2uwV/TxJlqGEDuax72WDy1xG+9Ic18G2qxvQzGf1P5cb5uLBOvkeHsG
wHwsLg6e18ZHC2JT3G/d9mPfeIyjyFfiQQW9SEV9Of6V+1ZRiUaphL39jUFxQLmmTOuifhho8wCA
2zMPTnVgAyYxQeES/Sl3Oq2qSuj8DTwcsP0CZTgFtupXeC2zaU4tHvQUULMOBQ/mGYMCbve2mxVq
bFnxhGnJ2ztzgLMyjtHwyAgWJTmO3m8WNf93hfylbBLgyR/OoVllwGy/2dzws9wzRlJzbJNF1GN9
tIt9y9Jk6VGfHAE/C4IgdopM2WZmtbDgRuBrjN2stbvIgslDQGYIcdxtxL32kg6D+XPLravsbCef
7g9LephAhVd+2NArtWP7l7sZLVAXVFwF2cN+uVUojFhLXAQwawBhDuUW2Z6y/it0Kvf9rlIBLQRe
49upBDRcC0ZWtbJ2XfZiqszH879DT1Y0WpWxmYwGcTsu6BhXhx4gUIdkqlV63Nqn5AglOEfkIBJr
EVZFaVL43GXgP5sZb+BfvIm1HgZ3pRFUaH8M7w8zwWFL0YqBhn3c9lpokZ4/lx+6VIxhAat4jpbJ
TCATyFQj/V1PFtiRZaeorccQjzoYkeY8HwA3PgSG7ioYBPVbYGI+/lhSC5WgnaPR+wZGjDvybQQ9
LZagaTB+lI/do6PamoeFHr/81kq5zoQ77lgGQ2b+MbuiXu8hSz3o2igZZQBb6IQ6S0y1eM+sZ6d4
6LWGBJJzfER11T3fbDLRm6S4zQi4Locvri6jSoaGubwBxnz0wrkL0WxvVuYKZV4O9rdpBUvpaL55
vrsleLxEF0UogImVYZFa7eqocHNS3pOzXsbnmPBR53+Rdcif6qqojzU92OTzZYeuWXJLY36hgCCx
ud5LNzhKbBthp9hlMWWdhj9dYbYJFiyjYtKDTQoy271ZxfhJi80B4BxECfPU4bSMEB142FwK+z6/
orlkTzit+hr/ifqcECt6sV9hEv+PbH+/h7OIvd3n4uxy7JCJSr4OzQndxAv0j8h7l54SkhM8dsyP
67kKxquFLlKf54eXb126G3lAbTiRVrWOaJcxou7FoH6h6/guibnsDJINUwunVWzr73Mzgwfe7vTl
uFNuBiegA8g28HpLqkJvvOzQrdzy05T4SfW5a+HTokn41y5Y1ZTcxvZeuOvKLyTUH5ZyO+ya4Qoy
Wc0jXROAaBQ98tbDlr9lL8bGPFVCJfhYxRM+oXuC0O0xWxq/PKu6NWZKdB7Sz28Ap2WjxOZK35qU
xQ4gZTG5Csm9gy36H1tsOGfcb2kpg8Fm+RWrFoGidwsm+97z4W+VO6vCt5p2bCmojK7U2I3S2ZBH
yIszsrYpjNppWDo/TcyEqg9g8AXYnoQtuJx5PUOceMIlOcskJENhJ15FacWqRAkpAWch/nGJdDyG
uPzU2oSN/UsTJU/132XrrUfSZG6dTtxJoLOK8L4vo3euTMOvh3s1bEsWweCWuYgDXBfgRGyoT5MD
k7hkk7VxJxkV/6KboqGo1XIjQ0Av1ye8vxkL0FJSsE4ztGiC9Mi+vt49YrJNpwVCgl1TvxFhESuB
p/EOpbIVWom9FkcIp5DIcLdj/jK53b0PO6j7CkKZdfht19e7/wDM2COC7NIo4NO4XKoMD0+eRnLu
IGAYodS39D1h25GjJ56w3mHeDcxCgqEcnQsWqKQFk77g3fkdcvuHTZCnlQPGlDmJftXxUhze5nu3
16SiZRVY21qY804eNrHC/buj9s858P732gBn2GMGlkNI11FFLHl56YLHK7V8B8/ZL6MgVTBVx1cI
Vry8c6YK/u2kaN7A0DPRSLbrJnHvKZXCWBc+w8K5VLV6fhrCTWO4eqpoVgGOR79gPo3Qow8EXdQD
BqnnHGNeCsqA9h4yNNfsLMrxJObaSnX4SuGZ0G0/vg93ENC+vPWbnpfMwkF1sofuxk5TByIxlniQ
9tkDys2HdBO6JSGnRTVUA4i6fYEICz+gJQ4pWbzmQMw3so4G0+FzYpfnwO93jIHsmmQEpSdy5bcj
b7JPaiTUXFBCKZDq08MXrQC1G68kHUkT37EYtfr4ZLUpuL/kjItuImjDfWg/TdaDKJ+Mun8MkCSK
CgQW7dEV1gcny3LiI5gkiZ9yaNTYA3GnTeYGHWcaKSTfwgvOJIJmSy0hsHNSrOFY0PnXYLRiLEZo
TSwWJkBNveVRdJVvPnbKnAPo6m7PBUrWixLYNX0UelFDKR7Zn+iGkIMwP6UjsD0tCZf3rWecTySL
J1VRAUpwjHyFVI3f+67zm1BAqY69tfx3xCj6teWqG7gmrsI4mKPbMnNGnuQZxqkL6jm4EIxn0xSL
gCVAjT6AFeC/C5EpPXj3Ul4EdVPxKc7uIUd5AMZbIsaTRJSrqyc7FceHlU2ZpMEIftGAS+Sgfvhc
6v+Hd42px/MjoUteP9RKpfHr8Q3iWM86jn8ppzAA2KHRiDUE4UFfWMkcd+L03VLldSiG2IC25VpX
B/idCFBsqagPGfdsH0y13ONtwkGplsNBAACmr5+qQr2z3+oY0TQtytG6LTzslTrDxpmxNE+bwE63
5QZVwHqaHzTXmtVw0YVo+A4zNRyuAVimBfQhc9le9NvihtVGMwoKWOtDisaTA0YTJPZ7NEsgsjX3
pTjzCRDDq3J7rkEwa7eSGku888Hq8TummYzIHkl4MfAqyp9qN+4GkgzLLYwZeAaQpuuIhclh6kqH
ZXDwhtTk5fAXugW8XUGVaF42Z42QdOiXsz1hTZk2xax1xKU887NgdEqLJ9/ifSTGp5qSEO65hINI
l6Pxrs6i3See7dL87S1tbjY/LkMwPsflUrUR1Al7Dr33B7E38DY8TRXcU8YYeE3oyOq2O32YtU5u
FLtfddjcMfsDZmgt+7+CkgUQkfTqmR9RSmjt4OF6lUW2AVP5WI4LJpATe131KnB2dDIfcmMU2wSx
3PZyD/WgzBhYjFuF+L/ayzpK9X0LOD50xOPZphSaHI5wWBwFrah4f5Rn+aE0N/7op+AqgUlE/VqK
CHKnbVkv43M3pZATqpGQqRxHc+eUFgb9L9EaBGWTSMQjQkm8YrsqMutiMPGJYJaVjq/1OBLEmNAd
kTaWHmrgWLjfZmCTPoq10a7JXSmQEuLnHbYCqwjTl63Zc/wS38bvEDSsZI91W6Uq16bkZNUZsNVl
SvZPun9NNFm7VfnVcnBtv13QrUSRdIJk2mkO7CZNmKzcSH/ZG1tvizecHcqLdbQMagEF7r/FyBwi
4ugk5zmYx5aTahrnfzjHdc36s0zgVlTiuKc08LYGIXryjzOFzL+sFDdRsqydAuAWcppP43azqaOs
EUiJYp0zTUEmu3Ymwol1qpYIciJZBriqwpuoR1MlmH+W7DQeXNhbizm0xnM0uqvyFu086yuHkV4e
wac4b1IqBS7AI8iU769amntF6A+SzijQgw7e6Ln7Kb81FR6H1M5jIiPcfa/CfqQV/1YT5oqMiHBR
7QN/zb359eBukTqsFVFzbz3sdGYjDDrUZstm/jqkdAgvo/wn4qv6Ij+Y/cpAA1REPbJTyiFjsiem
JhVe154e/kQX+DKEZ5gRPPuQgZljZakIRuZvMiYbby1HgDEsOysadMTpLEONBRcNbnB+POWrtiRD
Keyym7lbdZeIGELf6SrLnm+lk/Pb+PywUt75heFbap1CO8n6mlc3769WrWbTzMkj+dlfhgYMwXQI
TNQkyzCzhRXTQ/msTn0K00qY8E6YvcBprXr45OrXWJHxy5ei8pYU7AdP7GzpHrYY2XjaCzsIdUKx
INI3n2pnrBCidIYKsYw6FwTj+pEQHIvU34w3LBuu4P6tvG8GLO+IWDCWAf1mS7N83s7/2Kdklk7T
M5Eke8eDNKbljJBo7YlQPTrHlxSCh0qwYyosUMDsdXm+rx981bqpopRgOAcQ/A+rmlL8MOfiHn5I
Hgrlh4NPCl78F0NSwk3W3VoOC4IVMW67i60VmLJj/IPvOCMtsyyXzRiGfkz+owVjzGaKU+B14+rW
310tvabz77HN/7cNuCqmNUlrqyNF8pznh2LKqvZLaXzR7iqhNaS92Gl6NMhhwj/TIKMZzydo7W1N
PX6YsZXCVGNa9VmY0FbizMZ1kXmiAR68buOoz3h68/V/qn5WMSw4fI/AmcSbwLMxF7nBSnSxD5cA
pZy89CZlecaWsAeTW/Jc0kVKDDwudqvaeY/Cwvx+dtByC49mhZNWBYFAQWsTZ3XWuOMCNlUagMtm
I1tSs3g0/Dq9qc6np7gOz83UIk4XV8I9Uttn1U17EawZ0jKG2hePaALSgHjSXN3NuTThTOsj7HkL
Vkt5JECLZCn/eWtQzc8x2mYKpWqgT9Vw4a4NnPK0o1YZXPpr5nUrxiCXbbksAUBWDtI++GmXCrOY
K7mu1P1HDDvM1CNMUAoAvE4QNqwCPc0nfNVxKYkvZgSocsJ1JeeBKKw3HlnWobLkOX2yfhbw8s+j
3rQfQTbAXVISWSJLrln8hKaKDnMkQXvUY4zmtEHB6w65o+dopDN/Rqi1LFrtXU10BpL0vaX0LUKC
WqQsVUPpjCXM3ZJKGQ95zuJHkr8vDQFXu1gT5BCgMzDXWnsuOyHRpAMHDjc9YOaKpyTGTyoiKdeI
gN262tayzMUpMKrszCavFfPzFU6cDh+7WwLebdCEKbucQPJwDVs06xz8uw4xLp3Lt01PYD8YCyFG
StKZeXKTUIhiCymAdHh0Qcx4/S8HqIz+j5iDQ4BBLczZgCIsZgcKjgCyFaEcvFr3/1fENd6pBg0s
yg4zzfue/1RkP+PSwY13CmyfhWen2KCGsQvdB5lj0OJfQEw+JddGzUTUQ4FAolB9gIndOgzs4Kq9
fy68HZT2pDbJ0VyOmWJYET/QyS9OR9jH0TLVnbddkjlHu2llCIcoIKBGbq+232CipQdzgLel8mWD
5uMP5R9F0FF20/PkTSCzZnzoWPJcGBI7zEPssmyNsQrROVjAgannt3lcejfYi1aeUfc6FhNLIX7z
/qVtsWFnaY88MyadV2hOcjPUWTIEHEJLrejtAFrJ7mE1w2sjeYR14J1Xk5ngGq7yrvD1QMIcRwiL
Qj+mF0GqGBxdKN/NE8sogB0DUCRXyIkG7ULc4mXCL75ogrPsbuy79tfcwpqoJMMwmRAY3gxxTCIW
kbQj0bxzkAAI+Rth5qw8ZcQkYuR4uprKgKtP8mg1rJyHxFNT1Xjj9BjHYORVgHvxqT62cRrryPrj
N/ikhVGS1OIcx4/UDJKQiJbz4d5gDiGqqacaY70xYst1VnAcSWBYX2mz7KtGbSBlwK63kGS/r7Z3
mG+LnduCno9ElMXR1GuHVMWQFBaMOnVWemKM1EfQ84dw0ODlJe83v6R7J0hayDb02aGOa0nRWqIw
Mbmcj1uZZrmcqBbsL99BGE2qlXBlwPUGytW+dlGm50tk4GwEdmQSv0nrkWyfRUmDybgcKU8pV6UO
H4aqNLePu0FuRW4x9nBlFHizaUGNCehroJ1zXLSBTkINs/JtQlGpAfGnloIKe1vRqdIsdzKLb6S0
UI8MYNqhm9t8MTMqiCBPvYoVZ0LLDhmtLQsfInWpl7YfXbVJNZWiL2TqSZ+YuQek0fUBliL+KjMb
zhAWWxYV2wL2aiJLe5zZHQt0MtMg5sgD56BVPbYLxDq3o5MSv6Z0PkDvgVH0QGRZ/vP+wjDJdnP3
QTku/y/yWVUdkIrZkAiHn4L9UMVsL5Yf5IJVSGqs0lv/un7FJHKcGb/RVRS6gTM3zVRm+YIBAJgM
XQHl+k5Z3lMAuE8zyAvJs+sSWMi3YaXJ08sTU/ge+DepF3pNri0LKe76IqqBSf95k6f3uabJDB1A
6fCzQwbSPVq7uHQH+YidQ/AOrzTyDxASoQjp7cT0FqClw5nDN+DTM3TdQ4Dt0oqqxr8/9dvVcf/1
EUmXvPP63Hwnscr/7qRePGsNhIvJp5nu3Mos0/t/kcjHDbMmJZ71nGaSZxEtIsMauZerdIFn4cdy
oUBr7fb04tN9jhomocKYvF+iOPoWU+E3d6lY9xs0980V+3f81e52k3JVFZFfvb2Sgb1gWDo2PVuf
QH50/0tBENHU5sqgCDQwVGlv8CGetnj8LDCb+aCiTEumDB20QiG10zqvbfmVmistbPls6/AI6/Jp
6SedpQd/wQFxOdTWazrO8fKptvLYDT/E4UlGnIwpfMMCKO/R34ebPPknG6e5nDlHQrmDObF0rzAg
Z0fl7laSPRv8PFmAlCZRCsGHULiAUFhM4S+1mdwISaeqpM5qVkKhjfRNXh3TvitIfdT1HrK6s8JZ
xY3MHPakjG5+ft6yue06Fnm8BTPSkI1paNKkx8bj7Mr1VGtpJeudZMh18r626quwZxfpRrf2XryZ
isJac28TyqYKupcnjPsnq+870eHjTUcftC2MpRh6dBJDAhI4CRVxThnEwzCKsvYGdhsnM7YiwSWm
NkpkHlplc5Nrrwj4sfTRW57SLuiXqiSWcckCrLNXKUIIECkFdNcdRT+tzcbgZpFwMNeYGzRE8zpS
EvhLkVdLCwn55xyHFltjtkUJdccJdeSfP0ZGa5hI5sP37OIkHesIYgYZkZXhfJi7sW/5zHdDbG6p
ICfIxmTtg0EMlqPzskiOfx5AHiPvYpEHdlsnNbLAlqBBs/LJzkOavVhEjBTQL5+tMkehk+FYLcpR
fHh4+iekYOJrC654oHvuwuxleQFJhXjEZCFakiFWXpXT2NvU1qLNoXu4+lN68eRfaknfr84gr0Ft
+/8kEYl40S95XqvPBThP8a9QXJNEU9sFMnh7v7PX8un1Gg4/f3TVpJD/XCOzj0Vf+gMdyDAvyXus
93lDjGt3pFNs79pRToRWb7EziDbxjw7UBSD2UrCteUmC7GhEPB+sh54Tn0MAANMwXLUokxQxgFWO
RHBI3fwOQ9rdx6BfYRWDsBqSSWR9a/5LOJiubmsoI4C8F4ptuLDEgOEuv9X64ICLwwv9TQPHCS3q
VYIHgYepzJx57IDAdIs2HXHwk+v5a/0wkl0GxAvv2PWcqsFB/8stzB23xAWtC5qljkSBmP87+reH
pPsUDy96xYiKcJDXlSC8Gl4tqcMxtiNRo+RqeAuN1Qlsgr/dSQRmAzZiL9Ch0O5yjhZ0uboXEK6U
hUfh1LtOPVb53bnWz8M7N3X397U1ZHAv/XI0nn32YA9tcYefB4ajqSGuwVVonE0ylweiXEapSAIb
hbid03mJIEjgsvMrKzQ+JpJShSBDhyLluNZkf8HxaJU4BrszGXOQY9VUlgQvQy+RSW18ttzhitnw
kAL1xeLuOWXq36UAE9kfrw3TmM0ACn7qUgzZaFqNsRMALjz2nISEJlhDHo8MwSybnh0TlpZaTkSd
L9f9WouMxClpRT/dFPo34qJuaaUlpEMssX8QSTX0BVQDXoAbElQAXWs5b4X0QRZEEnWV2Atwibra
wYuvX976hVOKLqZVzwwHcIgn8AIdvOr6FYA4qNCMlICjFDbX/6igfyPi1FwL2BmMyKp87qnGNOoI
ijvkeNXxUO8nvkaliFZR0nKR8C1RW7Ug6WGg7ZeweXZBh+p6CQ7fxLRpG8Acuksbb6yXrQFyHhq2
m4sGpTIgnRgV52nokwRJvGHmn7KfhBaPpTLHhCLCFBlPcTy2Xw7isnYY8bUDs6SPYnmIc///qIMS
6pzJFFvOWp1u3x44OCLYs/LZxYcRBLaxo8b4W9UJMs9IVPSQJhIY7oVG/RN5uFRomTbBhHUpYzcM
NrTB/PWr9HQG8fGIqRuauYeHZ7z9rHAKDP1B25qSbUzmYu/cLIi5WXEji+bhtiid29HVFqPq5GKm
5p1/Jj1FHksSiHSkmkU6c7C78S2PDZSnTvDt2rLv5E5YoGPpxVxi/N6NqeETBnmjKd85Yw0zIc+O
1faFDpfxo+KPrE6gmWrMgiIV2B30BObqk4IbPyp+gvJanoguSBpmBxPDXGwQ/FI09AiEjCA3H3GY
qxdi/eEIdJpJ2JUsKJ9zeusC0qVFRSdhW+GZ0fFYTvnrvAthCPepRUKwtMFs2z2wJ9dGrIPsC/+q
9BpskrffSqXy6QtOsVpWbybXrol8haLBCTdDWxniUAMwp4GYiIjsPUfi5dTg6iDU0FJEq5CkXLnV
nzI6e93Z3DXuYGdLhB8vNai5DBPhZluOYHoz5LfGl8DMeKM3QdciTT8NJcxpPENKEugGCI5q9smg
Rw4uKCUBCWscN2gjAKABDZaPCylMPXEATh17NbN/ZIVTPA6HrcVgWEN+85G6Up09ZC0OTxNZ/KLk
r9+oFr/HOAqlEHHaHi1UbLA4CCvsRnhcdY/cz4mCJ1MLumTkQIXjN2H0igKCZET4bzQIUnhGEIbB
KaAcI1iu+PAUNF6lVQdkbtNc+0Dv4+Mj+elg7lSus3tfhRzndI6GIbZ8gMc6Ja+xdFNZOey3hfcv
ZKuzXlbf6ItK0+QLS+h61IYrnsnn9JgduulDI83QGUjMfL+1tGRAMCwvJ2Aps18k9HVq1l9vMlBL
FYmNHm+NQvB8wEuFsOn407n4o+4xN/IoEYgfXDfrUvno9pKGJWO4IDkXyuOTCA5ZwRBC1Rfe+CEd
3cNYPrDVDoIQQUxnWhE/88CEPoG7Uk0m1gCuU++/g6EjjqCBdmXoM8+ZXhm7PATA4cCXDKWGjkCt
xhhGZ5BInY01S5jnOfiD0U+5MCzqG5wOaaf0ns94Woo+8wY17VWzIbNbByuF1QfCbDg3bGMKIkGl
CCks9GNaYkXB9rYsdsnn/zZq2OvpuE3jcmvrqOB0/esxnb6M7xoV2Dl8Ds+ASJELT/8lYfg4r1mI
ZU+M/h/UEgwSTp5ZaKJSpza763w9XRggMr9hNowpcw+3hLDj9CN8u331CGXPcnK362BflJPght4k
baYKWRRFnJUN9ZBI0WoSlw2loVrHOXSTIGd26z1+iauPqPgLTiCuHw/YdH0fVoGHegLGpEsOKsut
SUW6MHhyq0a11XXurDGpN3kjICOlnFlwcd3ax49IrKCzzpNpafmN2pd+2aZUnMMa7LCAeveGo1B+
9Ds4T25djP5MP162+6TRE/i1BBAHFdj4vGJ4KnHz23a6ffVjOm924+gecy9JY7pen/kW76NRGb2c
9RZMlWH0prE9LNGyzhYf2prymO/ovdgoK+l1umxjuU0Uy6HCzS3FCp4KDhaVtPbhRRWWLpI2YIVy
Fr6hDAOu9azmS6fQBmZKlhohs7WXvRwnjtxJvzKWYjWbie/fPpt/n5Hp6iVphuEr06v7toJ9Rb2c
fvbENzjCnw2jq1d5+K658kEd88hv/hG6ImtnH9xmHnLCxApwCcNdHmY8kVQdaMj1TgBw/ORg/O79
GEcPSRP/PNdBgMUVgr56vuKtoE8YmdxznIfq9CymHD7xK5Svid/7b75Y9J4eV7dck7/kXswxBt2e
OmT4BRFylj35iF5O955J+uGgqCUurFvmOlhwVGaZw9wv1RtJEa5oGISZlH+LAM7GJW+qF9L/VyaT
gPSldNbrQiCH2mGaAl0Yi6sc+nTJxGIVPkR9cfD9E/4FUwTP2NVZ0eTnp6oRiNK/hsPpifd0VfPJ
0FYDg3z9P/1/KiQ0FutXhmz14t+YYWztJnv+Y3tcPtpIvbYqdZBBy8lgvDqZFe+eR/JqBYO36u+5
BceUmmgZlB9WBIVLLDdTmJONg42JZ6hAt3pfpx34pG9MDKwmbk21oOfIv+mFJGgPH89ERSprDrda
GXhW9C203zCCHieneORUikYnhQ9wTnWG4HzTNfH2J/CcCUpq5UKXRb90OzYpi1OiIwxIP1PVVSAL
qfwXUeUvSnCetDFWk9Hsco4WUU2ec3imlst8FFwIUkggn/j3ui5S5mARpu8owsuNQGsPSOaJ7y0d
JM5uzjicMqqWvOSR2Qv/RZMrytQ8b2xp3D7LSabt/4Vli1mr1USslchjLJF2+JMVCVuYKGC1MjJN
KFyGp7ua9S0/zlP8LkfCPxDe1zkw3a3FwJUTX9q80kDwysZalprwCHtnm/bEohFQ/nCT4Kg0jC0r
ZHyoQpO2m2clUncVW8Zq6kAvwUGU5qMM7A5cw1jApPB9dU2MBbOAdgl63yTB9QGwKRTFMHcYrZ0j
SwOTYT77SwXNeTfUNmlkD5+bH+77l6agHYqYoLdJQgmxyIgdOnLkLvHK5eb94Z724NClrtSrQK7X
VtcReHhn9L9CNwqfpEZAyDRrk6xAmcvzBPMepay5fDJ9PpK9puOgOsA8CFl8MYExXstGShgfTLZm
ZV2Zua96jTnXMY1wktvjsx3PcZEnaxOrwNuvEQtHRAS2XbEPt5tuSXsydIr03UYd5rywUKRIrspr
iwBKTyxl+NcKp0in6ACPToQB+jsRnUjtkovXK5LPnI9IR0h3ezmRLy1NEUoJrstZaqUWLA6DUz25
z3ynzRgmjikvEuW3pDt0L0p2Qt6WC4nefXkqGnv+KQOYP1+okgnFHICSGXSU/Lc0NebNLLEyE82Y
14X2Y+XWbzPMKjsQ9gQTgWBZsEatTU8KC1NV6aTirAzMJV7WiN5LuANsaYg1aCHA1Kd8ZaM33cEn
p6koaa6kFT0YFU0mEavD25HfQe15jWXSv+JcylfDQxBAaL5v1ClZa8u1J80ErCzEnud0567uxXGY
Bt8t58ZB8uFVLeHIJjcG/lWP0e3zIghqcje5b1NZLh1NCQrHgca5UJQk6wx5dBXOd7rgmOxyh+rg
hfdu9bYlDxwK9SDQKCbRcEHZ+vaTifT4Uu0JkgmY4JOwhMXnHHnjcvbVQ3XhKWMkfh1eoauZGQus
MOrVHWPgkKYZ36gqJQG1X+e2kxcn/IMO08tFhfp6B4+L8XpgA23TXd3ZtihX/4qPaxu1w9BYRcvE
ZC51i6dsr0yLv+6NFUU/2h/PWuxC7NmQw1/4vcHK/0UCz+NYkoGJnsr+1m0mppuwGhZFFEtiLXwR
vzrbrpXu3ifEEjYplZklIcinXjEulXYUM2wlMIyLEBXIY/H4e136lU2fdb2QS3AaOmcLFP094J4s
cvyJ/S+n4+rWzssyuySXp298E8IT87UgoaIzL322n+Jqfu+tadKhhziKRq9M4qwc3ZKIltWCvKmZ
gTYR3ZcydEDOQb2hvg/ejiazCp3QcvtT/yE2jV/yogXw4MrQiKWyoPRL+Hpv4br7KxcSncMjdDu4
0dr6i3VUpZIj2pz2qvpoGln9RCG6riSemI3/lhBSEAv8jOLnNYUEYEyp5FEI4Z+8SavbHCwX1pNB
6W+zKqjmvyD3V1g9JslQkcSsnKbgDYL1/nFjN+ySvrVVcS6+L32lDjefQAP89mNwHuLdzFQq9to9
i6WHJfP6nAKh4AxlkonqObQ+u4XsJanU8HEJkVCsjOK74I2MAuyAN5wfN9/Nz4OweOleBKLBTvrR
YIVAzylJqP8w3t/bmOuQ1up58P/9QvIvXuSCEmMjfiM8cjLrKzLfmDqK7CDunhw2Bg6FFAQqbvjm
T/iV9Q8iSs2jpfBwFIqtUZsgw/qcbcp2JHqqPcVJnih238O9uJU9oZU1xD6cGY+AYVkpelik8rPJ
nwMrsdVmwsdumKqm59a0fO0rCxYnj654cTCptCBPRb4x6B8kbM3yl1vPcQZsOMTdKxYFl0qQkFwh
sHNcrFEmcBJiEL5UvGCFO1ezlMnYoPZRXkZSn8UWNe289WBaJtRhz+VSj3EDpAJYAXLt64RDaIMZ
5aUep3AdtVKGoSO5Vlb/S4dnfIiUtOOZznJUgD3x9EA/eQ99b66FrWOQ3rP51pswdARpDRjXjaLy
eKe523PwBmZsS3jEccLsrjbg3cNkdqsRGwepV5Fd09qvU12nByqw+PFsM1pFSwNfHzO1J6fTHV6Q
b01NuOkgfbXKh9NDuwQyQK68+GQ8aMlrOlBOkyNGRST3pkJF0o/2AmIfVNFcHBhQ9VEQ3P3WkF6Z
L/vNvQNS2Vxmq4e3lwDdgkSH6Ai2EZg+Ovd0Dgdvjp+9bwtVgDcJy49h98ergyYemXxRkHDXgX9O
rt2EQ9DuDKDSTBoerzCRZoGRGcYc9cM6FeQl9h8liRDHmlAMSnvCiu0gZ2pof30FX3D5KOK/Ih20
OlzMijbFyumW1EgwmvW7FSHzuRBXm476RgJlJW+FCk4kv8hxeIecrL0UTDz/C0IqaKhQeKGZkQ6/
kR0ou19p/lQme2veVWcnFjF/X698N9f8Uk3vx+lK8Uv5b3deFcbNrFrf8MKvrOAzR6mTD3ntu1ls
trhW6CYhqUqdhvm1ps+h88sPFnhupcVRbZBiV/xAgVOR3+g2kSe8FicmS7ksy0CAJNfmx1uNOHD+
OzsmNny40umUa85FZslbsp/qyT/PEslo1F0n+c1cSBqMms4dC3gVgkD8rT4GC9haYkWjw+7+yp40
pRIA+2O0EnF8YOunM1suDVhTFfYpNOWk3mYKqhGnIL6ssssorbcos07Bxgoh6XFMQ6iPsfsmaQVX
U/4bFVRuzTGOgxjWTNs1ELtx7cfLR/93mzCz7tpl9bXi5jIV8gd0leElLuL8pkpPWov/112avvxZ
OhvRCzA+ejcNigWveR3D6uY/ZGLvWM1mkN5ZhZxKVzE5K1ENE75DrrljQoFq4ozhFo6jnCGogZr/
FnnxVMyA1f3sBm1HK6HC/zXp9RMBlK4iYPuNaRcJYUYmgLw0aElm+tz072VhbAFTl2JTKRRHafc3
SnEGGIpM9CbfRejaQV4F3SWLauYkFZNYIcSB+61z2PNrezNxp5lpB+G6qqV6q3InOdnwiuzQY8bp
PeXVgj5iEtOajIfl1RV9DSjyRXhkgnuHNPFVOKM/BBaLoRWqwK9XujSnb0zKS1nObXJtF7ipJiwt
BWvpLfi0BZik2CaS126QsCaBoDoLsVpXt5WaJyFlTwMWzACUTD7RjA6L/tQio+j+GSjDlzT1BTKb
W6KuelNAX+7wjJXVAfjB8k9YE7YdCd7YPMPSVvErDSl1otLfp543O/4HRcx0nFrtQIGeXR9Ae1l4
gROo/1EvVsNLUNxwXwfdDSNkE8vzaU+9o88JMLXFb02AoIpNgGreJ4nnFFAM6hP2kgUn/WB2CUa1
FnsjS0qFsKBY0J3ErrpRS81SgXBkd5jSbFrmaS0LwS+P62HTAdYb+9ctad0Ef7IbVCPq+Ji8YPmv
g4ZQtXU+yIrc0LebS0tMro7FjE5CJcZjHwIqoo7mHiZXZw80LdVojz06lrrjwlC+4osT3C4aE695
QuoTp1oeobQTos5akFWXy/nR3WHzWATcZFTxI7uAgGnev2YAI8abw7w9fa9/+jOTnbBuBkHa0uhH
j3uoMbnVJGKo/VQUkaXswxvbuqaPu+LA5arZ0iQjNGpHkIqp9pg2UBuxhoky8h3ijT2eZR/zmflV
mnbFQKSAPwyEqdKbyN6zkAUYzz7XfOUr9VdCdbvU6+gEs7dNVZvlRtJ/WkTSoCPvUXGJMnerrCnU
Fr89gMwxv0C5+oDYCm47Tzfr5wKHhYjsmO25gteLiqn0XhVbm0zwM+ypSIr+SC5Sr9nRcCDh63Sh
9WKZsKq5cwzOLjvncbEqFFGiR4fS0qrRQfl0C9bybXsAengXhY/ySHcFIeyJuygCgvosB7QyEUCf
eyVSLpjVzKKz5C35EWihXiWkp83wDC7pw+cjMJEw2tO0wGWyS8SWsMpAIKE3kI021/fp1H30JA/U
Fbrc+k/yw5OVlDOBs/VjyFmVDAnkRVZWbbqGw4g4gLxdWKSlq8t4bUHsamXzz4xuJY48np5fS35U
a1+NpSke50bqEVEOeB08Bjw1yQOLRjcfN4YlFd80hyDsVvbUqI8y8KRBgODhYS63x6UJOJB7Vz7m
rctqAKT/pEAWYl2ZGm4wMqEp3Qur/eVidqSNKcf+1Lik8SVgjQIvWkOIZWj5bjD5spKrJlT8TqZz
1PRw765gOJM2LbMCDU7uH9dJB9lgVhmYM3a65k5/n7M/7vGPN93j19W/1EXiZUKM8O4ky3oh1KjH
aiW/hpp37Lqj4suHlMnR1i0p9aE/WfQLgpW98LIrL7deO3yiT8XKQn1+aX3+ewfYBdVwhfR+yme9
NO6ItWS8KLjTbXyDHrWNFI5/HhvimvD0t+2Wymp1e91y566Uvh1t83iDzqrbwIfwOAjpFmtjPbLy
4Z1qGXz3FQjHinSA5Y9Qlm4EijN21pm1a02eOodWD89X/ERygLJ4oDxgWOpAki95LfY+H3QQ15Fy
ne5sSMTavTWFgjmYNULjcfKO/j6HYOtXMtRxOPnQB5eaoA/Gtl0Nro+h5Pue0VYLl1EVbCEqK2Nl
6grtpg/O/1cni1w8bn2nTEleXk66lgLiPIaagntmbvGPcvpff04JLi1p+rmNAaJzj1NxsqeqDUd6
j0RY4kSHXgVrM5X0/PFkkmzmdy1UzSHZyXjA3b4KYvJc5BNJ0viY6to8INOpFYua16yKNhw4D8Qm
pr0gK3O10Dr3Fc6AMzRK4PDnQ7IwdXS6lIYmfT9zsqPhgoZOs3QYKVMNmgsFYxPDWmCKC1jVa3FG
nIMI7LTB+USufiPWnV36KkcKewARXJo8SkfQoxKkOd4W3mIXkq/Co82cEprsw5zOrdVFuXLfuJ0Y
XRfQ9X+beddNHP4ukBgn8fQ1dg2u1JeAlImGNsU74i2ig5refsbRXkjOdMoUbJw5ya5EkkzGxocU
VQpjl5zRaIY2uv7bIdgHwR0vYcrYhTaBU0mUnvoTIMDhUb3eJ5clri2pnE80qVFX+i+yGnsP/E4i
FnorYyE2dqESo1pd6so5d0wu/PSyJp+RA/myFfIPBG14IqdkV5zzn0bd2jx7ZbzLA9H8D/ujkwWw
xFjUV/agkK+03ODEhO43WvmnxjB8w9OU50dxbCr9aqeqwWpHy8g6IZLdS6FJqD/FSpiwjN/VnhfT
NfsGrf0ZH90mG969/3OkZTmzEvA+9Yv23JiN3GzN5M4rieCRUmMb1Z2kq9caDHbXd+GeZi5LpWyV
ABXKZXGBESrgNwLTs5pSMasmyRlIhcI6uh9/8epzk8o/45o/RVfX/BezCJZLgyiXGaAaMm2qH5yN
YQFvrzAb06f6VQaKYLXUIrAzjWfUno7DHja0znmuKybp3IM4WTYbwRD0ushjjSd76APVCBaTPphy
bXWTdDnD6666qXgmVMQyDDYJ6jCsPB+Ct8YLXN1SE+yaXOaYSHr4zwQkhX51qnKcbZlpi+KIbS10
zwqQXnGhuLW9I2ApRpDUg4LJ1S7UDsVSpgbzst2QTa2UBMQSbgClpFiGMuOXWhg1aDdr3j+gp9eW
RDcdsMIp8xfi1kY0JxLnj1ExbBnhUWAZUOUYy0CLhgZWiTSDrynOuc/MmxFXmpwVsIf2mOkX/qJ4
ZinHo+OzVlIK5rV8ZYDYX55ZgIF9fE3PJgzLfy4wa6V7vkbQQuVXQy1GkCpiAhHAu6mT83UtA1JN
JIf6gv0AuKskEh0E9TesG2RFz4NYB3oAhvWTuviBmP2zCAjXheYm/KkjNSozW3GFwdcThV2F0dzR
iA322yg6PfpDu1Hrh0PwrAgwvFfmMu6wPUaYqaJSDFF6KdhXYWYJQIFl/jfLK/xtXLGdadrfTEPi
DTWl1cPEpomMvcmthX6AAftYxudosDgsGkGkqiGVtiZ7LVQnX8TIezbhIC/K0Wh3aDMI7wtuQdpg
JhlTU6Bu1jfl736h9IMzKDk9rjJQlp3zUp0T14DTzIOmiuOQhNmObAYxP4aL2de07zM5GhiD6YKo
lVeBv3rT41VLeI/9DulwrrZ14xd8kEAY+Mo0KoovhZz875yUXUxKhmeiV+dEjOiZIVaqvRlwXTEW
TJYZ+jfBDHKLxLzUmQop4q2JPSu+E+NimC4fOmlgW++wZrf26uTzrTN/4SSblNY7oeM0KERUROma
6ZR26+9NpWMizl1PGGze7elsOeqt/3XHD6OkL6QRW+ea1RTIjjHABNhfI27We1rqJ0t15H/3EVFp
Wzb3gKBAnFTF9Tg/0rd7KDbP3Wgwk2324QksnVT2aJD6401nuKNzINI2VihqjOYopE6jya7fK6dS
qBsQ+RM1rsCggLjYhZW1qzPTs/tuB17jVh9b+XGfdP/VkdcbEQdgDq9trNB3FBWnihYKzQYFiPHU
Oct8eEX8mjU+yMLAsnjNbkGScHJ6U/rzHMY5vwjWajYQwXFd5bNmMRsm57s1EXSXU5DmMgszKiv3
w/VsgJZqURbtrfzKau9sDvNDG38QjI9abnTWnaw+4cbunXwAPRKr+kWUmEV04VooA2yuIRh78nFR
8dcSRtZYD25ktybu7MmSOvsgJ066q6ZBenPjjUNkqRvBPK/UKt6WZNc4lMP9dVxo2kEN4MHG2wsW
SFf/aiOai75k+uyzAVifuOYH4y6g5JmJia2Y7l9YffgYrQiG5KU788FBhnZmWwmIde9wwxEjoT1/
LjpCdEQhfKYoiC8bar0f+X3e1Ti1iDBCM9EFN+wcvpJTguKfbxhE3SeiU/+5s4PQu8jFbGoLr+1P
usJ9Qhl8q27x4szMbjTc36hq94mwqY7AiY1Ny4u6S+4UQJebMg+7GxN8DP/QemxPI69W1edv6Kvy
DWuWnGpa1WmsJ1TLEXRxUyJAcJM2LeloRbg4Qv9/oaW3ajTGQ7qCkxlRFbH5QFK9TtVClJxbJvcf
3eyP/0popjxg2I36bifwCJMPCYrYg8RRNQA/0liVMGWHs4QPp2KsKG80BTKyhW8rwyNSBwD8wBfl
RPR52PcQQXot0N7OhOFiyYvinKGZhmHsAaHkSl0qxQnqY/OZtWXGklZ0hIQqiu8FQEoXVgyVerno
zu0AiidEWOD3je6um+bu5rsJVQj1zQp5Jel4G0pRKgw82ZPWAhaMRNf8XsarpfyIiNZO0U1nEDJx
m6A7TkYr8nBNBgJWSwDKXFij58nIRAX5GtaFYifEDJ7ppsZHU+ivIQiXH1ppJ6Ou8J9VDGHH/QZG
jZoNefn6VfoICJVO/tJuR7om5LxkUwVBxoTKMO8uHOsSCXK7NRyHkOa1F2OjMtA3U+xX9z6Htfor
9yYHLTfqd7yhIIZkTQmLc0IzbvayanSTuzuZOKSyoV+kVZFUZsvnQBYRR1+kltnLkrh4gnzoGChw
LcWWVxji9U+5TtlKKeQUL3N2U4eCeB4vsKVG0Y8Y5wHtzdgL6IHk9cbAvyKx0yqWcXBUP5952qSB
aGYhptS9Mze2NbdjtizWYoGmEAWcbE6R5atRV2FGkvxEElRBXovh96u5e8CnS9cwxdIJ/qRtnY+C
zY2EqJRfCl6wz3Raxu851wAHfCT7hsq0/TO0Tvj9GfIYfqKobBLTxPfk9S0+YvZ484xj8kLd5tka
PYDZV4eIOrFdbsObU4sAckZr+zo2u36RqirTPMTeTOIhaRQCjq2MmpEz+kEx6V13jcqttrUMMbg9
HxAE/clWIrmU98JTGDqZ+2z1zrUk//7AnRpbTMkmLe7PSXdHfosCzJk5qnR1DutndwTd0ushI9FM
A7RqhsVB/IxzvmiFiuqDIbt1GSL34BjorMm9M48ZLE049IF/ctioAaVSGAiqipInt54xm2NjkJIi
mzLcNKH5FUcKLG+W8Bq86Qo628WVdFt3IebXUX2a0De5gVUDm2NItazL15dmPKXLYLVwrV8B7y8Z
l5WUYuPURk8hs4JKUBD7lhr36+/zc2n41PtkSm3xJ0cCN9vn57RXUAWetxyqR3rn1emPAE0VAMbV
n7jX/eWU2RR4cWeaVDYjOOlrrWYwUsaIeSYFfC91UUYXmYzCw/PdTXn98N58elGCBn31VYMj80oV
s+NK1YDfxV2nZsBm+cfvX2XPzJ5YWA2vuDBq32Y8NF1rYg2wQWF0DnOBMryfZRmW1Vqq+YdQ9WWF
XPc3wBiiR9rnec6IxiVlb4kOGcwakUCsF9X/D1iXodPi/kxADtxiIp2CS8f0LYvInd3kWNLdTQrx
AycvTGzxBhWZVVDZn4ru5Y2x3G80tb/M3/UGMkGDGr5Q3iFciTm0KdSyWjNSuABJgOJjS6VNAacX
frQLEZSz3Fi0qK3UisSvLAIUg9725Pvlg8NU2/ijtQQA5S2cAqGNdIz6ckzHIhohQAbdKiuxsjoD
3hWHGfwY3uAOKsJRLx9gJ68DcNOJDN4fX8MfcCF7KP44pPOlPxv0aRRDNvPiIMHNsbIeXS2O9GyJ
fTfiXgnP40bw1gxiQGr9yBZ3jNmK9/Tqesda7AzqBnHyoyJ1Or+CByjHZhvS2i6azHGJDvyjmwGk
z6WOcH+tpYeM2W5m9yhhFdZ3/z/WS0S8evEnaaMk/V+AowZHBsN6J+0ZOaPM5zcs3cXj/tv4o2zp
mfIPc0OgAOaalxPK6k+Ua28LZeLGKoaEX8NxXL81zvc1yrHHvxNRRP20bNzci6TtAmiDchSqG8Jn
U+3AsVHYLRO9wm8pdFjohpFCc6/YRS1zSXnnvum8Zwiac5H+priSm771Fb42oElAUhFCJuR42LLu
Iy6o+IsoOvRHVfHhQhifnFU6w+1IE1Kyks1NAJRLeU4YVBHem4+BiU80Fx4Wbi23Cv014xBXDCh8
koq0Wpxmq3jLIn40CnYt3G9XWlZsen2+aE1GTdoviNReHMspCBv0OIasKm1qfxwV2rpF8hVuXEDc
jotNTOaz9eeDj1/PB2E4lM+MTH/hb4V4LRlCd9LOYnCS/ryB8Swirmkooh61Jj3nKlYwgQp6KBhO
78OlLGKtJRhEI9ZM1riwohxIjlj5IgKp1jXsRwZsJsCLbjeK2787xjsRa5LiO2X1yGfINby0EL7t
0YHawJQG0o1IUSK2isyP5G3g1OxsakCcUZvyPdJ8qhTb5+bhbE5ssy6gwoWQGgmVAqt7eI9L/+S3
eK5pDycdaMx5rtvVsEydqP0BLEw/QUr5mggCP/hEj6fH7i5wJ+0C6YDJlXBXuCFp2jfbpNpw61+C
7q736V3XaLdND5yozOIZlNYlduIbH1SOcbd1DD30A5c6uF9wFpnrbwBzN/1TnYR+NtcgzOk4efmd
va9Bb79PYkIKDv5WdkPk+7ZJLNapT8+SF52oKQCUjUQ0HfGkfNDJ4NYGlxxBXZ7AyizpLobCa1ET
sNtX53hpnidROs9m6nPoda81fvEBkw3UqK1dRMdfb61CQSOtb0VbmGCCWqwidbcAClR7nKPb4NNc
W3/EItNtncVsL8z6TIDjydubRMC7aapK0D4TL7ZEULv0P6DLLCtsjgKrJLoToH8tpCIKUarbZtg8
5zNqnZcANwybfCAJSPI9pXQEF7TLuPBD7V+f0Qlf7avl1O/zf/99EXIpyKLq+QfeTOB9pFHZH6Eh
j7bJdf9bBX4U9oUgOno32vKG1oIghVp31VIwV9mahandSQ9OL92XjcZi5HfeY9Ej8m45DKA/AkhY
484YSI8WebQsSlWFqYAKBX8UBpoc2IjunxJgLHVED5BzIOlp76+oTRhIuutcxCyMWWK+qMxNWj0f
qvpYKBjuys7KK8fChE12YX69k48Vt9qnNv2/NQuwzMtCBT3kE/Lp1Z2ZCrFAf3mIlWW0a6UKBrym
WhX48I1UdX192JrBCArGP2gwfQeEAVDUpuFjEXWFsd1CRfFC0+SThcLo3z41ghV6OFzvoA3oj0GA
pfAX69v9AetvGz6ORAIYxcnyKMSk3PcQyIYbjmw49gMXec2QhjzfNjEG9/bwtvNgqvL+IZLsh8fl
WpsI3srFoXLMZ5Q3CcxyIvoWh+6nbkKlRmTxFVqPX5sqHecYeym9YlQe/i7bPPMmlJpmXv4xXmXs
jHdI1l1FXdlmU4TqEn6uBmypL2oXkealV46LLBRqUUp/SQTrUtiBpeinuJoMK8/kjQ8/d6Sepneo
blPkJF927tiqoa/5Cr8lspFI3DktMasyrGKPjESpyZXcvHXSKsmdnOXGCHuIsCTbc+q5OMmK4scA
cfdk2apPKwXbpgVYspKQDR9CPB/eRNg/O5U/WEZAeJWg7Zg42+9AubnjdWwxBth26TF9zdNCrJDT
kM6x97shnPLwRlTqPpxfRD79tX0QVsVF9fWFHdA7uvdgcwoeBf0mAxOsqwK6WlNIrgKwhI0M6cpN
zAparaid2Z0qCcpelI79pt1CB/af46kClLcN2nwcoKEm225HLPNRbuZsLeGYZhkgQUlLFiRWA89m
IQXOO8/GmQnUZ+w/tRIwmWqpd7bjnzjQo2/xHcMscQl4+/34iRSinYty+/X/3A9qS4OPHQZjSSlU
X20cxZaF/MLigvNPEw4qEOcABa3KHLoV0BQEaDqIpm7b87CdFIZ0rb22ewGZGY39a/hNnnAvUwaM
7q1+nNTTbfOxdNYH9zLqOx0XS83Bp+jI7qhJ5ByBw16NJ3V0lFsKwGL4cl4qhpFcLCEXWHyTsifA
TKaqzqy66SFVG/RXfkRTMsJiOtUjRtqgJF47CKbr0Y6TspoI3djyOkW3uyXqJTEdGomfkz26PkbK
jtoqhDwovxJw8VIgeEDIVR9etxPorDVL1T8To0/QUsqi7YHvdgyYRSxzLRzrtXu7swHLZcC2crSW
z67Vgm67rP8LZonGy97jgBwmkgE4DDPLjym+IDOVdoPoetZYY1CbUXFx/S1sxicLJ3ldlQYFAoXK
qv/XSPPsKi6VMxmAV2pEp8bDfvLO98Pbey9feFTzquZ9qSAmfh7Cfk3kRMLf97YOInvClwM1IYGR
MawsC07vFKwBSX6ISXpOGkbT3YNJztoHhk+xMUEXpp4cu6qwHkf0hZaQ5tlDYZ/3d3Q86cjhXhgV
xtGqnUVc+IeOaO0tnck22O7LegVupjgcxxXV4p7Z3kKvjXqP4Al71DhWkEYvimiSwhLvld2Gu1Mx
JdKi2AYcf6aOOEbeCF9Obiq981bqOptZOs+8qrD7b/p6i7ZYKT4DmwOms+OMVBg3ecqAnQMZtTOe
xN1AWJAh+KlBBAaxv7JIfoXZIOgw3sUoz8bWrQ0tvDnT2td1pCanHFkX5GGbaiGhZITUOdHuFvQh
pUl1PBALwyoSAi5tC3gS+GyPTZx/Um7d3Ox4S3sGNcowwDeHU5cKoaifmW0GeiAT33G5u1soOPZj
FZdVAF2HJI8cSpzUOozsMqOf9fei1tPcHBWMmQ6lkoXOmWhr3nqphKKESw4r8I1uHj2TgNzX65g+
37cqWfYypM+uDyN6xkH7lnaTaIw+u29MVjh7dhv1DgUeV5/bjwxPMs8s1ZgaIDvjwv3PMnuzL51M
WwP9je0DJRJpcvK+LJHzo+/xUFgrabNZSSOywhydy61elYHgFgVSG8r/zd5QAhb9hyloDI93FxJ6
V04zgcz9G3qFIE/ZSkbtSPUIZXMDfqyk1WHhyRjaWtK0cjHU5hbdfSt1qwuWrsM9Ngf9p3JAyx7h
5Tkzgj+8spS/lY8fh4rvqtbWVW3rdlsyvN6ay5IE3wSA0NKG4q60G20Y4kPIpwz8J14xdWQW3AGM
McwQMjKViukN9eQ12BBCYOE2PAoeWFXhX7FUyeYN4HoFjKmjNh8dzptchy8UxAZWx3Jue8jV7E2b
AxIC7sY51TssosGofcdkQybwMGl9LDyOZvOflorpHiJpPpJRbujMP6riUzR6r8bMSS1V7nrw2Or1
X/sZOJgvRXjl4EJ4q/q2mK778hmSvBa7UHB0rxALFPOv+bg1qAFmLNsMng+SzuEvetBa//qJfxtR
MFi/oGK0UBVwf4u5AVA/CNegjH2IYu6t1asfgLgMs/meunO8HFZSVlqtasa7LFe/0/gXkRLxw9qV
9gTyut3EjtyMoOvjENFfR0IZcO2RhBAzQnNRil50R2sP/EFueL2JwokNwr59Myqk4O8k0dlb9qJW
9bpbQw6PWJ6B3wszB/ZigcLWNEJK7fECwky0k54NBa84NXk9r+AiNqet+ZUUay2d2Ar8P60O9Prb
TPAsrB5faQzKcpbus/p9KYmTCqYXoc4art3p7/k/6mcKQXZulILotYFKref6r2nwTt4nnfEAION5
W9qgpJVwI2zSiTTKxAsbElSoiInETcV/NX4GVoz3DYYu0HUFWKI8NVixeFsmjcpbUMal5bqGumxJ
4Uh3mxOGD+v5FH8vHIq9Bgg0ndh2SWjxJdA33ngrwWpvXUrLgvdKJAPwHWYQB0nUCUSQWYZDt3/H
9pfASW9+oOFyMekupbgo/Pbdoor6uCOMDVhUqq0xbdhbl7mHJXO3gQhezB4da8byEvl1gr0Wap6U
4NHQLrlurXBOhaCbfEqw03/DREhX4kVS2pTLikOariClMAfsxa/8iQCZcnuVFch6f4ky+LZvsgcv
Rqm9VrBBMew60uL1qldjByU/D0glA+6jpv5XMd+IODnQ1cfp66h+GaLsldshGSYJRZ5BYXLGyiTZ
lW0vli2WM+HstTMNJYm79wM29ztJt/SbZApXlDn4l1ZS0LMR/P4kZZTYHgwTvgYLSWvLX6tXjHi4
NaHDtob/uWjujE0lPwwH8VOVkkseX4YJ/mTyY57cGamo2cwispUgU1xh3IW6fyhzRNfueuZdn8q6
yDR+OfgpLcGh2pHtKAfSXq7cP+dmxtmKwN20RZ8K52awCaqS/ydfWTmKh++wRGuUbjeuH9u700XU
ZCRNZC1Sw7KsKILvjf9eEoooNrb6Qw5fdLUtNNGD8I7BU1w9u9xSkv5jRIJjVunK9a9cwB1M4orF
eNogpta4Jmu/+66QdKRnTqxRk3yBfSGYFVcsa5kyntFKhrGlyfyYK5+bvPLegBovcQj+/SheD5yP
FrkUkM6X5SAGVX2a8+fbBJyOuLWi0xyrxRsPbZNRxEGZdFil5xjppVYHPdstyJyCVGw3PyIPAJrP
o94DhKv/qak68mfp3DOaXUe/byg5GbH7iStRehRX+xE2RykdyMMhETsq2ZHiNhMlSHt033h4gSt6
l0dbM1BXdI9qfwaRAiAevO8cB8VD9afA5XuVmY3GD7Fcy9ijzQrQAoaNDKsICbdRnal7uaPijf7u
M8QhmV8fXyRn5sudL8G2RKEOMilVlXYsvpUWBggMA7i+Ho/bH+rc5aKxasBBr2QfFJB8wMk2FHdQ
opJt4Hqqn8k9o1P/6UUxAbpvofuiMSLnRQtQ/LJKEJ+jy1CJnIpiIWEnkSDknC0Imhqn4XUHuitj
0p8k6mgvqLl+RRfOzMiw7Pu4uP+FlAn4hcOfHN3Z+rdUTYNxJt6Z1yANPl01i8HIg7l0nqs/IbbU
DhXCD8YslZ6otTMr3l1I5vrmsUd9t9cPPAW7Uo/kUkv+hhDTxIsqR2xQTHbVhd7oeT7dGC9EEvXM
iWRM/2V51lMVVvG/K1wwh0Atj3tbLx42C7XPm1Kp09bBQ01ByDTTbCCOFZ2gWczekdBLzLHuCUrx
ITXR3JP8/SWNxzJKQ+Slo+mBuZBHZF6Z76bnQpv5L6Uba+r14OvbwWwTHZ9X/5j1Uyjp3KUISDa8
AMUeSFopzpLTBEyJ+R92x6fYFAGeVm0iW1iMREE+XcHh1h4yedSFpIalONf12iq2ui+ztWciwWsN
FysvZAo5/MM7gWky8VBU1c2Ds3aMKgeJjPiQYJIq1cwF3zF6q5nFyg5rnShp/CnOTzCQynt3J1RL
4p5TzKqU4Asz0IcRG+BEOWs1VblQ6EO5SZaItATsJ0enYtt5O884UTGhBh05MU7lOCeMQ0OvThhB
QDjLqlFpKhfPmCSI0xo3fGgN+XpeXm1cHihlSSUlg0ubr54OkXjcbqusFVTMGw55XSWftD+bjCfO
pIZ7PFqEJFi0ZElKPyeydEmsoOl7CmBskYuB3IoXHTwH92uD3+y2OdpLX+Oh/9UUjjoDzj+OLbgJ
PbkYeHwXCOWpf2gTJvwIHDz2jFdAU0PhFxcocUPrbTiGuimtMTE0k9bH+TKUaNWnMZHdSpRgweRD
gjRCUzX6MmaxpaaiLUd3PpVj7oNKlFlolXYV+E1J6f4/yqR+v2NIoanBFM/SLzOTFO6Lw8SRimyJ
QzgKYm4YUwnveDEREL/BBff5/uVycQkzi3FYaAOTRWSLwjZ/PlguMYfDsjGBBp69eovsqR3P53Ub
Krf7dNinTKLfAc+j7ma6QUCspgwaPh1Ny/HuhAthUj95YZui61FHx5An2BL8iEBcbJefOEq1hzjN
MTaHozc9/j1XyYJk21IeZnqfRi2XQ9q1/BQkWONI6VwE1e6/FYI6A5YGP4whN6sE9Nj0qk3/nLtD
sAgzKueeu+iF/zngSEUBY9rb4qFLd0tS5T0D9T3THG6uM5JrxyNuFvSphLjlYPZi4CV+9biRyCUQ
o4BGXw6f/g79S1Zr2gpyFr0cIyJQv1wCZRLr/3JyF4yPPgDfj9o6I53OL5DN4bfodrBtfs6Rkn3C
V2n3geOKdM974ivRGRXFQrm0stREDAxXohywYoINJkv8oSpCZwFqmdxXkPxAcGZNefFBrY2/9vYv
XQKxgDpeHvNNkbCMteNEwn8oHpeIXpjXq3zHHu7prUS1QAqzWwIPvlZqQaA5GUlpWobBSUsBf3AT
zh4u3HcWtWCcKsICqFkiN/B1Iawd5CKYuMcHeBaaMPJTP77ugFcvJNc9tEZ+E99WHpk7Qb0T1iwf
ZyZ1FTyQUUBEj9MQoHY7voNf9zvLlsEEvrviel2b7U/QesvYSLnnfJA8T2ks+oCuJ6eSX2PeAGB/
dn12A/tQXfWNSQmEcfvnKsLcEoAhnAoDWSS/1xTEoUztIuJudRCA7BWvD6WetxhNf6rcdz1ot48v
bd3b88tLcPULO5LNuwIdN5jX1mI5x7LMNJ+DsuXP3tqd+B1Kc6GFd0DsduPAR1oIewsFsDJ/6Rto
G9f6TMFBBGrLEHaRqWS/OMI3LAMNJj8rL3cqQVgPNJzKNwM9dvNuItoKYILRv2MH2eQkFzsXLlp4
X+Xh0TGah+0t2ezcq6K95Xb6Ymke0UXt92HIzxOxlfIbyX0S2+TIx6Y93DYQBTDIzfKnrTfCwstm
ur+6ERajGGU7dGw4WIHCZrcl+DNOIIWGaHXpHPBnCiFkZw8Q89c3Y+mgTnY14mNo/N214eL3fOC5
/zQknBf75lebynMU3FrzKFA/v7Xzs+PLe3helqiHZYQ8s5shl+rhm7u3y+NpwKAkvRrWi7nksb+U
Ljb48DhAijpsJijpljERAbcmIlOjn1w0fJQ5J84xf9Hbp5wGb8q2elK9nLX8D0lQHgAOHVCgKsvN
qJINOrHJHq8aepQmTBDdjwaXAILRFYFryHmxy4H4wOoT+8CQps4G66whHaQvpKWBxPYoxNUKcFlp
JyZN6T/cAj/ks56depTGkOVVfNdy2MHQlO5Xqh4nolZNcqzNODZEGkxPfjDgv6qXNxViKnaHOA5D
6g7pSnki2bgIFrAsf1TYMquMOOYgmgHbOdVZQNrA9fkKMMdqeR/NsQ2mm+SUJOhz3rr0tyIduS7q
NpaQcb69ZcAUgV7AXqXil/xYbJjiL8PXtO5r4/4xiJeYEQqc8cIj8L8mresokm29mMhysc/hm5mU
71VlXsla6M51jY9ccmBrOOb+JhHE1zjHit5Fj4ukNJHOOB6IgaNq6/pDi2jTBjkrTnty6kzC+m5E
HBINfxZzHbIeifHoe/W+WSQwgGqQEp/P7ukyb+r2WX54zQ8h6lufZ6h5wEoUrglHc2pKpQN2bRKn
VUi+B4r7/9af1Xye8B+JLZ02Qy4xD9jXRSS4j4hVU3nw+hzgiPGyTlU+7m3/wen4QKc/+CuN1oFD
grdp/W9+wSpge7owY+lTWABgMlHMRINYGa/WBoTUqnIoRtouYEk0i9EgfG8qWE9V5M0uy5yJBLVw
PwYXlvReKT2EiNve/vL9rzJhF6vcn/Zfp/8thiAMDyBoJ+E2IjgvcmTqAaXy8Iera7TipUy9K15z
LJfVP8wzfUmZqpEs2d2cHQDMZfvXGmRFlPsdRnKxPueePs4UH4byplrBAWUFe6Qq8GYjCnNhksZy
SjZI4P+jvja6BGtIKozqxXblSnsnVDF3m8gAEbfvRJkk1A5lfcYOMp6kdjUC3JrBQ3WlkHGUk9qx
3UOvycoe0pvqBnlFXwC7MuxxcJaR0G60l5TiRUOoquqf1GM4bpNgTrWFNZ8vKyxgaa/ioY0iCKak
Y+zNI81KdNFFy8FDQVAheR2DcRaIsvMeZa3TZmjOwiu3AF/AWofBk7YmBmb6w6HUt6NdpmEU5wxs
mOf/bb200fl4apj2BT+d6NGu8V+QaojgDLIBZyJFSZ1JaBFcupWEBk2OMqbB1OaXOYn2nOdhb8o1
pEAAW6ncaniFXy8IWjdxe2eGYlRdNCAkVZxl1efEoHviFLbQgAhBQToP5lKDgIymJ9Na9hV/kaaA
cqBXwdZHIqxj23S55x2hvpNzoyJnT8G3rZaumtbWOxRUNYclR6SU3y3FRiNEv+kxczYD8TdSS16H
pJA9YIwA2aOoHneFuwZG7L+1iwNdOIWYlap7K/FVYd+hCHMBEh1WsyRFI5NEfp5ibtnvB/Ko8kXq
8JWbIXuzHZa3qTF2l/1O4qXngRmWqfZBLqHBGxKdrpjeunlN4TBXYfIF8MRSmzvSssceI+nL+0fk
+X2wo7LjHhH41N7qDepiBIl8VoxksP9cSXbcnkt76hCGsjJOkHwUH6g3m89RjzrlQ0p773jUyn/t
ueU0EN0FVUUQrO9CfiNdYOyJP96euG1dOVnIyhRoF3qBkckDBI+l3ZQx367G/c5KTEDRvLgMAvfC
WpYW19qNzS8YzJBKxlJtlgHZRMQR6ALtLn3o0F6eGmZwAWZ+AtJGq60TrsInhgNx9qDElvstuCCZ
A7dL4M9oPu/93ac/71aJ7WUYhTjeYrhF073YwlgYhZ6q7K5fhcDjh/tRbsPEMQ/jjjXjqtWaSa1k
jDd/uCkb92UL7ee26VA5GY3putnsb7cx1ZOaxVFAEXHvela+WqCDinBcqtE6/TORBF4ByzofrCbE
8XjtTql0cqIlaxVKdoMweCJIh/NjLU+Ms9jCXSyYXKsjdMWilP/IJFlj0Y8zR1BrVqrpJdLSfMmr
9MpUO+8O9G9dTLv5TL20W4UiU/WPUUggBrho/UXbpGzqexyYPkaeyoxdzn7NL5x1XB0oKvVzjASt
2uHNxkg0Yy61/Oi2fTwI0CHsiLQyByE5e5+RzMpwfK9rUhPWU16l99UapYCbKMZs63vA9A5WHBoX
loaVDvwJjnwmGfldS0n0/w5oTbC1fVwX/O3J4Sxz705PekdgwvJepzYvNn+iKAV/JTTuxW46lUBr
IpIwJLzwnCRVFoWZju+IJy8CIYrKGC8B5lzl20fTXeqP5l5egs+LLa05hvBAP9SYQj8l5jLV+U60
LWtY6GrPRGLYDOZVHnppL1J4Jwk2HWQvDc9bA2wqAKrUDrKOswLrLG7+1JbPAps/AZL4EuOB6kDm
L7u7Nu4F/28vrZU4fYqjc1JeLn/H6Cr02lJ09m7K4ZgUm7izZRu5du/ZDyi7VGCj81mJHuPUXJ8J
r5Wez33c4L6NHF+yQlb6POycySSNCVBS3lnbMdNiy7yLs1bZbT0wrpOlyNIsNtOjdut2FgwomToZ
QAuLdAn5qHWbeO+8gc8UF+9rBgykUr7IF4E/4H1qKyTSZ84+z9NLUZn7KREc5vTsiqiiEPTzpdNu
MVemujgf5uuMnuUUqmLwIeaKq9eIKh5ztJRKpsD1RnFRidlwcemNvo7PdMENsXfqzgPYPaqKnh/z
w7a1UK3t6FAISI1uPCE63s1EDCmVH3mPPVoQEhDhE8ueMJ768watz4PIyUpM/bdvaGu/LBOrnd6j
jMsUnvJnEOSR4PS1UYFbi85QZwsTnBfahvSs8GEdntvQs+T/cA/mSO3tfXU3zywulOSzQRzMJP3E
bCYt7WnQwuD8RDxRZZsoU2HfYsXyOadCxDsAcEidVUcvRyf1h4HB7P/fkBdOx7Z1L7Oa1j27VQ7H
Og24pSeH3Rbb5kYeEyUOcrPqBgztnT5SJECFTkv8RYAp5sM6oPMNsKh3phieLQr1jviE8z+reySS
sTrHDOUzXQ4WApzRAQe4nx3KcjgLDGB85WrxWJDmvh83/tKjeI0fsK4iHLI6H14qDeSyXBp4KDpa
tCGOVNDXns39lT/aAp0o7TUUHkVdKZ0Zk7kt/YABVzG/i6eaoOrHg0t/qdgibO//2128DIjg7meO
KuNFVr9/IbHBQjCsifl0dIHvI7hKdS790QyYNlp2fOvylaHyCskLyn4BD6QPdwyD1NufdjMuqFG4
TveXggrd7E6sOC2nFuDCv/zhkte2ebeToOANJKX8+sBWcJZpf7lWZmpcdrOsQXzJeOOSo+PjuXlq
7r1DlaEdr6N8mlAycwVJfQw+0YKDG+6L/BU1Qag09An1c/jQApENvW0w3aDl/qfs7fpM87yFi8lc
qd99mZoomtDLYYYD6xNs+xLqYJHXWm4qs+S1II0PDa7K0+mTp/6rCn7icGPMZiavCYKdnZZWV0+t
pkj1mk7OZ4RwD8gxO8MbNODqqzW8ptpzVQo0hPFMKaFrY+EtsXSw0DqWBU5hMWyPw28ZNOcjZnNX
iXfGcU9qMvVIkTmW6osLbZOvbXVLi+8JgoP00NJh3v/oVhvcBfAh4ISFY/clfpmSxLLP+9psGSgm
Q9nWdQ8WUvb1vmQvdPaeyx5ittI/pjmS4JXQBf0GNL/WYbJKrASY9U0i7++UyJzzGrk8lpmL7Ab1
GcM7phVI+2MG/nu8EGVNG3IdbtJu24GDwAV6c5ASW7zqud5Y1JCJ1qZiA72E7ik/k5AQ8tik/ulP
U/db5WRUM0FQTJRtPFvQmWXVW3b+hFr18kxkdNFlJwRGg/oCskihBxPRxdA1y4B13LApF4S7vyz8
0i/rHFFNgZWF5OsmMoyYajBEHqrgKvw4FedFJgyBVjakFS+GEmy05y2/oiFct8sI31SIO6wKxS5l
3Pi0Rsx9z69OuN8zPdfTDSz+1/Tc1s8NWey9kN6w+dvMmaGymSY5ohSs81IDBrAONVsaSmdxF/ti
7DltI3EQyLDfWk447T1OGOGPMDYRy881nkClMHcIjtvzGmVN0Z1EE/4VAaA2LZc8Svk2kAwDfQvM
aRTBs/ZqJKxLDi+u+9IjVa35oa4rcUOqa3FxjSA7/kXt6Z4HesrjhqY5M+3GRcphaHl8in75v+vF
3vYblbC/uUxSCv+F21xL69yqsz0rL7VbNg2JgGcAzfrB8yV/e55Jd4EU5AuJEyk2IKsxTgOtNWsx
PQoXssd3lE5YMVDYH/04bCJuvdgqF/cjIYMVcV/nJpC5aEF5kObzwi02Nfptt+EGxAeHY76mNuPI
2CPiXVjnTq/bsYQwgy9kUTGz/zThEU/JrKPNEeS2/xZjCZknZ8qrw6NxbKuEQog7Xio1yOi8U+q+
U17ByFizygimZS9MzqNks3t7cohxA5oPC9W24wi67V/3PWt+ciI+q7TyfSakkRfxyl2YhdMV9XzU
PghTSSniQ/CMceud/7J0NhNyBOvGF8MIDuUWQFqA4FhXr0s4UJcv3NLFlPZq6+orbDYh375FSiq7
52ZgMNK/w8i6sIckniE4+BgUBLwXd7ln5ZmK4kppKPYDqHxxIxG+yBZ+13InF1EOO+P16SRPqsc3
ZAxPq2rP2DcK949qutocxT82dfg/08u/zasSfjnI1izAUAzs13gBjuGrOXp2UVgd4Kz4hdlC08Gh
//BLG4xr6pI0uPlIT3KGaBIzEOOcAlDGSZ3uoYgFO+BCKR3DSBbx3zCagNsatHRhPmPRmaSCSCDz
l+fqK1aKelnopogTZ1Dj3woXivsXRD5E2yYQRbVGl59/zNjFggsJ51wXXjDiN9afuaq0+UI40oBx
4AfQbTLOeVDG9UDYHnXaHPRhVIYCyTKcMPkVgeZF7xWAnznHTP0kKz3/pNsQYqZsMOTH3LlW7fxn
N/uZGuLVq5lxL0vpFMYhSF2euSB8nafgXaiYOgNCjkAOyVQOKxn2GFwC7Pmho3o72FoX4NO7Jp0W
NvdqqrEOnnDbs4iMn/QgvMVcb1UfMFoF0fxRN2trc5RP6A9UL7WFWSSh5/++m4oGf1EmyihArBax
xO1cwxKm6HlQPcLedf6nJQYmlqJsaPYUe4Bn5sPomvHlxwaQ/bwcv6ql7KTPeJgjcrEV5RnrqJ30
DX8MBM3e9ODWGYI2LWQ7wu3/ufz2FdmfogGYOlaFkYa0/jM1b8uKK4rIfJnGliLbHgNLTmAWryYU
s7+/wMSm1z8ZFmZ7gV6BXV9H/0Zp8C0v5A9hnE1vlpI9AcfuWGgN+yZjyoNsYTE+vFDfoID2aZx4
ht08RwgGWSEXt4wQTiADRSM/1NoIfB7b5N6I26V+CPBKRCPgUEcF6mIjzllWH2NVBMdip3sxNnYj
tW19bgOVcixr9sHyoEIv3PC1vrQWM3O6EFUl2hLhp/TLGp3YFn4r7P2bBS+7YYIK8wLAqBY7wAY8
fnr0fFBD355TuUTm9ej62C2V06C6z+o1ChMdLIVctF3tlexPLgT/CycnoZ0Nm3vk3BcBfLmd2XTt
Piv5WCzuPiToFxA8wkKEjSQroounuZAD9NBQOFhYbdrjCkIh/f3YzXuF2d6ehOnsVM37fY6FdjN3
S9fY8wd0NrnF4LGjiYCoHM22lj9iF87qJ03rFpZCYljq9l0e6Udkp4rsSnokebE02BYZ/sRoBZkK
EF28uwR21Hne/Gd6M7d38Io4kWx8P2+G7t+Fp7sb1xX1Y/CYGsxl5yexHBttLIsWd/Cm0LXFR7/j
lg492hyG350zPZLrRfL/PeYjzrLDLdseEZs9623NATIRuAE2JdvUCyWllxJeZJv9jQ8fiQQqHkeB
QiChJSMysu96pt3xH27vIY9YHBFApufg8S9v4JWCqKHU0bmWQOhN1ZCjRgMyDcojjHqwZbwVTbhB
2n5QpjO7muCyAoWUuSsPkW3QFOIlxnwCEQcueiwgmoeWFMZQ5dSJQkh1CcyuU8wB9EsXfEIcknUd
UpaL4XM2AMTzeLCCU45g0Q3tHW+3L6nfymufs79JW4nqiPY3js+1qm80GIRjGotNlePx+bccivKK
vUM6YHUMAQfpzVBSk0mOXIladpV3kUhJMREvBjR7tPj2malLrfR+H6e0Ks1wX2v0PRqVhSpSNxpd
nbzrsgI19KLQRTynmbHJS/Tp9q9N0IH9MCYgfNsJWhVgOUYByEhvOMP2kwCEczlKcjZ51xqIniRi
RlQ5f7bEJKlYegdJKNDbM0KQFtZl9SlPmb0Iq1loBv35B82zV1BxZOcDdoWOg/hoYHqeg2OQqM+q
IFxeMjsgsvnlvrpDcPdujJ3rFH88gRy7XTV3QIXx8jclkSRR89ZaLQpTtIv6iIC0XddTrWKswaxi
/RTBBORYieknYFU6+xSyCblGpc4f21Bjme4AUaUWtpcOT9JDpxoTyT+6C9SoQoqjK5+7OhXrk+W9
Ah30pn4heB+NrXmQ7v4JU/I4WZpGxTK1cKbYKk12lLsWnVidfFTYLZPCT7d75E3uwvVEXWYEdfD0
WzIt+VdATFcJ0cv1VEtZQu22E16tbitfm9zFaM7riWqNNsaOWsejPV9TQPWLZITCODbUhxdaC5Gb
+vX3qybKy1/QES72hhT8rZ3fF+lDwEu6JHSwgyn6T0J55+g+dBrPv99RRRxgGBkWydZoKkVOo9dF
iPLEFDjhzp9ICBiNqYfObU5Z/t5nrASLHPYAVBnrVDhc+Ztp//imPabBFXGmmU6/i9tf8chNVlpV
LyYFaDOiuIEKZV7bYxVonzdPmkMGCGNS9IM7gtAZ8cdTHb6flU5qlqhsLcKiuKU4a0/JBkmkO8Qv
GS5z7jddsZvXvzjcM0UsE92SoK3rsfbkZWKJqtdivx4UFjCrVLMyvvYQAwPksuKQZfuoeutbM6Yl
BbaPkBq17EN7HARcsaQNzkRBrexUi1+N/ZpYKdcN/JUxUG6SKJIE35vZtTS8uBIGuu7C01V9LTw0
WfFK5m3BotwcdgwCoVXQ+fS9UQqHMaBYAdRu5OWHIk1tuobcFSohhdPJIiMFMky89ctU9kZPhBpE
uI3iqbZ9MPr8NY6injbVxDQmpQcbhr3ByJTLYY+2JQHW70mwOvbBRzbzG6xh7rKhtwwTsd5DV8BM
/56fIn782VRmq9yQxYjNppyX/64KUydWUSEOaCEKhxpcUbLpzDz64cxk6culEb7kOpy/gIB410cO
8jeejnsTAE4sTKaYwulnbXPMXqoaqaLVrIiMWsFqh9LEoyQ0maAukBLrW91AZwSHNMlh9Lam0XjL
vOV+Ex0lDPlNGRtGaWqiGOxQPAIbLV1OWIFiu1UzA6Ne1gvuMTfVZb3MUG3bpC5iDJ+NHuIirzGS
5kdPvrx1CiGSCKjJxTKlbl4J5ZZUi6s0wCld2yAUznEwhToIuHmqXmvbmvQNTLeImgDOqvkKP/lo
16e6ofU0iNFcrkjfi/mSwt241GISMQnuqAGZ+eXC0/VDCSHrXClq9tbpArYx2gNYVHoiYZ30bc7n
ipC3HwO8DuxGkmjeKzkxuJIRS2hsK69LeLexliL7zrgOt4w1AfHAaIA/168bJWp4R+N7WSMPcAOh
OvkmGzAKiFSgoB4spwXGEzdXqWELrtKs+pUZqeFxD4zQFVRl4NNCISXpsR+0MGpq7kqnsSrd2YSm
Fnn6nFoeA+81BxrBXiLHYo2a+RCajzc0k3vl0QHUQzWWy1efr0M7VpX06Cvka6O34iBqdTJyrEDG
iKLAL+9Rt816U0RhLoP/Z9Xdq6r4r5TWjHzLTTjm7mG4dJ8mcI6RtEEf04OTx3esETtpE0zdtszB
isVagV+p6ZRvBUqq3GHm/291tQNNgvglbZoWO/QAVxa03mEGOAxkTIxBYHh3ycNn4OqcQ1aHq5kr
Hcc9vmiwDlNPbzZ91QFk52VH5HJ3sxEC+r0Sgv6LmcYcZJkIfKPj1Pu7R2uYg8YOWfSpUWUk19yr
y0U25MhqLh87/p7MWKORgfnJv42cm0hHeuEim0fZDrJVPG8/K5soTHYs19DcIqRcX74W03eAn3BJ
E9ttNn7E0zn1D/FeeTKl+r4N1Vf7EmP5A7ggIgCCVLx78UHFcvg1KI1OXImC2TXClsUYUaHs/DYs
LYDV1ItLCftppgsG8VlyytFn6t+UfTn/qe847qt5/xImjg19tYRrG1rxkjaw1Gc0R6z9Hn55ivgN
70wRDr+Zs9X5b5GvLBQNE8a5YtiwF1sBzM7Ubm3FWQXQbdxKf4kHrHINXCODKo+CFHQIP4npru1R
wLyosUjLI5T3FF9bOg3GindO8yCh6ETlToPgFQ2SlEvPzawetcYH1U/a1XTPQdd+b4lUReubin+7
C9hJJobVUZn1iYstD+OyKAZ20OXsJI+Rzayf+1euRgPEbVZGSS8FzfpoA/ekMeIQC5wIilk0RTb2
Ap/PsmbNlok+AdGeYoV/qeWjbNESYKFpB1hrKe1L1YA5aDUMgnENjlrF85Tge5Hhje00Y+Id45mY
gstd/DXpwSuafhmFSRt4BRnUaMoZPxZ/cT0h6p2mm8nwEMFtDL0kdksQnXw99RjUYEBjGT6i/TzH
josgamIlb6sWV2MvAzMOLw9nAIpq7hFqJETPKo5uYkDLvQfLP0sDiqE3UZJK9+WmZPC3jCywr5bO
OQAcQ3adDBDXMgYqFBkqD2JHy7gE7FyQk8+YEtBTYwJj0BNF3xlYQfrauBafYt5bqBgWCgu0+aMT
7FfXTk1ZxET5eOWDh0qEriIoiLkghLL1KukxPZyChEiK3hV2oiyI46N5Q7d1MW7P3tLVpkw+jgOB
LTyQdvAtg5/+WjztB9w0PXtqkXAWHNwvrjsVHJ7uy8Av+EuGtrVYXAHIVz09zpOBvtxPzn0XUSOL
7P1m7V+yW4dKf+EpmFgfi4IRtEnU18Ml6jDLff0HiUrDuqNXZNK2cHRtIV2Dyh/uHgjIY27urE80
qguhnAEXJXFfDBaFgIgFIt2K44E99RNVko0gNalceRVqlWL1AJSbnUC1MdVpPyYKdH0O6tZtdnnh
f4yXeEAiS3KDgoUmT41jjUyHjZsgAVrLU4MsNAmvpIOrLeCx2oGeTNS/akPk8ycXwNBPz8r5WneU
YNeYfH6LG/WnYu/ztIsxhyneKNDZ1lFTBIX76ZqSng39nFnIaMsZUqpUZ0aSs/RVrav2XbFMiFCm
ZF+76tb8KwvSmqlTkCQfYvMpt7rD1QlRvKTebggi+pq8+FxEQ2Ol2gJHFDRso1fR4/HFxCj5yftc
dfYGtTXvTtihkZOx7kpo2H7svKMTt7S6grYQAiY2n/OqbouuP+Ptv33cYRgReKyHf44hf7vXsWS0
WzlbQfJgZZOpFQYSla02EFoOEIUwT8TDfKh8+YTv+hCnL3wyrqDOUuliWb07pu64zgvWDv5QzahP
WP5eNCfrWp+2DTYww16C1WQoV2ccNGQ3htzhX9Y5FphZAwkjA30V79lTPL6NCubERP47189p5k9Z
UOKn6wJ9u3qMg5KIaJvHtGs1jmcYyDz1spBWsBASRLbjj3cuBGPCZGRjGikiluaP0znSI6Q9wMGP
M+R5yA6JRH36AK0F2NPfI3tFG3ALdJv45m7AGNzvcGT5t9rOsfZe7Cu9xB6MIDpAjXMVYfH9MqXS
yENuYBCfEsCA/BBiBGNl/+Nf3mS6/KipZPhphlwgNCrQZsrIr7FvO+iUI2lP3wt/kIltovgZCCJf
EDijUTC8H4B4TeaAAY9GSokdxf/SyJDHAY4sqlFfCenDoRaHkVQvuzop5WgnFq9ApyjvYw1fsPI3
8q7OB76MUKjUm5KNa5SlYJWmUsa+aLhacnZhzT3Ovip5CFeU+x1LV+Ugtb7KreRsa1FDhNmVXbXW
qr9iXoDJa5eUK59dDFNFUUxissuI98rBYKZ63rmyrkFAvCK/HhChgxzPGSl40UPU14sJgT+mg8Gh
r2r9fcFl3bdNorF3DpmgY6CB1nbmRkFm/YGhLlWVHXSuID/C3MMidZh6A5CXpdaBkPZcSLrM1q1f
5uM+j47t+gX9k+mnPipvOKAQEap+/POrpdgyFJ8kUlx/lYohqdRQtULPGSe5uH4/3XsyWbfTgtUl
0kA8bXeqS5C4Wzxl8mdMpta3GIdtm6yPWv0HfQKBgnawUvDYRk1RVljz9NiAraPSP8FVO6Oj5AT9
SBNy6phOMEU8FwP9d66lbYKrv8hfIyks6hhjjKOyJ5w/QrkNmGlco/v18a1Oe9q9kG2wxX6vcBzP
vL1ZLSrWZvDF0PLXSCRTYCgOehChddCo7uis3sL71s4Vv1Q/7PxzkgY6G3Jy1tJJnyRDRqKe4B/L
33pnADIqKPYzYHankKcc7arAECUu3NwaZxect/p2MPLFwIrvaziMek7FWLZqJQL6ZO8gXWUyPzWD
Ym0JMJV2g7s6x3pEzF0g2IR07G52RUI19XC13HuuQ69eTRnfkkbXZSu7G+zgBkO0ag6zEP/R1DsX
uwhL2ousHnEZgOzfiopyHsDIt5pX7w+mYDRw+VB6OQgxayU5vi8PuS1K/dlUSnY6erx/NBfDBX42
07zsJU7szpDYQPIBwQ19gGt9vw1Hm1p5jfk7R+PxVi4UXQB80yL3U7BNHsjjbW6QTcfOe7+t/0V/
m2Exye5mbiQ2CbAZdyVfIu/mdY13ktjDbIhqri98NIaubjMggof83dTBauC+gfGA6cZGbetXu2YB
rxdAk2Y0wuVynUADzqpPiBN6DJPxMc8oomWEZYvgqmkNgNDuGTBEP9B2UFWAjhcDDTBnhIKQ4PJ3
jotL6T9xJFyf1Sq7GVz2e4avw8tdXt/yRMlSHe6ja4Q4uBvMfzXDqat5/MNOKT3KeGFkm7KJQTFV
7MtBVo3ZTzqnQuggWnsrtRFfdxzU3xJGTKoHM0LwKf51kCsdw6OnisLiC3uwkvUl1JWut8ecqnJt
vUxhV7sPjRqGhgsS9TjJrbL3DkScofC0C5XuZ7uh7nvP06b6Rm+0EO/H9LCQZQKSc6sgBUlJBgq+
UjSvKCPPzYFC+IQMmFc7PNlKZhEB2+Uo4HqEXA3L+JFVs/mpO8XtfzbxYikTSlh7M1Uu6fbpUmmR
ZoNSjL2lSWsZKxngf8q/eh9cQ2VFZLWFuvsk0gIE1EPB8vnclV4+dRIzY7Sz+5j3t9BPUDfk7Dr2
MHj9K+CYavH5LxGJULv6EpszfUya6I7tEBy6VPNDbGtmidgUCPywckMA0rA+sHbYsskLx1HeV3Lr
FUAXw1fJU2htvd0bI92Lqrp4iz5Aakipn4v45kzDB4HhGN3+8MnpxEOcA//vb83XMt+zKQB1lJa8
BR9YY1ZeoVvbEgUdTzFRlGwolj33RWdoCEMgUsCmpVW+/GHzugtYMqGveI/G9Bo9eNEbSZyOY+Ax
EBU0VzkMTP5GUy3hud8Z6pvwNk2QaKMxgmSxC7v78YQGuAwDf0NdlIHrLN1Oo/s5Svb93Alw8jgz
jDQYzdQKDprF3fkeJO5tvKUNnU9DneruS4SRYa2CCS1OAdkaOsoE4y6scqVqolZCA/ZJqJvfJZpM
wXLlwaPHFulLhwLx/hw6JrjCWu+wTmN36f2rokNF6qHbPafHE0f9YmI6JYUpR6RuYbMrWztpt3yy
htCmyS9+HujYlEc+iIye5G0PFxLcJD81Df1oAyi50YFeBNtGO2MvHwt546Dgndn0cgaiMH+juAj0
SkiX+EGsicMI2+nZMweU9IYG4v0QNgWuCoQAI10IyqKjlP9Ex0HMGNRHvtHn48W8VJGJacPyc2pa
MZDF5Il1AYtfH/hdFDxhw5QVvaXwyVv1XOK9/epW9bpcGpbdtZpY8WcIfg3H6Cex+V/0Ra9tjZ1V
MZplXIP0441e+kKdMX3sq8EEZla20WWGM1KEuo2cVbmetSIzZbeoXh0uxVT5SQBrHXFcrjpx0PnV
MjpYrLFewK7nto9JFL15NCep0K9qZfRtwJnLrwEG9oySrhdDM7GfWhwardGPVE9Ok1hDH9/ne2b4
PbE1lthwNWBzkjKF25/g4++MdenmqQ9JKnUi9zoaw7KUBX9mcWL3MNElvRZI3fmvL3LVJJ4hGw6D
/W1QvyCBcGoPr5X992oOTvwFM/DeEC9DmT0f9+fC606bv4jh/y9El3VRGeV5lu5IFMoBtegjlSTt
EKvxtmcEMF+g0n0XUZMkgpp9/mt6xzn6Ro9M3657BIbSdbRsYiarF78srC8mQI5KwPDX3rCAQBMd
eebo50Zsry/FeEKds/d8+R/du0lUEhpJr4kQnI4sMXTrdgk0nTJ5fyp8CwIOLFPSKaCSriuXgAP9
9/hvxjQq52Xk9bauW26algH0BOSRyKDtCw1eE0Txry34Zw1QLe9DZsG66RyqzdWs1nICGF6MmlGp
+p3pZeRaVwNpI5bWeVsPnCsgMvsQA+a1tUGOmmObYEXfIDAdCqcR16w5rQriQaz5O0n/ZWUvx3Ps
U6aUHftRWh0Kip/pQrs3OI6LSm4qxdBuNd38kmCY6nKBsy51dzb4LfMWQohsDHucuYHSrKQad+Ps
VjMtPpo9Wr7FzN/tjDOB4S0/0CKpPOsPuk4eza4z0YUCs6CKFKQ2QNJLQ8XG3qDfbgGooNhSGfM5
KnHgSWAaDhbgVG8W1uaTC9zztails05E3NC3TP7r9V332XoELFyHQ4+7eCW/WYRIbjkRiGUhrbCn
k6Dw9j06a5BM2LRQmNKf7GE+dH48RKR14kSTEb9T1xtnfdZhtOShLEmob9Rr4uNaN7HNEN2ujRYD
fbvhNUMJ/eLSn8CDxLarpjst3jRCLodA61HLFZXvVp5I1DC+S+xU0QII9FHOJKb//be4tMWo24V/
qGX9ZKVV6VBUH2j4HQhZZZTvGLNWVXcHgFHdSCuy7gH5lThtxDisOOh9wIBRDcEif6NBTjcthXs/
lOJ7a/BEZPVDooeav1wkG8Bm+/DLcf1vflcjXeQgFFl0ey3xCFpfa/Gnw1wviDjU9kieZKl9UbFf
kt8h02PTZh9DEygeGKfc+d1p2SWs3OU0WhVVBhQz+m+fkWaI8RO/qqPYMyw8rahtEixbMDHmkjjA
J3O3SO+iUasXdM9G9A2PuCxJok09xWSFE2PtGPxovJoNpoTctbqOO1OlyhATAT5MTpIaBlsbCWTc
FvbsMCCsRFicOYd2+DX2CJ3bVeKNHoqk+27vpYLyKh2wXI0TYyND0oLmcL0InZf92MQWqG9RtY25
ZwGvx41N1jJeEyvblH/te5k99glEtr4UGhdIo4TSu76k4BzoMys2cvFVZBY7Nrf2GXz6RN5ctSwJ
+ZGM9Q/AmykpGIgnTYrIoXDBGLaN0xhG5FEIipI1zyprf1SVIlKePP3fkXOokKpVToLWQcLrdoej
JgbM+0WBHTp4TYm7nz8m2SEEznvCDgH8nKfA5Be5uqOT85RdF8BXQZ8L/g64vS+eNTUo8lzLteaH
ODTKHciIoZ53SgAlU7vrliXhQiQeocIOufw+E8S7aN6MrDElER2wzD/VsG0lCewstupSobtNS+Kj
A9jvOV60iv1lDKc/g1y72IP8ZbsFuO5lfGXTAYaJFKPpVhXW3OdwtmO9XRGputqfkOgPXABS9uga
87vgbNPmuozzD2zmE6CJ/+fI7oypy46JsTElKegBaWXjsXLr/ylyPMoQ3Tnhaiaow05pVHkCEvmI
n7n0IbSVvv3F8AvHTn51yiRa2bsfn7wHQZKcnpGjqSTsRfn7dV03lHtvPXvyFZZW9KBY+5Swimga
tIbudtb3RM+C22pJmZAM7fJfdS0KkYmCVMLp4uQcX6MnenPPdSjGn0kia4AnXOEH48wR0A8x00dU
JdrvBiH6nSoPR0TJz/a5fEf2yWhP/9MYg9YiwjnQwvtEMLe0qChpHrGmzv5lG8OwitoAjfEIOAML
mlMsTEOb2yvNeQBlwjc87gionSQ5afAOC9y8L51mULzLhKFTYsaizlX34SbzknRi2dR+fvtqaV+L
yatIVsulFDrKF4I3JEst3v5aS2p3K3Z0IuV8N8YMSQBfot/5UrEecJazwBb0xCU6tamYvXq3f++X
ILGXnD3uXKC1kxOx2bcKD3VbO6B8jW/2B21MAWIHlzSB9lR0DhmQ3cIY4fLPpEUNp8cB/5nyjFoD
Q0qFoq+Dw+evfNBQGuD/wa5BfJG7545mVYeDIZ3aacBHiS56UWkOcCAGiZfnNilOW42BjEvVPdR5
SM/GzeyvdJ2S6wpxBY6RQprqJKHwLxBrMb+Dd8RMGtsviIJFLPbzNLcGrbChOnyRMDDQ5WC8VnzB
0ZmqJ33mrJSLlxVSo1RKOyRMcZ+fo8NJ9C5eT+td8Fq/UH0B4tNC6EFnzqLRa0LzkXZt23AMWb2N
yFYos1xjRJ8ouvbiwvaSk+2Ob6VX/zNF9sISFVFLu27gakrvQ12PNwL0kCXQL+cauroz0iwP2I9G
NHQ5epmNjA/gt6PP5g8rbTMKIXiLDM3LMTQecKbdB+oBWMBLoe3Ko8ev3hLNg4RKu5Exwy8YzwzW
RVAGxwzz/OGgErCegGa/+TM36jNX20/viFHEQ6ry2mUTjxIjr6J7Xv3IPuavvvcabdwQKFNt6BQF
W7oYBYKn91CvZafU7OEM8AW9/XpulDU2XKEz5et5aO094XEg0cCWgqFFVGz9wa0HUdFw83M9aPej
Kwv4ygCEkFpz6NtLqBkyq6KPk7HsPcAZbdzOW0wH7cmjgy9oWccze/F9NJscaQCwv/DCqZyE7YL+
8djiwkcHVqci++p0yWi3e9BF6EeQyWxznzadeWx0YfCiUoAZdDcPCsVkX5EEWzavEps5E972mKqE
0WphOPM6P1DjEYiupBGD23389Ll7XTMUtsJD9hw8zqtt6wgW3Dg2upSbu8BG0LCSXjG9sXcdNo+p
mpd7tY28+tXXDW89o5JCZYOmyyozUGIiD7/WK3A11yyGtlau/cx7fXASVbyTjNY0Zfd+SWgMOfCi
e/rmIrkewimilCsR/BjX98LQLlY4zn5sv9JcggISvoYUlqalwJ5OQgUgxVYLU2nOUZM2Zgqi8fYY
7TdDcoajAKpgjqy8OYWzOBkz417Wrly8Z6aoQy1c+0+Oppm51X1pjs0ma2ygQpzbazIQzwjFjvaM
lY2T6wr6i1Mp2j7KBDwhbl+v8N8Vtm2Fqy7LJr3idjV7Jp3oqdzz4tzWMzqDpoVtVdQDGDaQcY85
FxHH36f3cxKKSkiE7MWWsewkh8s7ZxOL0ynCJb9v7tAb0RYxntWQLMQRlH5hIQ2bYhCRb4rRuvLW
twH8Aq9FKfkNEzuBmdX/Uwl8dYbHCP40/wSRPXeHe5l/Qvg1QmOnLifg5IyhMpZl5ba11uNBy3SH
+j6fHYdnZ2Aw0XnK2p75KE3JH8IMk8KyW4LsNLGNaeNsVrZFOHmKw6n8UdwzEcUIO9c4x8MrEAKp
BBZnxDzzBkoVTPstHeJPXSDQa4uqcmPrhXqALs5Q3JVQop9irr6KAZSznR1XgGbEvxjCAshRlmnJ
VjZBn5Rd9r92307hRN8Ue6tRQ4Me3iPFg8Yj+bb/LfkwZV5/a2m8VwvMq9GtcsFXE0wz0N/QxurN
hpRLICfKE3HRlmfYed7y2Ta435EDDt7ot+zVeIF7UK8yPVyyggeI+xK23T6BHmZkGV/Ffw5z88iy
uELiWAM4RNtebvX+vFpXpe2KQ1HbQ7xzCSe2p++DnIVZ11OjV5dl1f8DoDQ2/laScjqWl6Vhx+ed
heEzPjmJZAQfeDKRHZCOgoJ+hvo0dHMLLrFzx6l/s/BxfZ7hvtk0ckrws5rxw2ZoEG10udwUcFOQ
h4UackShjQa6iRmraLMBnS1NpHFO+FuB9G/yLKNc62RdsPMr+7Feamcs03xmG9+WnmVIV4rmBOUD
Nld+lrr30SpwbugVmGuA5cK+NDZW7PmNuA85vs2Y7XhfV+NG3uCOu5j9myapcTCP94Mtuyg3OHgz
btOMLBn/f6oTvIog9tQt+2YJuYjBjdZS0jPgOjYbAjHD91I8X24K3fAVkaXoUERSfchxpjiafNXb
UfLZLsWGMml/BQjODgVGQ7p7d62Lk0+L23M6VPDoThfh0AuR79idBQT2Ln1PMoe9A4ozPNPaZja0
SUZGQ6OycKfVuVAoZSAm9hu0Nt8/ivdEmXBZubh/hPnmpoFmDm2ShDF/G96JCw41r2tMlYyuBvos
nrtq/cqKUO1CNfAUx0IaHuNw3sd74pD+61h7KiqtZiKYsIYlT5eIWZ74hP9rz+WMIO6UydI7CEb5
C0PgrAq+jGUES2kClhZFf/47N0RDIdm/v4kg1F9jCf/yYPm4XVzUNcBbgxcR/0U7knPH0iK14TWf
QRC9pr7BuMK+RhauBjmfbPyM7/m/mhQFvipk3H3TEL5sEw0GiCNILKlOQ7lc3YsRroTp5QxEBSWJ
TIrtUTqqGztS2t/jsokBdRFkqGhjU1iGkKMqRI5MKOHumo+qqZjqc5dKsL5cTkgEpEzIJXSK+VSs
nIWoL1kpu5H3yzwJhklr+u7jwl97+/6dFDhupy++JyKaH/mIRRvGjn4E1msc0bujoCARJU+nfxQD
8fxP3u/e7u+5PAovmiEiz/0HuuWK7Jsr/o0UHybfzTmnt+WYSCorhzoMEDXw9sz89ZWAqPxZ092N
D3l41M5LZiYNWOk1pzEnlV1E/fCeFZp4jyNyd1mjoSyDb+PzvkXJqMznL1AQW28Yn5xb7VyefS35
/Jz3/8z+kX6HtOTvD4SFRuSq2VoF13rc9PMr7b3Ey6C9F8tTosLMBli6lCZAQ8gLbIpmXRLnJoy0
6wbugHBMFa5lFNA5s3PEGPgrSVR7D5j8EFHnHRyU2fa48kcw6nMH7atgaUhF2P11xwdSTZ5flcLf
hyCDneEIhwsEen8Y7pJ5fE03dDReqoTbW5n6a1ha9/cBnFSVCDbD5kt+/d9FulR47Lscb80e2mhA
q+YwbgrkQeuspgrAudGP1at3nEQxgZ8h1Gw0Tm8BGnEg9W9m4bFjnkeKTJhNM39T897JG4iklez2
j6jyyRjrRp/FHQCTo4uYMA1CSiAY3wAOxbklX00p/Qzgcna8K8PT3fSSxY2PM9YFjxDo6rhjjfa1
eFq6mTtG8X8MvewBc27Banj34bFYlBAI47h/H3LmHqdDD5YItWVL5mfGHROUDSCWGi1/JOhjzU3h
+WJ0iS6oIKLGeop0KJhc6lPdbQIbl90JwdrQDbzg2DugS3cIgue/FGY0k+cRfo2eYg6+dWZ1VV5e
OW06GV1098mTrCU+PDrDr7lE8rxqnfZL6ncwXbPnvVWzSRJz7LofV865GQWAnIxAPY2/Ua4LK9hi
oJhbaH5Ibd90Y5AlhCAQRISczv7o2CO4Y0nA+cY9m8QTahz3aFpDXOtVflRyHaGBLNCT857XJkbY
n+GGSqiAeS9c1MLxtKBVeHnLWGUmQmZdZDmyfJe+rLJKbXh86OryhOdTV2BZeAjCEIFtjzzfJK6R
8m2XVdyr6BO5xF6z9v993CUOXZhofxuhvH/eC95/XrFBJWhiUlXWpBdfAu24DrwV1cBtY7VA8WwP
wfF7iR+8rcq1aZ+44j7plFetlurFo+DgHrysv/4q0y72FJYc8s7PLXW8M/YXx8TC7pMWSxRZ4gtW
akUOZZ/XKRg7NanT4AX2DgdfwTyb5OqfDEHx3J4f3iTza5/G5Cs5VGtPqbPC74jTjF4JzDUH80f9
hWopJIqaNkxnXUsR5A+8dhCXGf6F2m3uZOky2KvQV4IA/lgn0Y0JHN/z8SdnPXRs7WixEhA7GHhS
wpTDBgXpaKIHPQPnUSg6Go546+l3cKYSVwusvHFjDnP6fKXBfRhbjlTsUpLCkYUJjO2ZJ8h3/TlQ
sV1hNFWnQFkgXi3nGdUE1k9ABNR/c4xxLtlr+45mtVeS8ga81n992qvs6HpfrQ5rq9CHVJAy96vG
y8al4URG3yg05oRYefIZmE8TpE65EpSwaZRPFQjrcL/inlWFFc/RkPOqFSIKmvEjiOUln9z9vQkj
jPA62L6k+q+qW6gVcEMn8mPOYVXIpBYd3FHkFv5mVbJQhJCbUosakGiN7ZNzzmizdNpFHoP2+8DR
0bjEm60SUEuiXevVt4LgA4Aq0Dhx4XHZFIngRDZSpjdQIQzKLHvE9swyJNvxsLTqUZkQP/s13bv0
mV5R6rfR7SpjtnWfVfhv+aU2Q45lW3sndLv8vS/WOiEWV4OCLDZJYHIiMUYhfH/beIwKSu5/1Mnd
+5IloZoUR4x7OeJCqYD2EHp8gTrgcvtx9T2QVKVLVn5f+aCLGyGhUSbL+1Cx5/+JnA/RuvyzBtM9
bUIW+/vr8AO1EQQuPLT57w8WJQPZSBI1n94OdrwybKxlzaXienQd77Oe/PpwBUZbpJ4LV0DwzWJ2
bs1JIQGLUm80wYI+4+E+zBBuYHHAWZdjOVdHvwj0WdUQlsv1PrzCHayKuf7tnGCiEburTCDvZxhI
T1ncGjQNw6Cyc4JJcGWphKzP7/RsFfmoMbY88qSnLansenuIaF8LdOKMd9P09wFS51P3NZ9OLdax
RNa+xIxGVYCDIz+e54if7WFDeno42gMQDIKh5GsKY1PxJT4T+BbE41xlVzdkR5BwHre0d0Kfy0PR
Jc6PbT/iwENWdultZ4WcGSrWQ+dTXHt4iWeSWh8kMNLtzGkg9ihPN9WRRkshL7V6xF/XSjZx/z3G
W1Kz5x+M9wMmSGKUTsi6diy2Irf+WG2eH/B9f8c0pMU1x2Pi6c0TPBcnqKT1zfJl9Q4eMLUwf6LX
/9pA/i8ANj+RE2Qa2o+epoFvAEJY20dbukCuczSkrBRVhpGQ+lyMbaI1pPZ7kP1TkkxkDdOgfVjf
VM+YXOT/Nk2eZWqyF1tGHIhr3msnr2I0OH03vAOEn1QBVCyH+fuTXtyWWG2P/QcwMQ2qbeK3E3ce
eU+KlQCYWFDpeonVzksXxAk8p4AACvpLbtOIaIiwmLVtM0xdkElt3nIJKuOlJnToKYxyVNwrsFGZ
PDBH8Ao8OslEqfkeQBf7fwLKaZMIntN+Ra9Kl/7/psIzbSwDQrkrmEuLZE6GdC8mlAFBfKj7UWv3
LgvwsWR+bGkja9QSLwljzvhba3Z0/+QiW1UyNmAEP0TdYTNCBjaXgSHpnwHisjsNSWWSM47GOmw0
YadnHXL0RvBHd9GHIZGkJ5fKFqmC51JdjCddgQC6nOF7pQdNs2HLLXiKpwqAcMy/3Z39eHTq/+ZJ
8wirdYqn2cdIuea24gY5lDjTSacTLmwDXuz60yEwa/36gw9QNUWFZVN8KN1BXgxuSk6vZG3HVt5H
CxOLf7mAMbD9MgXtc156A2Wk+chH81Tm2DYWljI7FDVq8Kb1U03EDntFiUT1cd2QE8/pLAzB3AdI
w1MZ+KQk5HsxKqbUKtE+A4KMmC6hitvJ923qfb3sXBnQpzzwYtqMJG5RHGY98DssPDrTnBqix1XJ
Rv6O8fEOh9XUTECEkMx8z2ggbqI067iW6np76gfTtp9WdW7GX4JD1OAUNHFpW7sTQr0cHOVqrQvd
qPbqqb/6D08grAU9EFhmZW8xmi/cxvJ0RFMxkRLT4ViFayguVx5WCUXKnXyUmipleC7wXOsTvHrs
TQXgINW7gsv2jIeH9pEMy8NwgJitgkDqXydnjq9+KJWuMHDEVHzQoi4Y+GqkK4OJh4SUZcSpaXyd
Qn1O10PPpy9o3uKEx1c4Twc5bvefFv6jzFAuWgxtQiCQs1zFj72cK1JTZzbOY1WUHBiRMD2PRC2b
RCDe8fQ8UiRYonXPCypiQ0+bqdfWK4uHoXD84RCcRUV+NrVmrnTZyXUC0bVKtnEPKOv7lvHQkyXA
0ureKfISDctuuoXzjwIWAnm2EOHgZVbxnS/qinCfmG7u2Kj0mNhDgpXZzBfY2ADQ/8R3YvYb6u6e
edYl1+UOrN1jZNkBGtFxbgNcb5pjqJ21kQzcHW/n9eZdOr8sIWlzY2R/mg8sOXAmdThAJhpSz1sl
Q8XLFGkVW8AGptMZNKsYRXoIJw4f4fTOtuYr1Lr7NVVyBpU8/gy7B1RHi2qzBAmvBF0+TVUovMnn
rr5Ldum1h5xjWyPdFz62EkeFY9Jku83JplPGhkzm19IFiPLERz4mU1DIgaZL/3PaNpX+lTIb/kg2
slPHQ1kTU7J2kgiIRus7OcqKge+lPOmG9nlnRKLNypL9jqzC79d2DYxuaOLD30+LdbEOsTctWca6
difjIIqr792ipYKRdhD4H5RIfaA3dm3gplnW6ivcHJxfp/orS0je/C6unQBT9hX+XIXsFksIy8mT
qopGJeKbifW3VHMOrTdaT7cBuNqIXVv1k4Y5emuxdKPdxsqPsHy/si0EHFceryiymrg7/d0D1QNC
EYCYXW/Gc5IA0SpSKAs7QDA/E1AZ7M1zWzGIdF4eIUNLjpIeaZlJQQxSKswgrjblv0NBeS4pMtE5
/cjuTo4TYbB3a5s2nVAYHxEy1CkvcjMkuE+iM4yjwEW/n4VWBlieEd8rUtv5Cmn6BaWMAZCaremD
of9sFqvX/KY3qW16ZReGUzS2jXvgLlj59Ablpx1xHbjurGLQz54vdBeAxsnuTqTrucRQ7IYNUWjv
bJ6nIkcvLigYzjJfhwee6jCTkaY+D8Cpdgz3zgtm3lqIcsa1Owi9zfnnVZvcyo6+r9N0T43pDajY
kEYWUmPtyARFG1Q83rM+ZQpnWQ5f4crQHfRDb5erelrP0PIVl7zjG3NNpJmw+25d5NPD7HkXGx10
U/5ABE/RKu6+VKrClY1gy9I0U47xs2aotSBQwK1NCA8E29Y1kSJAJ4Sz2RhjN8GN/iG1iCXspBE8
Ff2OBBzC1qE3a3sFYgsA6niJQxuff67eKlvZVFA5hmWsebmb1buvxl6n7ENipHrln1jMfpK1JFDt
/L73+pkoR7YSEFBK+au548sdyvqGL0wy+A8OAmn9s1Swu0/vLTKa5XM3vS8NkmFsamanU6iymgQ8
a0rqXGQwg///8G+7p+WXD8MshzTqpQ28+Bk6bMIcGs0js4JSRX5e5FbIePweTd9hZ42FinRz1hW+
EPzrmKW9/bxxtgGaFi8BgWDa3qqUX1vHUlA/3VqgGDu8CC9gXE4CiuYaOlfU8S7R7yCm4HeC6yQt
K/GMjrDsxRK/0jQkJ9fC/E5QlhDpfimNeHewRbr/kh5a7DwymXOQEy1sKEpozMrr3sULuqvtn4mU
uazgugHogZqFS7MK5n+uFpnvQlE0ZAZu7vIoJj07J0Xe3YWdI2DXp8I4wvX7CrRI1nI5YbPZ/N33
suWDJY1TUfS/dwbx9t+4UheR+Z/XIL2DBHkLa9nLYwasyNtCDkEtHkpGgQVKolJKghJ/fSWlYHTJ
M/ObkS7uSxiGENNPnYH8pcWfWhDonxZAuJ9xZwuvrWG9OP0siqTueo5CZ0kil5jHKLh+Bb1CbdnG
mmElSXcl5Xqk2VgBqR9H351Xc6TlFBTSVfB4C8nlcXx9whIwEty+mNfIsLMFBtgzgRQxRRBAdS2r
6a3DBmnAqYjm0NH8xHqn1XGiq2BHF+VJc8n2qkwGQU3/wgmv3+B+n3RPUSbLBtN3XxhngIq1lqul
BuIlet7uxw2yBB3NEYxggfabOoKSmj4/xdNvNzs2m2Udt02oRTk4vbGJAEo/TPqA6LQ3rWGn5Rll
Puo+iGatyRhS8mJKt9ynx/rpciiC6lpte6eXGxXGmex6WhmjBqvqAadADiAyt/LWssuluiQnGLhX
vpez0M0jjjE6ztutYKXjxpqstgmFMrVHNm5YiTN2vrREb397xgHiGq51Z5m5gPz+TI/iuZQliXpr
vDzVBUbTwl/EoUTbElV8p0TfSG53xWeaLBrb+dp4aatDDt4KmZyBpqJVxPO+ucZGt4KFMgUeAIyc
3TeYbEcCWvCy6oAfjVI9C5Ps58ZXsGTqWsM9wUUYu2CMHcUbB8sGdxdsEnCY67nBpGTauw228Cve
liIV32Gr9v1fbQBBxP1ysgjCYK2kb4/eH7q8RZjqOsNzEFSXMtok+ngDO7XZ8SxRPHXOx9PTirMw
FO8fZyAAfYGaYHjLl7y/bTf+OHUUKT+qGCS+eSu6M+R+De1bckxk5P0e8YfbWCJt63K8dkK7KN9q
0H0VyHxzyJY2TV7/YB95KrkJhSLFmi0i7YxMU5HCWuXGeH5cBTGMbsaG/yJUFqelKN/c660X1UKl
ZZ3f50mME68RlW7+jJNIrON7BzTEaXiLM05sziwN/gKSGJonmjtaHbmj8KU2p9LSEgshfcJGt+KF
SskTOjoeeFiq7WANhfTVLWRrF6+67A6wvppf38woNPNcoXUlZ5/D3Bysj0hLRK0+ci3N7rUmi03b
+GSsaD9l967gNuHvoXFe6C96sSenUTvonRb6uDudc/+PDY4T7GgWwy4LEFz+oPYP/l5TI5FzqSgz
I2PuhTavYoOH3DnJr/lM/jlsAx7MkhwCqyAB8Ze5Djtz4ldRiq80i5IZMZ8JBEqmnx/c7KduqXp9
GwySDa3LbOpQTh4YrfHr1G3c9IQu31ObfNYmfL9/v8Luk3vIEFoXnUv0xaJy9Da2NmJFeUOWKf1M
k2vx5N3FO2KRxMPQWZ47H3MfUPyBB8APp3xwL2Qz92s8u49c8kAOgwvMtPLDeWidDgPMwcn1LgGg
8NZ0jJF7FMCizwWhqRXZu+9a9oOcNG92F34wUxED+TkXYKWlofyrqmb3WzJrDTZWthLS9jHK1s4I
nOTDXo3ODw2x22BwuMfZpRWxWEjmNWufH0mo0Wd9f3+rZMqhr85tj3A+qHZVvzHPZ7I6pPLOdjxa
/O/LtmMZk87f9BbA9VpdRKCp5je/hxPlXgg2S9X1JRlgvWrF3envEQvv9+O4pDYOJn64JJVnDb0x
eHECDeX+MkJkOm14+XtqKIlo9x8YMbXBPxKExcLDL4Tu1VmBU+38UcQAAuPL7f95v6WT2ki2wTtW
x+ik3Ck+XqI+ynDT9Qr7WfHRMMKU2QrWVd5oWPb3j0KqjvzZwp+z1qosC/wvMXmhOj86eRwZSOep
G1/BdqXpjIj8ilAW+wJY6KzXtmt7aMKoHnxwNwA084fX0nw3VvWfyZcAHNU9R5ZrQAxWRIKRpPZT
zI1AMx4omSLZXWz/DBUqncF+Ny2I+31tQyfMeDEgrp2MY5jltJZsiF9dV1cgV66u9Inf1Gz2jOct
TsBvpnEvp35akwArZK1p88onECm1Nk+3nWnj9CiY8+8fyhReNQ/d+wEeKRerFKK0WICF1eNF6/cy
yu8UVLSpfJabN/v3fluceJgAS9JRbKzt7jtO4B2CKeRTeI7mZWbHpjrrcFDiu5hz2/SY9pnLCTw3
VuDU23fiKrRR+Rs7UK5KWR3rWHmtfWmFYeZgmyPH//r4ke0hDvh+Lo4yWo7vOujpyLJz87P53mmo
5IfxZkN0Zrvd2LTh5bn+HXYXVifKCb/OM6YzK4R0iYarnMGE0ZNGvRHbY0MdglPN7nVSYFX6s01k
eZHjKp+f345RkhOR9Vs8wi6kpivLZbK7+vrT9+mDS5Ab6lQqst5USXeUvzipsswDEcFDdtGe9z+v
NE0CeWGZVHRPFcHY0ekCWbvqJR9N7xD6WLwqLFddR3qznhdejOJg3eVHxK45BAFiVBJL2CfdRwqm
CofE57FspRAiX1uphiDA7g7P92iY5K2YMwTGSzcGoX0oR5dGaFbEHPYa8l8uv1bxvoJSA04BBW7V
w8xYMbE+0WmFYElUpvcnwYypT/oI4caai0zSISAi8ytdObV5jkGTXF05iWScLKZ77YkiYzug4kZZ
YrAOVsDu3BPsKRhs86rCFC1Aofw1VbOpFPn6PW5K0CY/aFYUllQO0jLnI2VMSpo49v8phremiPnN
elxDYU5MYmE+1yxH7hvP0SEiXK3eeaxiNqmBhWc1Nx8yy10hlD21zcR1SQLtEEFtcAyPUEDZCwhb
+PZzAubrCB9U45WpzKDcAV15MnY+307EGWtcsI1UfJlOHvRtDnJhWt6bkuvWKuibFaa9E+FSsIX8
oe/+4zSrsBByQATfP2anLFDyhQZsjOZc/2k+2aQzz8++rh/trLNy9LXzKUqTsxBKSIvw3rRna4G+
7nrKK+I9d1kHq0+nf5nqb/gm0BojL6Q1k0/0Mv5Z4rNO/ekiro5DJ/lQlu397IAeUYpLmLNlJCGo
82TcpS7BDzdFfxFIscIol7T/5G0xvO6sJ2p0SRG75OlZH4D/Jq6KhzG61s9sC41RpxFNywrge4m/
gqWvtRyMznjpnXy2iGGnARJxqbEnnZ10kinzYTGNWmlv2K3UsjxIjuaFKSMtdSscikEU6fezYJ5Z
82wjmuXyBDGoZ3eM2YPqQxHKnGZdkXxuNzr0NzAYeFQM6YGAOyG/8hjxTOm1pHolpEh10b+CGV1z
x4qOxHuuKXkcUsPDx/sHhNFXleN4wheZVsepUiIsgPFroT6cMcjFmbFg/921hpSe5PegmjPaRPSg
SuuGTD3ZQlIHNI8JDvTywy/owg/eSP3h+Nl28XOw8GWnNIlLxPztySrqRarv9AtEkDOHr6us5X+y
Z5HaFebvyzftSOnE8cu8+RTJ9aqsz0+eDtCA4RQOTwEuY8L122aZYLA99zGhHVTx7CqkERt/Yb2K
8+KGlmcMXTWw2iCE+4GjcOtoi+fs+ORHj8Mw5Png7XYp5os43JlWX9qLmw8XfSFzbk2/bCaFyy2A
fiqev7+Gnlkd+i9+g9NxK+4Wetss0bCWYNEqfu1NHX1HOmEwAy8Xn7HrAJB3rQIY7OiaakMxR7LD
bKhfus7wPSpzglvi+QcSLW/CVJx8Z07m8onGUTUpV2Fs+FqxF8UM5v+IES3Agr1eJj8leKns8JYj
dmoa6FW1ZZb2yUv5XkpyLBbVS17X9xXr9/jZBkhRYC3Ze3yEACE02Kiz2auPsiVIaFX6ve6+pDWu
NulmrbYqgf3mwD5kTwqAIIeYcyRnmMO3c+FaCQDEQxEGcnReicL792O5xkJX0O/enc3BYHdqfK8B
+vkQ1vdmJvgNDzG/0dD0thCTX9tcfN+P9gULdh5L1rSCNq9ZLAWYQvlrw2TPnk7ZPSF3GmmcyhBD
EoB/g+sPg9OVf9UfmhfyyeueClH1HxTg4p+W7iIF0BMBk9VTRvgzuXp6QUte/D1C0ZN+xjAMlsOE
DiGZryBPOb3d8NixiVHZOabYO6n5q/YJp6Of0mBYF2xBjz6DAGRFVBtHBdnFdVAbutB4h0zCtQNc
bmfBxfj2gDoSo3mPcKDO49H0bZY85iLe1VV5FIgUHLPmdZj90Wk0nScnCzUQGeEdkQpXvoEiD9bQ
IhN7kRmiX0843HQgwCvfe19vDSwxQHD0EKW087vaePcHIfKBcDCVdPqwLMNdXbjBZyN9SONzHtfh
olNZ0MEFudiqK4T5jDNsPzEGrCkkZAFxtFaGpa1HCZlRzd2iDEjOMojqZpV0SGZx6pqTkUUz6W2r
3qYlMc+oyH/3v562K9+0JRpl832PYt7yQNaNsSSHtZpHWpTHRNo3J04/usokmcX2xWSOBRmKbrsQ
B8NmTkXCwZz0qKgP6hINnqqQ9kH8SpwRmqPtipZT80HrYU3Lrxx8Bv0Wd7lHpAmbuOHAPSV7eWcn
kNPwDvcgm7adqMaEpwBovOS7tTfDlva3obJmqWWQNgIlfsrExG8mM+ICHhGfvDrQLpwIUqa1+mx6
dGdELyVyX3RONjI0GjjRgdRBqoCQfVsk0+sDjsevVPGtON+q+ngWgkkSsvlhfDQnyHrO8SWVxRhR
CLXMwFgDIkh+7/kolWb/VPvVEdcTG0pYnrBUtqzvdUxA7QhRduQ9BqHfqEvkOsznUkFybuO32MUp
hNBvvj8ho16wCw4QoMJGr48bsRdzD/WGH7diHF+uZ0WcXlxJI+Haiza+9bvcEvW1hbXXsqlkd89+
eMAUBHs768TE/68gDs2KFc/yidm5D2EzRsRYm3n8kaOppFu/r5vCKUDPIK1UfQEMhpoosfu1Onq+
gKHGTTSWSeeK1JwCspr5kKHjO03ieJ6AOtU7lJImormRnZGUNXUFQCbaaVBcWdXywQLlsHfdh07O
BSvcEOwsiRcIEJycTrwUFz7sHwlfhY/u7cVWdiLVZj62XBWmApAeSn/O1DeaNboMJk9IblBc3FnA
54wdkGy5KZmnm3gIH+Soa76QVUuoE3fMxMbL8rpPNiMloUbENvjb55n0+y2g5Ps/AsyJmaFIPzWt
NwQt82E7+BGIzgXNsCbYGUJZJzPpE7e35ep3PkbVoPu+BJkCxxRmiVlgZwS96d0w4iqN3Y8/TLaU
mw4IZKefFmSQw7jqzwHc0v0QZ1PHEwm2gaf4zpAHggp5tvm7K2vQDrFlexPW+8GjPK8AlFnSoxK5
T7d7wJZ5yIJtw6pX5HZ3liuYkSgu9Dnf0xadan2ZxHqaV9nSCovBwJNP42GH7gVR21TvUoY2O7qH
KAQjIUN/IE5mNstKUbtB/js2gfC7Vyr1ZJKJs7UX1r6EJBPKo6rwqVfRptyXpp5v6FEsz0V9fWOa
Srhy0ux4tHExjPMnjrt0u5zL6+S1G1eL3C65SuoHDI9k9ShJRWZooRgDUz5QE/ATOrfpWlKMJoy/
qXiLztAYh4NuwbyuIJsg/Rs7i1Jvxf47sawZpRiB1jBFRYvT1eM51kTVT3m28D6lMZOc9ERuzbhZ
kIpJ2QrqdHONIJShwsLFaq6FuSTzxqVUSwAvYGiByQ1u8LCdq65nryrgh9oR1x1Brvzs1Dynercz
MmYH+RDg0lgv0M6WzAqb02mYm/hod7JmLS0UzPbVsDFefxVdXi856ItIdoIqdn8Ql5Q9me+NQIoy
LhNSs6FkTQjFZIJglcR886VKbjq/NvjElgPTDFMZjTTHOCoa5tumXL+QL9Ozq696EM8nFi+zRxuJ
Vzpz8xRoGh4cOJ3I/vRN5dHt4Zsg6N4WsDAhLeQDaXEGREj6ti29PzK7DuLAti49tjKl1gWkgw+q
H7osGBJm0z3bhmijuR5Haaf2pIkxyvhz6uzu/pw/yNsMfKZYSrJljQ9CG7Ij25WCpn9F7ERH2/GR
6aHfA19b4AiELcGxIJ26Qp8lWhoQraV30bhJ7FIOoJHzaTTic7shgVtc/fjCoq3oLSsKgv0pCSM4
7Xv6cLWjXah54KSqpqiI2WMW+jiiRas47Poz1KYWHR6pBlODx6V/+cpt4uoEbNTqV4qruW8uB70z
5Wu9gpZ5MeovL861xTLNzZjITvgM6EhWy/2GMNOx2lwa2WqOd5kxsocuzKYNwD1x7bh8md1VD2y4
QlfweQSLhq0HSb693gEz5CCJi1w7o+KjsGVFUK3Us9WBSeerWPsHcwiGbfjoIP5qp3THpj9xMMwy
kt+Yrueoal2s/i7QbpsVaDqkhMOIhoAXAijtwqeGF1txlr2DJTVH2PTCO0MvT29wQnTpzYY1wNcV
g5bNMbdvN6fcwfMZfZOgPGqG85DYSrZPGT3JAr0iQ1eIXsK2GFUlH8w3KDlY5XHtlcJci7iIYSj5
j9wSzbwFbM5cgAg0HudrJf09ix7rXF2GJtnjDwdQTmLco4F6BU7uiNbtuWxfiC7Z9JLA4Hu6cjey
thLaw8MCLlUw9uc45xMwLrli1Aa7+tkMHvzxJBYd9Fw3lUF3381RhE3w8HOWa4uJ8cbv7TSoWGaQ
wTEhmJaO/3r02tVl6oEWFLO6ddg3gDBzwh6lUNF5i5n5YJfw+BGMrSRNGpFehjbJOMi0xs3+4NP1
BV8n5k/PowUNa7+vm6BSdkaH2iebQO5o4C5oKTP16Y3M/JkBOFUMQeT9W5RUb4vmFsgwWh3Ji8i6
dSpwyp9dNaP0+Z2G1T7bN1jlqBh4DKkhBpe9U3PZSmoInwwVWRLSx+5d2R/QkPodjYzem2dMP41T
32f2Ot/dUnbQdKdJXGCOCVRyMVJL4/EKM2o6DKOf67t8VxlVSk5Vy1BxatdqwWHGiNKoPUtxws7g
vwbkidV5BEqVmAf45Fj2Nm2R5zlhQPzARmEPWnCZ51w3xSdIgN0N87/niCBVMtsKvetZUSIoCwuh
SdXs06q1RLGBf5fLw1aXeiG7fir6MLv2Dm0sP7joGQJeska0KbF437lbyTm1xzkeflgiejTO4aP5
it815rL9CUSZJkI+HEKQGftRyOBwk74WGRY7sZ4qzlu+mnRPcBSBy5repGfiHbUr1qOd/lxc89mQ
axmY3f0ovJXoso1GLNzZKmIF0C9Q9XYEuWYtEAGJLk/R6JhCqH2UnmTkaNWl6WjQqJwBZ/LsqoOC
1bT4k0R9JsxN464uHXUOzGnUFcUwqCEcFWnTKJ0iPiVZ8i0k1L4FDjoRSWnsBPdTw9JsclJKU5f6
+wzmi0xJltmaMMjgPI8Gut2CYvB+q+06Rfso/iBqjfIa5KsJdSRAanuqFdOjHTYJbGwH+NpjpsIa
JqAs18It27y67LqGiU4xb+HCIsueh90WtOyPD3/JUrO1nbUlb78DVAbeumKO0Kur1GhscGy4y403
ihYZjDQHQiUO+PeVAo43e6UgqHYoZi9JymKD+N6QGTbRwhF7/YGkJUKV5gc++zbyaUX6LibWyvXg
IBIJdsnFmQMleVzkIP6J7WrLZj9mGfg+DgDS8rGequugSrzE2nBz6aNpRtN/U0HFj5IIOaR2+qYm
FiX4md5k/9Jie9Jw2SQ80so5y7lunlhzt/mK6F2BaFwCPWrtEM5lkdlDP3iVaI0UzU0VTJYKA9+S
stNReGfb0lv2mBJPOvuxNo8JF+RICNg6MEfv1WjvLYRy8hmMlbLEc8WqgMm/eoF5x85JWmnaig/1
J16ChnzjiX1nuGov7I/T1T/BI+2+vcE2i8oInRk94AlP4hqTVcQ1ZAnF6wjLRD3prbgHl9oiB+bQ
6eGlM6GX1fTkgIwpZ+Cx9sYw064y9SfEpwjTzaoLUFAz+YYSIk/mQKseyfo3a0Ey+K+9HYjwZiDs
mpEZPeFuKAW/vXHwJAX25MkQp+DzIAj+W+E1DxZZiy9Gi4u/VXizBi7usg5Whbi+BO610w9sCnUw
xp0pDP8SM0M0s4SBJzBNWTn3GCOa7FKDq57jffAHfJrACHzLEjTlG7aI9OCsuD4/2ZkSxhBN67EP
Tpy+/D3CkIprhsQIaS+cH0mFxKAjpdXk99Qbq/RQbs91L5e/HZG9kMNFqlutNL3J5iX/KQY3n6NH
j2t2zyKr5CipU1VcJOFrZwsn4jC5r+a8nzpzWOXyPd0Or//NawjLC8Dc9x/pbzUqRbm02lkzfGqU
6j3pisGUQH4+mXXtRpHcxH/50zFAtoiy/8SzHB3p2eARmEcg6jPBweVDuQFWx4G44AN+fS1nRGtQ
N3J9roYBY8od1zyTbLrYs8dU4L9XUo7z6Phd6ull0QZ1HwAPD2M9mdit6CyDx9j4UIaQ52dUEPrq
nDlO8UcNxoXuMsxjb23RVPsEADbZYrFJ5mAfEVGK1GE+PUgXn2+ANV0haW/3bR4Go43cx8dRNml1
6M3Sk4FdKtclxvdy8ISf4LXk8fK+QhYoNVCVe0lpWjdT07jO0LynqlLJGMdoIXzTUT+M+Rxh9axc
3yE8qUviTmTz4UAPQ+MIg4sYO61IZ19og9LGPWi9jCJSnQ3VCZCJZi3CGo5GI4Zp3avZcfNAa/fA
62O1ZNxCvyxTuLvn47F5LktIW9k4Kp8bju7KLcmT76pILK6CXaUJLZdP9joO9+6A8O+JdAzds80G
KRWYUD4BjTknv+FJK5LzqqwMQrl7HTeiZPtzsiI74do+9uj/fy2RCFB0kxDCcXnGQXaZ2w3rLZr1
9FPxVziyx4IdIqWzwqXuQSMJUeVEJSfthZQfLqTaCsH2YW9vLJgEQ7QioHBaap+N1D10qvhk0ZBl
req1kX49v3w4mgRft8wwOAidxTXY0cFfSJRWrXGzd6pVbajsIynyIfLYupZ9BYGx2XjcriGgLpzv
5+TddKUy6zFDL5yCS3NPVU1L8onkM6Xq62iN/NVDDJv1JJAzbYAFLuWxwm/ZVEQk5lGyK8cb3dcr
Dg4UAvYY+PjnEPpYMU5BS8enc/7DbtiK/Ydoj/XlAzRMxZHt55oaDRiTrpq9ckKRUuXta8KoZBcU
GvoaF4vnc9A/5jRY7zQ+XPZmBcNUIILY2KLCyhkik1zaiEqKx8eGj+xiLD/pQdj2GLUW4HwoRMzi
PBldX2jVELjWg2iOghvY0dcnEhJDVTVd44kng0Z6u3iVoBtqATFc91/tEWkGHIFtGQsrGpP1j/HT
hMQ415M6EXz9/A3LgNAB95h+OuO4d2Sbj+o5jLc2Tf5b++96JI5gsMmTQXalG8ZE8rOLZg/3TJHb
BPS6WLo+ZN25KHCH4cKBAZ+c5VJ9On0d3CKCwi0xhLBTZzfaMlYS/iohjEXaQoGVGfykVPJiATkV
ByjoOoOPb3l0HyBD0Ro+xp89DNfYMiXiV+XFdkIIsaosSlUFm2A7VyRy07W3C1oKZ9u0F/L/we2F
17wrVYTBCkEpX+Q+UaXaohBq9Vlm0fgyB2pR/Wa8OuGcW6VEnZD3jT5Bgk9pUS01jI4+ODyLFvFC
Dzf9R8quKqRrUiuimsP3r44R+urDXDa1ddA5FdEu8vtM3Pj/ppLcnku8DhjG3XR1lVL+79KZROgr
cSkHfeDgxfSPk99a6RN8bTkJcDrVtQUU/vLMidQ4LC0oJBy3PrQwREA4tpknUa+wG55eOmYCREOf
Z4QyO4v69B+fvlHCs0hqv9w7gLc65JGf/R2Sew2Wzyp5iLQgCgo2W65eAZCpegYy1QQGA+X9npru
vSw03iOCsyhg/W70sV7DECVgxx6Ic8I9FLGAo6CRVQIk/3RWOmSIgKshn5IJFRX7R7pzbr6xgZdv
Unqj9I+c77IMaTDvx0b+fgXhYG6MqT/64jLGdJbq36/1K0bKt7KAKcu2tvrkP+MYi1WIsybLMEjv
c0fbynD67lY5WeX/0ipoCZdSMtVnU40QGotl2bwq1m1lxt4G2AU8u3FRY+qorOYkLrgGXg2+66MG
wyMtDL6mq/GYTDYKmiN/MiGpSTueiQ1pBbMdlD+Hufb5dgULjEQwkg7NG6RDMBA+HWjqQHyYDwnV
a80oFMbadYtE8TUi8OldFzwilll5TmcUeqhYM80kgNKJI8IKZ1ZEsUH1KDt4CBgUzZQJzdtoVzdL
uDnzDZe28Zj7q+RSe9x49lZpUqFAcrrjuDxdwz1p8EBJyxG25pqKR8uYLQQS2nJprUlYiSwwqDFt
ZAyQDgQg2VcHUgAaFsjwTOFP9FsGvK+nUvyLroiSjXQdc2qYNoJ65cfZ9lSB0h79oah1Ah25rdpD
afCgow3xol8Nr3FsGQWDLaF4L0AFl0UplgT0i+qN+OlLmb2GoLP1IDWh3COywemDsOWq6G4g92C0
TeJx/MpzgZ1on4fkI4ih+Qhq6nVVStpMnU0o4jSjpZ7FWiIRWMvuT18gAvTr5L3YAeWgtnw0qDvH
DORkM4Xj8Bolh8vOipGst+nlroE84AFGeBxSqWzPiBa4y4mFgM0mTO7xng2zktNohIcQUiCQ9WFL
fXKjzFwC6DX0L/NkaFODkvopX0Lrh0Pt8uP0VWcBFa1LQtyZDnt2l7beZH8C4kVH2z2legEmVaQH
pLsnt7XUboSLs6V/rTojhExB7CyL3gJxOzfQovCcCVDM1lxGqa1PiaG46VFJHVd4m+Z0x1JVdvok
0L+sV0xEmTvPCXlgrh5zxkTvpvJ8niL2PmMwUXVUDv+OTB/uj6uipQXtwJc3YSKQPiWAlRn4fwsT
4wulYLqaWLhXg7GWfF+F2G84yiuA0xjXonLX60KQsMjtrUVXlKYAJKOq4I7icm2TMHLWt8u9c8IP
4mX1pqRiRNzjN5+TGy5LfnjmgutBI8UYaD2VCbX9i2io7jliwN7SfyQhf9uZaBSapmKw6NSUCYqD
guzngt7uzXwxqA4oAVJ7VU/TkZTYmET/O5rmYUz9y/X6bNLEguJ0uXyWES8gOhJ8gnaHy7MFK/C5
n0wGP5W0T+rDMpV8uPlFzezmmlETo4u70PLK8R2GJnzH8dqV1HFCFQXWdVVD6YzTur+E2evQfFEQ
IkWPOP1sWCYjaF8oy2tZtIc6utq9tclqIQoLMLszFJ5h2RtvzVidg9V/NxZOQd+Botaip82tp4/y
JGxBsA1iKZqcL1VavWbnltvUj0sHEsyvjWTjSNhpMIF+H5ugwtlpVvALtan45yZ7KUNZ2n7WfMLK
GYJWdkM3xldXE5fiqpZwSZaMpHyeCd8i20bvFNNYJwfnNNtly8d0xWRNiS6dLzH00tg7v+z3Dkoh
NQQqlSt7VA0kUYSPCuog8cKf5lhTKDnyL37BM4kx6v3yuL232MVp/m/nNyvWXkb1y8SwVHb9CkoE
nR5q/wOuX+yUV67dJlIE5g8EsPjGCkwsDiDuxtLbsRxV7O91asHEOG+gw95FcUkqwbGUD6Ja9KTp
dPDlfZgdWIboXxgAD9dvTEF6Q/U1qDzN4p3ZFDsJA6HMZ5kvFEvKgMjh3fkV1Y/JJiEwA09sSLol
AI21vMLM/+o1tQoW0FkgF1Ia45zYjvc0f3k2SfNHtjox5/ihMRmsiCb6/WQrnXbJmjNVhNWPQoXx
CM7ej7QcLaoTONrgOxEmXAbK9h27XQ8MIcF4PLAPQhoQ87eKCquRE+2cEVRYWYGCqr40d6x9j33G
MGaKByHat3LZLH0iEJEEp1W3EvIrVS2Lx786Iprs2JL69wkoMmbu1UXOVo6uurah7QNKb5TiUD2h
a957kk23TpYouoVRJpSSraHWivwmxtKiIjFhfzTOEde5HEtZL/IuIflNbrcYA3AsysP6/kegooMc
OR5miUBKDXPs8NWD2VtjpALQDBSKFMdM+eWfGnaQI8SsrS4ArZ8PvwpHS5mqxFtA6I60UTr5KlkC
kDPOzmosIWlCAtyoUYAGFxn4mFsRGVkAj9Jz/rJYN3o0ZTo4iFQc9OIUqaIvmSbVV55KgybDI3YO
HWAHgxi5mw5srmaeVxFMPTAs7A7PdczhFHo5VFAngqH9xV7BQ3QqyojZ1L/qXdIH660kZ1bfIiDS
Do3tBFzKmbmoWoDtD1mpNIc8WfKwDl7bM3Ru/XRIEVbJ4ucMbYu9usmOG+XmCVrEy5P6/NFKf1mX
7MNIDEXX++aSEjzxM+PHUjsqd96SLI2US7SNMrlfoPkF0XhxQgSRiihEsO8RToWVivKaD/BF0+JD
tfuvSPRaH3i3SVCCxGDrHXEydQ23GRp6kXHqgrku82zrG6vQ9dUoS9BZqYXTA51oUczYBu9uZySh
jr6AXyRjO4nQSPILuYpmvQHLEQTRnjnOz4pP6vyfyHmqUuJnXoR4X3LW1AWWPHaORpO6MGyj0G55
gCburmjGwhZJpZUGStKdsEAKdI+zoKrVf6wggdRznz0R2CBkec1DCSVNa/mzpTIsmhJSPhNggEe9
3+Lp0arAvxXapvnNCIg/1xmVq8o8z4YyY6ZxEjkz6I/KpD9WwXkOImEYN319mJE6sZ/1dpwnxJlF
dImt9gcjuOawCuyBkiZxFyCdBqk2cAMQmHYcae702maIUjSTrtQL95Lk5gqxr9HFAHBPxYiFeCX3
DT0zVpmlE1tbaLIr5tJ7tD+cMqNBXv2dhAF1hiYT2msyMklv8QtsK+bE+YVaGSS77ETyigq5g68V
ay8NvkXxoEFCc5t5RUSAb7aCZ34U446tG1bNepZhiWIEPwuQJbzZDkbHuqFxgY+CS0XHMulFGWTZ
Qs1AKTVk+vVB11Y9UVxjUUXHGpHggxd3vIBRX/kLXA9BS2MlLLAU6Hz0QsWVl5FGXNufhdRAFMgW
ZlRSdBjv4cuVWtrPC8cTi3EBmyVWaU1KKAeRnnNB5hUv6O47nH2HPLQQ2u77Fj2l0jhmp12wrOEX
I/3ELzDNYCCqunRiUu3/LcnYTMUUeASkPZu4XnONHdC/3xGBdtII0mMFA/JM8SH63P05aNck08/G
mg/i3cFM/2JH2wD2/VCAwxxQjkrzgC5xyTgKl30M0cpTuhMxjqddfWTFo6WscxAzGmyzyaGMke1c
s3iuLUuSI6SHmbZ9oFOUyJb3rKTmperqY/rZEjY3C/frR3hYueBDLL+VdA91dWaAfoD1nqsqZ3Wf
QRE2sQWAD1PaEGJ4oDI7d+tfd1ZJHSRngKYNQaQCUGosxczCP0kw/jGVfZBUzV+kspxWQQscWtzJ
08G54sywKERu3F0ibJ6uFIO4qVrWqscXWwnd5HWz49FXxk95aupKClUwzL0yhtmWDrseS0NPtDA+
kHgxsgEWCJfILceMKyCgE5UEonoKOObOtJhDrIAVL+bQ0KTchRj7MqREUXt1hd3Jc+rm8SXlciyu
hPxFa5vAysQEdDUyf4f9Lt01ZSIZV7OeWdh+URUrncJmdAUcefFql1fwySXPru0Qkkqzbm/s/8fq
SwAHPVe3bbHvL6ND+QoG0XimsoxRrhgRv1FxVdUSStN/2+5qcl208ttImddGJYl/H5q6SVr8fzjh
rRREU9ZlHCuyfd3RuS/bPKIbHu1BBXKdPXGDTC7B8mKISyIvNZck78oMWMxtxzLGZuPP6c8T5/JE
FMmdRviDaYLPnvUq+9lVcPgUlHhKYbvHkD6eKl4AWtTALAL76kmtF7QqyPBpQ9Ur9Xeii03Bn+4E
mTJyHlDu/8rblokf58hlzXJTBmplxZtH1g8CGCXhObGAad21ZLx2wvmbjH979Ew2PaiXTeIjy+AB
jHWNPkTKof7eQEMRg0sBP40XjHsjyHFAjP5KBLThnY86TXERW9HlWSN9/n/QvK0S4zsjBx41xyVj
3+sucwpgMJIpviKAwqVvJPlJhlo3opk4+uHvjc6U+ouueCTo4NQiTRHXPNBlQvnP9PNoqcJNmNIz
q/wiJiO/3unvv4PuC9AYsCqSNHOY0zBz4XdZluUvvEBcJQ7zJty/UdXLupb40UkenbgaS6sy9JGI
GcZaiEsdPLR1fC01Vc+oU2w6m4D9dv8bbUujvYjBNBTRohKV1O8QJv97nHLT4aJC5QknSoL0Cnjv
t1IAgf4gcVXRnHM5KRJdKBt09x5uDYJzc8Yv4lgnRU2shWehVSZ8E9iPNzjlFjnz9riuH7QKXg7z
f2GGrqKYSMG57nLjXQ6yEvO1+pP2ICviNtQ1fmOyruS2vSMHnMKQlB/QOvDIxHX0bylyH1ihF07D
M1d34LH9yfIYUPxIQsJcQ7tyIXdJH7m5jJo5YdVSQLy0hOI4MxW+gpgKoQjvfnxkl9j18Nsmz4Tc
vELqWuQMBPiOWfRG2FrskZpRWjA7jzIRPeAEDjv2q6PN4NJ1qeyUwR07jB030WRmNgJ63gy2ES24
pRtp5MR0QLFOd+BWHI24j61o6ZmlzPz68tFwZOlgqSXw1H/ogJIuhmnDrka3UwO50Lz8S/y0P6Qk
YbwVzWEIYcskB8b6CxrMyncaxVkxd5dAvOtxKxuxjxdmoPdsCWPQi6ZD69Z/2Wbhkm51unCsvwaG
tBSeT1zTlea8CUglQ5JLLKUFxUdmfEJMg1iicW81zwicARmkf2/Fy+LLzgyJ3IxzcIeWNufUs0gf
iBHf7V/cJt6QpGgd0TXVxi3POXMPW+VgB4s1voKtU7AT4ALzqAtfxORQch7fmn9NpCruZMQkuMa0
LbZYMm8fNkC4H4TEhlc5BNURvWrZx6hlhkiWVy7Aczsy9A2a03RI0E7fAjsRvBwzvW4IHM7+Aq2J
ptJ1GdqC+hO+KkDugrJ1vsa/yTLlyMBAfUPADszQ3oWcOLM9QmX6ulzTlpFMCNEM21RmeU8rtbKD
lX5DbJIFmWlPzih/crPHkKcKZN8rg0HkEyIkKdJ6SJ81QjPdfjaXZnZIDp1lAoS0wcczyMesWPVo
6gj243RQ9WsL6kmGhITIZGpwyHvNXvaXgb+vE6OvP7h5xnCV/EZndbVUoI/lf0f3yILJhP9X14HA
e9tbO9yrLWu2Ny2klYcpXgwiDFU6tkO+KC3RqV9damDeUp6odQ5q4HHr+0h9bxoK2IrQZulzGNLK
qxmugljH1cUSp6JUdqcguOgm6XgxFAYnpZsXKExmdmcOK5j3FzoZckX/u2w6HItcAHBEU8sU+f4F
RUsV9guJkKnXbfd6xc7jVQCmTHT/LqtTkwVMOi5Y+LljiF4tlWTEhuz/vwD5zllDHrD8uarAaoh5
sLg+Jxw75dT34hDWH2RXO4OxlQTVgeEjBPR+fgmJpvitTzudxcOAfwZPHJ9tEaBbLQ9ByEKVxAeZ
8+haPfHNqcP/zFXXsUMzwumJZDa3c3z0q+F7uWzbVah51urz2XN4V3KFgHC+NH40yjtSWoxUOT68
tpdaE4bZVvn7OMrpMOwMgjC17iSN/1J03HjN9f5wp0Haa5hqnAdhjHNfC62uizHHKG9X3dVYI0AD
DIO8oTqOlvks+qFwb2bbqXY4wkdKiRmFMWdU/WjUliN1QRYzOqGePSTKtIT3f8Za4TWSGesg1AEY
rBl95LQ1R7TnYQPOYZaasLqNnRx1P9QIgsKqfa7lq6R6begD6Ojx5V4gLLIuzmjmR9nyr07owv2B
nw9/JiwQsQi+PeByJ0+2tCY/s4Vkm0Ko/Fo7hbCD66sTOBvsiigmAKrtIeaA12MOjtfwEkwfx0f+
1Xwx3swRXKoHZmAAjtCgcJ+QWcYoCne14+2jTEoqa3EEebOfejwzNgQOouLiih0MEztOICrsGlbs
5P3oJX8zCTyOQe6wnbLBLIQ5TR8l3+e3a5HU9mV/gm3wPPziO9rGnc7S6oXKGJLxk/avtqDvzyoY
I/Nbi4lpTym336hp5v+/2ZPxEymQcPJsjEgrA/HBIVbMlNE8Y6XkNXO/KSRjGfqWvchVhbAFll9K
zg7EcQgjVu3UBr/5W6UreOlADC25vc5k9xjTOGz7MwyxOHGQ2z9EAu0Ha4aoBOFJ6V+KmMqNow4w
JcchzIs1g2KsQcRg+8BZq8QJKzO6hVk2jUCkEDum/6ZjDkTix2MOkBw2jzUPHHOY//2Bju3JBzkG
pCxg4kAK/ND6Y7oJfTo4WKwfxfvxzt/Zx94Twv2cz85rig790JDULDfDqCpcqK4ndnzKxb0sHoPD
vdVsc3QPqyhjRDxQjwk5N1a/j1HkfBoqxzb4tW8qF0o7AtyXdwIEO4p2V+G+vr2n9EsOQvkrBLk0
lCW0WajB5RBriD4Xdoc1EQyWKRV7A4yH2hIole5Rrr+GhkChd9GX7Xi9pYTfbe7AEtq7hgVW6UbX
4z/lguwkw5q7yeA5Ksi97R+qHxlI+4fpoIFF7RxX4RKXBnNeEa/AOWcXmqemdhTCrYorEXc6j1Op
N5Q4VoIhAju0wSkdZDzNjx25KSme/SCnn7ph+B20twFG8I8K/mBh1PFtof4sm6emZAnxufeihUrg
+2rgIhnNzzD2BFslA8lt1m0tmdJhM6ShEFF+/xYwo45iEm7idT2NxD3Z9pVPOJhuzuLKtq1WQRFF
7qFAb82UExUNnakotyjtZIXjVsc5kQEHyICHl+jAJjSuXTZNf7p6ZewMe1kWzb3eFQ10TMiPTSio
oc8FI/woxOK+QO1obJtYA1CpzEZLxCKVsRXlVqfDTLj2WDEJ5lPF3YhrwfXdL4Mw0/Om+UWzdAOc
HVYFTj/W8+TTosUQOKCbJITV/MyyL/AqRF35vNaCVUo2aEcbZFKcJWIBpXwIW57Ih9uNqZ2mMh0Y
LX+wISPpfrajfj7g5bbb5UfNZ0AC1PmvYJYOs16zbrKAqQA/1ny/gQ2rg/RzZ1wxC84v6nFd0uy9
O3PG3aPXldKnhseNm06SBInRpCtLtU9c4eQqACBCvOFMcajCxAVraYYISZ910nKiM50twg0qTgZj
joaonFOZLZrLTSX/ktQoxpi7dnvuyvrGdmLvlomNyB5vKvABDtdT/r9MO1IU/bHX3XQZF9EW9B47
3fvt+jrkhIj5VOTv/queGfUsg8tQa4nuRTgYlqWckihRz6p6Ot/paeJ1dFhzuO6dKWFPY3L+d4J8
ewTWB55fGETzYZoGNSUcbqlQXXjip28HgEDqsNpd7L5yiowuEhuc7qbsKsoaJuyGtgZU4bcJ/EoB
tLEaRIGwHXXKI+Dj0OkpAPNvTMiYUTiG/d6mzyv/pPJGlOsAJP0V4Y8XKD/jpzF2RLWZ2l3e/yfj
xt/bQoO67oApQVBfaw83bA5Hz9xs8VaaUwbDAnKY27T7kWVZUSFgT/93J4DufPS9RaPzAuS84Zer
VmM3RFCU64//5UvhzH9I/DKnYxF+IwLXRGf399jvAg/IwvlmXxDeFA3MPxp0PH3C0IsdyAsfq/x8
dt+HlACqslYbyKe44SZBlUtuyzGQ15ELNI1OmB5V2dLH5zCK54cb1x45Jh1rxzhAr8BaB5eiOECh
uxT8YwIqiwWekXTynw5uPng+ez3ebaBTdUAfmfRIZxVD/u+AQCUfFdh5QDkeWEmkujr3kCDb9Ndk
/zs88+OAPLoG7e603qfZmHLauYBoFiJvdV3+qyBQCewh2QMDADLx16sGV0uvY7ZkK/5PYuK1I0EG
zcv3UR4Glo282Kz7QXxFgkcn7W8Ykjvq44wPlufUbj4Uh6jQzn83hk7h66bUQMOIWyzWr3wh5CX2
lkMePH++qiVi4quqboLp6r0pER2+qeuy+6aafVBZ+vhTetrFRf8zZrhUcmcE5dmc84oZ3UfERHtM
JRAq/PtdlV/UVxPGJURudU1rpOSCd22jErJLjGaQadJL2DZ2NgNjhLHo0wjWJDsCe6bIOGGL/Nko
lFJ0g9aZsjWKfImMu8DhxFPQKEsQy1nP6MLh1P3soKdzjJNhxLhrsKbg3msODRItnEG89RXl9S8b
OENg8ZrOA1aAjwFzPAqu96Jb9svwi7hQrTcrGjIFrcjqLKN9Tm8leHwSFXsb5OSm40Z4sedMQVvf
4TR7RsbeoS6qHCLYnPCEzq/q/b44nlxru/i+285pCaMSAdhG0Ild3/jm2ED8hAFqBCTWYQGCdqWy
PgepGq8hsTg1/pS+4ygv+E3u3ayApRjSD1kQTHCtEoofuSIV2myjIuN6qunaZA24Km1BUh74cotO
zXU8OCL/Kj0iic4IrCdxBrLQFV9HA7YlkKSQMkgE9WdEEbxhmoyL4W9Izo8q/e0PVwQZtV5XGpuC
ecMhC+NAci8zMmIQvW4yOemdLeWVsfuCkC8nIX+PjyT8OTItAtyAOpMeU2tKVV26cVnsuJnP/g8O
THxHzb8D+Eqz6sLYlMQzfsVrteM1eulvol2Wv2lZm/0Gc8tyCXFTX8yKVgQHNMK3eIeoizizacub
0yxbkIFb/xwKHut1tU4+vL2QtgBuM7GTdqS+MG6QuyhyDMl2u1SEYZRHQPyh4jNHDcOZQNHfSJC1
opfYHuSZ7LAnJdndQLNl58NNREQ0WR3u94hJR94kE1tfZ2ab1IxB5BEOapEbd+puM9ZDXRam3/0y
ceJ10D+6DdHOLXGe324ZWQ3Qeb/Pqu0/pRULsGNvYuvlXwlUQEibsznUFioPBajPuLU1htvc1GA8
dZGYmxJqoMmYTkpLPZYe9jmacuYMofRPaJ/+rgwowBuUHARR+2dGoj0DyfMWhkLYOQMV/l/1ieE1
ss5FjIiANFtQ5fYhqTBxxE2B83SUEYxYcUjblsYgvu4wl1W/XtCcXBzUPcLIrmpYKo7cyRjR2FRX
MP8/GOGWaH54KsEuMN2nkftDXxyEUZMIKnWRb+TxzbxtdwhU2fTAThYR9GU48z0KDKjDVnO8OGRF
tu85k647UIMRVbl7QNgC6oOldp8vn8qUPR2jWp88Vhvg0ZLM0MDZKbhbzNO4Sakiq5cn9478mB6O
efryT27gx1qOPcI1AEeLRwipVmSPihZuz4AYKNDHoIjf5VNXhmr9r6JIYi6nE7WrdAYVkCYt2t8B
/6LLh+4Qy/lUemAuY6fyTv6Ntc2cLPfFTK0W6hxlHqzg6BPUJnJMnYx6Ap4jVY6tcZRSI7wDfjhL
Ca232ORvivTbvwEYLtzcMBhtHPOFibO+wzUAqzUNwxI3larazDrf+Q2y4bFhv2dww9GzyKpCXG2h
bbrDBsuuiZYxfpaGA2UPmQ35Hmb/pZ7dHCG2VpIsDvv2K/1vMs4A+xcub/aovY4bq3cc3KLIpRZL
V3bqRYL6AUh6jzzhu9XGgkBG1t2vqehi0TMus2CUmlTNoUThn1tsnSD3Mup+ovInyWMwk/YhnlgH
E5PcD6fxEkktUfnn9IFZIgCWFiDHJJ+0iGMa0ClL7fx0HrZEL4tX4MmbV6txPYy+5dsDFj7GxVPJ
q1N0iRt/yTQY4IB7yhinZddyPMLz/hnOt1YO7FtzZ/RMNelM+kvY07CEjsi9KCP3yd3b3A9CmFlt
stYp9EiMlw+cd001yxGcn6n9rv1o2m1cNUbzi2wiyl4JAYENqmpIS6ovI3x2xoBBueesZDxHqYnr
e2nw2qFMZLgH2+izPbazf7ZKyyZtnCMioUZKmRWVruShJbUSX1sWgmvTDRu9set3XxlLa7w4VzxC
dZjzAa3XNB0E6cxHAANjblPpFIXUZ/xYzV8bu7dmehmNfi+ClyI52GBpLGt8IFL3QXdR3oAU995g
4m0cewBBkT+w17jKyTEVyvvFRaCJcA76uE8DvHU/wD8Ho17AoGNn4GuSXiqrlxYNG14Uy+F4a9ed
xgJXQZnzT2UW47rLvc3KTMb9aUcpQBqwYt3KRy5R8PHvs9E3uk4QAzbtuAjNVcYC2FMZyOVDaJ5j
vQKbOIh9+cnvZxc+ZCagGRHs0qJsvapumJpVD2DuRk5cAu3jzkbt7pj7wDFUTPmXSlZUVVuIFwOX
3eW/+H1DmJxoQelRHoWm1AbDuw0/pQCFvD/3ZLyaxTzHBoEYaMwswmcDcz7G/EfoXMMl91l2v4ne
yM0P2w0D1khIkSDumVwqVn9oNhDEjHJ6eZScS/ym66cpfi39UkeOqz8NZS8q9J9W+XbcCdG6XFbs
FmgyLcP/mRw/BeCNVkvbnxupjXS8wRAJddqGRWPa93SBGYup4AYALFv+Zv8DKLV8CfLRoWdMqwqQ
4ZCoP3DsEVZTZuJ8q6nYPCUIfGvCNFldGznTMgywWwHoWMWGJEFPU8XRgyTJ9Ty/gC/H7EKFKNwh
4D9xiVvkLqvFwsrE7OlPbC8T9grrieaElMTvraSUrGhN8Z8+4qqbLtKEHFlRHLABlLd1r+nlQITa
fQY6Ymn742G16OREroZWHq2MepLuc/LiCWT/r1AwipIBNgzW1IuJNnNmxSbRpfKVGQT/r9a3W0JW
4/2TuZ8ywXubyPCUU/a0wGi2h+szWrl5otmUVVnE8cjFRyDUvKimeqXry5Hckhq26pWILHwFleUe
BkFPMWdEplzewqRDrx9n6rWLfLc9m5d3/OwwgVJwXUTlxH1gqJVx1XckvcBhCtppN5DqKK1+qNIc
A6KQo6ieXn3ZvWbm4HVIZgjjnYW9hbjBCSaYZV9An+RbSP5B79qxrP3JJq3DHLggSTjaDaZSuQo+
DZvyowS5f8KfRPKrxSm3P5EMhyzTrtZRPkg3ih4I/nAJDuiZGVXNKU/mCak/dqF1X+TvyuS/t5Yf
TsmcSRlUwoQqT2P+ngRcL7qaHbdJ+ZZABxTAIqel1JZ7v2raD3U3r9vv1sZyk+X2XDzB7pCgFK6v
LSJDBN2lWD2/vEk4BIwaphRzvQVDo500SaSgliYDY3jO2cO5R1EDr3hYjFBC45mY+a00EwTFuNHP
hoXU+L75lBxAZdEExggxLo03jGYYO9Ri/kwr7zHzDsh2z8BQgd7KUNL6JTEc8E5gszcDsuoRIZ5j
yMUuV9x3kAPR5JPjKj7LMFnrU0pMd42SFGcHlY01K2zhkAinWsjZf2UfCzqSSuZVDVJtzyFeOzce
Gwq35cGJ7XurkRdx5h7T9MotSQgMRKRRgFRs9PASaBSWot1Yo+XNWeRhtN55iG6uPm21wQvuptRL
3/ztW9SpLz136cuUIuy2xy6oBWI8VbcKZSCERpR92+u0BIi+dQDR62c6tEiT2QdI/X8YucUArh8B
NM2lRFkcNMD6ve/htTmNGlPEJRwiKk78zoMsAlUGS+nbJGhtty6+dD6oEOxTnk+s/p2T6LzY7iNJ
4wAbOSyp0ElARDuthxjSVIx2U0DOxNIVcY4uhrTW70NeRhvWrglLM4KJO2a6Y4upSH86f2KuLTa0
ygTN0Rp+fR3A9U+mPng/o31qKP7s36OgRKpPq4P+eKL3NqGXWcaGRgTA6uOEvjEnXxH7hIZVOXhI
BTIlDzTRU6yokOBfL90uL5h/5IQS/Eu5UyTWb9HaZZfSUxUe6vxIt23aLHIFIOZ2OTLvXxI489fY
fYkvF2/Mju6gzCaFgM8a8ZlW2jMgMd42QrXswSt6EG8PkbvkIfouR8qDP/7fhjdisRupLwlqWPma
sSkNyC+rZkGlSw4bL+iq9FjgxeW7rAuZPVhbhth+IR1iO58v/8SqvQBo1oJGjKt93bfSIKW0/+WC
AQBcjoVRqWc2CueEz8uOXqQjUuTvNEj8xf/beLoQ/dJR3rBR8igltL2tEb71Re3BFKVRSYndLE2I
u1XLf5Q3armlzn/F+IJY6NXzvep6qDQlLW3o2lMNlYMNErXqVKyXdxyuNQndrnQoGDYBXIuxXHan
Qw3NCSV42/tSrchB/opfAZN6AKGK4p7OVydPqZFN6roxe5N3gp7U38rojUqLFS0rSC9IUQBygdeR
J8fsm2G++p/7g0rguD4inng2smOdSpUHC+Qju/F1dKvdWypHLdVQub2T9JWb5yZHTNfLci5QT9dF
bqxJ+c35IawEWxXGsByj8lSsf8D1aUHFyu9dcgmZxMzcBfHBBw7+rNS0eMxVu1gQqXTHJIbSyHjL
lQ0Jcti3hl7Fb+2jkBWJpJMxwamgZpwYOis3vQ7hJOXeR23pOEHEE5WiFUeNoiosTqrUcskMWw/1
IlMG8yTEQ0swssTQ3sE3tLD+NscincGnmkaKr1Zr5fnDJzAPv1YpsufjGXd4YlOFed7ZenWEiAlv
2voki5Rm3UFK7ea/bFBjc5WpyW2bcs90RqD+H8Oqtn7grk2acDifCmrdMm27M3KzLk0x32g6jw9j
M2Xm3DqdddKdN1HRBgxn+JlrpDN8XH1stdUv4kbfk9bXu0LOlSSaHgs5sD9xNxpD3yW1ZvzbaOsK
6YJ2chfOfWMcMWSLLgG7wc3qraRAOGIKz/EqPuPbfIwBnn84aV1MfiO28ulG7ui4PuzWyIIvUxmH
eG4ICOpcxX0alS2enlK81M89/KshhEnYKHKt3/xcHY7d/chl3Cgn4h+8Rk2BJmDr7hGI1It9OzKf
+awXI71xirrsBYEjERFGIkAkE1AypE/cpKrGTMsg0rrzWQH8ZLqr29DN7ImWoIWoHmb35qLlNKbU
/xiE/D2SzftvpztxgaUacmob85GLw50cZIoCM4xdKQVoslaBBGPBWuj8irIkLeWoPH5miupfNe9F
pfUSYHAc4lDoff2FS8HrPcXHlbsc2SAWHz2rPP6Yc+Zwu1hBLBW2EIjWxtT1brI9p6XgEg6zNEdH
oKLzDi8MXBmMsMuEPdAw+T1Q9WezCVNWhmAR5swful5Q3ho0zyUkF4SF37dwIVy6RAU+58R+awOI
qE41+9amRPS5HLgDff+0lCu1wjDHwSpKZwBRMRkQUoLzD3fsWDyJJP9lo/2A5I14eQli2bnbcH6A
dGqM1XQuG9Cy/7M+EGHdX6UFPSHFXMBs6UaDkgHyI0RaPXB1cS8a+lljfJhPtzPCNgApCmQmcc0w
NVaBUfFTkdPRJVvlwFBA2q2DYYz3RAYcBKnLDVGzCLrfm72HOhyMkG3SZCWdBO7aJ1/88GAM0cmX
HcVfW5rldmjIkHULwhKYEKLGahvy77mE/Cmn1FsquP2qgJJTdyjOLNuOHdYqR+LSh2a+eplBX2AT
0OCZHzgxVySa0w1fLwd4CBeVgCdDuPRAMvj6qnxvR7Efxov1iZ8X2nXfnQQ3FU4iQWFkKXp1mdnf
lnYlMQsEkDN2OqaHA2/PicmBqo9+gHETEt14eaoin4urorG7eibF0BZWT2S8alOj1gqgWeC1Ji6u
Ve1A6V8zgfXjRePXbFRB6jCqmP7OfghuqKWFD2ztyzlDhbIDzGLD8ydxahrnsCZgykIqrzagHK7K
rE0eQd6ALNhcrkgD/mOOKKMnJN7d43BQr25PyEFVS4ybkasO09ssFUu2JqgwQcGYx47C1qVTJCMt
X9lZjEDd089qlfMS3uIkdMen9m/iFt84KcJKQfYBasrRj8TPJvbxsX4tlQjpYrpQlvRAJ3KjqFE7
LrWVA9BwnpYHCahRU5+7hoJ6VTBvljmv305qUad232lxCCYOpLcM7an4HrmtkebKkcKEh53TsQ0i
yY7aLinIxpX1I0dLfRzjkN6FdH4iU3DbiJKQcIdu25GquYZ0ZQxkDy10VFk4gGeL/II+8b+P3JAI
bItvwk/LGP4lynbk/vPXtqT3LaHL/R2qbIWKpxvyjfVUpDsAJU8T17EZtFiHEKMrnZqn6oKMo13c
yNyi2nMPefuNskIJ3nc43Z9Q7o83MpYzLSGqzdpdZfdnXSeNr4ewjZXStfutoaOe7dIDtAoQsAgQ
v3TNosSSFnvOZp8h3XuqKhBf78k5nyh7PzsL6r/ZNQXudw95q5tPPV6dPPcqRxy8SaICcyx9Qbio
EuMbs2BWM13y+kfyl5Hnj/sS2itMwxnSR+UVjgiBTr+769slwUpJzU0nBVggrBKIHteQOGwM8IFr
D4kw/vWKWl/NNBtwF0ragOvIwv/UnnQ8sMbYyiH5JHon+MQnkN3J5hr9LYbVxJHGVgRhwbNoZ7Kb
tn+Y2I3ID2Y9SUj61qK0x5IgaupVSnawsDiygj/iLJmHqr1q2MHq5ieaFFOAbdwV30Yd2EkuqPNX
DDShwQdyNdApkKq4d19s8mMDnb9Pke/V9lldPI1pjNzTOdGtSrZHkIKo0wlA5tT6gtWb7BQjIXiQ
SuK4bBoZ+/35JgGQVhmSv0yEAeWrveMtyjilWteKjrj7p+uEByC17wssdnKgbQecPcwt/7JpJ0R6
K3lGTJX61xeIHw1HgsLJzPA4wm6Mip+8XpK0+BWRi4aBBH6bcBSIXfkyMzdbsaq9f1mw4OCsv7bh
jk1YRrkGf6wlfsO4/QLdcOisx9bjc9lPDJvavweuU3ugLu7AGk4oyrU7YfPcnMvvM2RA6/XvSi9A
W2pr6yA7X+1nZi+GN/nvZoU8aU0j6WzbdlxI0a0UKYG646uvpr6536sclral3hN4fZcm+aOsDBjH
3VevaUDLqc8pxXWSAOhOnDeT7Ci55zMfSzO/+jAUBEF1ivadG/az2E1xWVg0nYwII93FsyowPsDk
x9EF53EsO9BsQ5ZRhXpbIfAGQsb0KdUSgYGHNcBYMnIFxnInpClxC2Lb+pNxw8tW+oIyEtYGre/H
aRD3bQMhs8Mw+VfKCwO6iqM0xFZ4nXqdcZMxTYC8eJcAR4dvKVYLZb4T6lRlz27bn+SzzVkLEEgH
Mt6SXqXlA7dppq+1TCFg6LD4wjAn+RIKzyzOJ3PkzeY+q9jcUd8T5V5YcPrFyH5R354vF7HjClRW
1Et+/puNKCoGbmVr5qwgRgigTHD3Ukq25w039IO8m6bIDHwdnENsRFbAarDBPYl90blvSF4TF2vl
FogYqdJz02tjPfNfwYKWkBpEkrDU5JT9Z5LzGy9T58J0HV/ZLKlCzLbQeE0KACqUh22ijxOTyxNp
Nh3527LtRa6W9qVE97EBM1pcRXOvF8FhnZ+sxk3rYgXvYtcGbvzldNoZkKrXQvwLWNCcfkMEPE+u
cryd3csvU919DhmxBnt17RA8AUWiDVYzrbnuV+RAWKImFQ59cfH/XvQroIvh2bYV12E6bNu07g3N
SqLePXZJCrNXdXooc6+C+WDJB+mCciUgfyrBW+ngM862KpfIGFq68mWROmNT4+FUycrO+AgTNE4H
nvqlc7RfLMAfDSKhVuaFv2dY4SiPlmsSsojDvvY2fiFnEBm2vqD3wkUfFJT6wtTe7irJg5ef5AKT
1t8ZC4VAlXJ06+TubyA2jIzVk2l/CY8l2VuZwVNGoL4+rYSRImu7lXiBJYhTAVco8oBSSNLVBh0u
5pXGNwvDCcpUAVTf9J3dH2DfGGKz4bM14bhbbG8rD7lk1M6JJspGeH2eyrQlBFuwgl4kZL+m7UBD
4ujzUvEP8I+QR8rVYERLLseYx1iKIa7UVcfC08WetNZIGEB/RGLy1H1yJ8GQZZx6HIJkSu1fHAqc
9dvN5XXBYL8zdlvjhnqHKV23x3sI0xMfasdJdpSMXmQTTqv1yN+4JVjcTlbWX3cyfdRWdQRA+Eh/
6zFBgKb4DjR2iK8ixzHkNp6jIid/jqaMQzJoJK7Umewuin0BWprnVO6EN5OpCxsglDMYzH+h6V6I
mqmiesuU279ScmvZkA6CLyX2+AT4wd6ppWiOsZ0cvGSPeaITp3RM+j6hli0NLNh+Jka3nqWhZJeT
ZhV/eDY5Bope5J+at9rL/UV1qDhPgMFBWEH7NEcsAVrxqZhMXM9QVuzFjiaw0INNhkEzfZZnWjgk
ZM+lTfILTX36WCumIq0LYPashndhI+2i+VhC5Sl4EYaIg67PAOqCfeuLs1IWhNR4TJdRZe/8mzsZ
mR7YfXlQfBtuCv+3aPceBrW1mcKjOTu3Rkf6zES3kNVq5A9UK/9ctUg3TgtYj27U/KhVCN//R6F6
vnS8MjV65j9YDg/ygw3qSIvEMeYnkEA9hJ9F5SkG0+87mh7Q94FYpY4ucLT4srVcMzHS8r0vC2T5
x5MtxC2L7lDilgRypd0pyvoQIN9fDbhs9BK8K/+TAjsEQI+JgAlv1L0yl3Dtni1pRImOB77m+Iu3
+IYT7Mr3J6YEWnxihbv46INpTxeQ5a1AZY6Nnw9tOw2qZegMt3iNNqpaWDIv52eib2tF8UrucAeG
LG/bkAxneKmI7NaY5Q9r3qXJ1AFUntbAk5y6XYxbI5G8cxEMHODM+DyEINLTPUafJwbMFhDph47S
RWejV/J7cIQdkXqGNKDzlt67g9YzC0sXln8IgTreJZ9pNGjXIi9GKrpzl69/nQ2tTHvz0GesDtgd
7aFUcqtiE0iMkORKp2Tcyk9FSZhaPSmMNLZYJS/YVwRDKFL/RrJCwg+AwW3Us71timG+0l/ezK1C
mdgz3EwGgbk/ezQYklkTpXL/exxPds+N5qlSGK9TSQ6PkMC3AYGlAQ1ts3R46QJZUqz8Gju0/VlX
TKAzYMFMasF5Uezg3ku/E7Y7RSK68tuFp2PyBFQl9wW+CnlzDBbVongyALqFbM0PemeKNncpsilb
J3DRL616Oj4mB8wJGgFxDKrVqMALIpHGUIZsPBufq0IDjZZYEYsKUCqckImSCz0Jg47iHdcvLiCw
jX8y9/jf0dn71Z2G0/oM1h1Dm73PGaslx1h5mMV8hxDCNbNrbxK2GwDUncfIl8jm3DDE/Q83RH3s
zq/bCc8SNPXhlX94jlpHJBgE4cCK7+EaLxJxX55GOoO4Isn9fDuGQoePsx7A1t7Op/GoDmlLuYhl
3XdyW6K2obiDmONx3JLzHzZDljgJxHszbuQ0GyJm89FvBMOWx1aEIkz0EdTa6mAyZXKTtTTGdxQ+
hyVG0XzCRtEl+M6ii+4k/yUTREi8auqI2sTFK9viHMSbUc3QwIPOPXCH6MBZhCjqYU+IkbkK7mwC
TqqUicAocdxPfokYBUOlBBPSOCif2dQpxXuKRM+gvJaj+yt3KNQBVLVAU5VOBZ4q4BagdlobALNj
hFeLVcyNtzFXMCCk5AbokOAaDzrTrCMNgsCFuArliPTjL4Hes/C+YaNPGXiJ+6AK+TC21QW/Eoeg
/i1GXNpos1Fa+r1xhLgkSgXjAAJvoWlViNu8uJkQOPkrH+gEH5xPDQF96fmr0RPr82SaS2furX21
XSR0qA57CZgB4imZ1O6Y/2phDtQk2fMdfDHKygJY7eGrJR3CkFtX3vVypT/eIotLRC1bjUxTYmZ+
plPWYJwNySABbn3JMMJEtm+3n2ILm9tYf7Yhr/S9G5oqtYPxyEOKWFDAAnUkZlE/kcrNtVdIoE3R
MDbQK2Ev7j7+Z5Q72xoeVm4NfYG8962+rOim2TIkXk8FBX6EJuSwaM60X0o4QITIS6CxGUfU4KZ+
knFRoLUm5B31hNVjIXCSgGDjy6IhTGbNE5F/PxtPQAJ5AVZLQQeXbxWSArVOH+7tKCiPrqJGifyy
bIlDEfWN8W0cVQZhC5wUDRbJf6j93HRFBhN4R1o8SXPcp89eMHgEGStH0S1Vlhj+3/dEbqkE7WPZ
T0mbwj7PMT5xDr8Svmf5doLPWR0UHrLY98Fx+qmFKnmT4AxctX3nl/Ug21PCGMu4QYWQR8Oj+hB4
PZn1mLb6j13FcZ81nTcEq0w7qYFjO85+DGMmsvPERSRznH6LGLHz+ryvZWS+ozwLjskr3IVpBrAl
nos9M6f+mHlhnKFI8/4b7usvzJy8ZHC4kEi10Gd4BST96/vehxWVh17QEIfUVNYMd8yTQAjGW0OR
6LroHJ/pR6dsWcF4/4NqWf7o8lltK3HNyM730CvOtRAmP+2dGaS46utRoUkVvnEYWzht23lIi/76
ur0CfPdIjmRWSC8bPQSBnEl9m5YzdH9cYuereNQMwAigi54/5xp7P3FzDV+n4ZxeEF+pmNVCBS5D
lxlYCwFFqCJnUOpK0JmHRjvsezOLqchmi7xpbFMoHyFRs93zBMrm7Y1foWo1eioCkO2qBJ8HT1TM
VaeYV52w1YYdkAmEU6nzRTZ8LAg2+ecKf39YJk02UhR0X2TTLfLwsvhgDQWnIKPmIli40vBLEoRp
RKpooqXjd9DSwgBwbh5gclJ8fXuV66JnAGP+44oUFRl6g7Vr1tsbz7iL8SilUpVRaT6cnJRBVSf1
m3QTNd+eZrweVw9i/GY/agQVSpG5P/INsZG0sZvhuNXFeair82TmV1gdAzpPosPhl8Vxv95TvTJh
3khteM2iuwdKwRe5BMOAMmLvF5N3DXfhJzG7EJFh0Xk9ZSkvWVOrs4AgItFRt1r1RhKfWyRzWAAa
POy2mfalBjl4Mt2LRutLDFZwdefAZB5GzeonT84eNbpmPTf/X37mpDHzFGqEEi3PYB/Mz5EX6gZi
+G06AEh2Cl0sC1x7+968zIzxsMf30np8wNn7oT89zl5Dv+X6VSl0OdH3IYdUY6hFsYWaKLwF+NAE
rDKbRhJYlliKIeK+dyutvcpLp0cbnuhZzNp12dPBEWw6jRb0fq+SoaA3Q9nDrjCVP1/cNmZ+l8OU
r3n5aZbX2dEMzntl39fS9MEwbmPpPvo6OVdkdussAvWE3PA9g6UD56xi7eu6eHOmSo5P5Hqo6BIv
UszXrKFICaINwSwvr76YMOtR14Io8jVfWPRqQcmYrN3YE88zTuY25LxVXn02j3/TvIooCj0iLaXQ
ZprMkXm2b8OfU5RhhMmuZQ7Q2Yg1GWisKS9XH+VcUQdHlDUfQgSgDVGHJzKbr1Z79uLPGnV9mHSo
9B8U19KjtNyXPsz8w8bDXazO/zYtG2W1N981tQ354by8/91CzL0EmQhMHmXDY5JGMZpoei2gCIkp
zS0gmmnRfcn3Hzn6CuNEkAkD0jJK7bpHocRRs84c9akd411hX6OHHNkazbEAPX/UOTQZer8ojDAq
lCnh+R4JVcVUajij0R1NW+LvfrgjsEsok0J8hNTg3r5qI1u9skFKlx0oRBfkv59F4/KmD4QPXFGk
CYHuN2tn4HNEiyvA0f2IZKmgmeCqsiWwRX7/AV1bT58PmfgSargvjYeNz6F98nnIsHKG1e8H8du6
bZj8hZf0DA0GBy4ocu2LbfIYplN09V6wr5+Ozm1BtKnfUde/0N2xJOhk9/BAmJkRa8/QwHwBqy4p
GDwnkkBaVtwNKM+znnEGbsAaHBkr8HKCVbXPQ+1XvGjOjTzOcscrXKTO+zC3gDXM7WhwVoXOe3b2
RZXFFDkcpi7F9+XBK/ZBKQg8g5d9xqFWdF4ORdtGTooFVvXwo1juoKMEH2ciXevsDTMW0RPml/4U
478Opp0+GHJMvyuWpEcAX5bRebOD/Gawb4CpPHf71BmiXTsrDzFdw9GKUIUDOJv4JBLtSvSWxWpF
rmxzV+P2AdeJ4D3xuxHYktsYdwMXv7WB7UYLS5Sgq4bUevF4rE7fqWB0GAY8MKkWBwpr65HE0UUh
TgRCjtPtfjwzsEmjYdUBRljnhSSAXbx3WLb4xxhHwLY3c97503xTghsbNFYQWRAen5Vie7Z9nwHM
8vRHaUwzyofwEXivpBxQsJTWJGGFLvtF258nw0WjfrZuH2PqJZRuLW2YHJ6ygS+MGOEpnJQw4/2G
XBN2spNS+nwm87v9XG+OeNzrq8D1TE1DUCFHVXNi94ebPnnPb8pG2jg2HEdVr04Isx/IizH6PzXj
Loxmgi8S2WDIXf0x4fcgwa55EIPwx+PjdjdpWsZD6KcloEcLRkmkWw7yiWbIRaMJHTfM728uGdE4
3LbF5/BKyHqluzTKRYMFvuWo/vexCjCY2sYJ/6I0CQGBXLokBRuTjWu52iYsMbz9RFGlF68Znzkt
6+0OxAFMQG3diIi7BvEx5E7+5ZCjdrp5YF9IGfQt2DXI/L9vf9VetIiyY5D03psk2PhRB2zt73iA
lkvQD23EyUqILybhejp00AssFJz4ZxcXj6IvqZbjQdhjUDT5rbvyLnRpssf8i/5fZbn7ulgHKj0r
VCUmavxNDfErwFHl6z2sH9/uaZpw+PtOirA1WIoUqEZl5roPF/GVxTYmBUUMptta834BtLDs7ymt
ZNxsH2/niJQCzr33gqch42jp2HOf1JQHmCI5FxilLQnIodT2m5DOQmqu1algjmyBqERxjA3MuCrQ
sQF5o4msFTPmbkFbSB44jh3KEIoqGY1N6NJxI2vvlZUpma9+fDmIEA73kEDOJ0CaqhD5uvLvPC3v
vBd5gZrx3c/EyZqqSSDNpgPKwvJYznG7bffUnjQmwsxfAGzoyyjdDI+Z38Xgsgutwr0xqoMqaCbY
Q95sC33YyBkEgeAqet5kNfuwSOjydT/vWY0eZ0vrBd2VUcd8RalP0pIxbir85X/S5GUFKU4iJEx0
n4Ygxyyn7YvqsK8MMCASfMjIY+H5F1U8PK/T0QXykYz3B00NIJz6tvbmaiz5T1m9sgGzMCWblhZx
nhoM5mEpvOwr8rZRSV5U59soZ3IQfyM/TpB4XY3BqauuEQEXCgBwZSqFY/ObW1zc58YSnzKOxIfF
gtuBCVnU4nSYI4fjZsVK0nwErQIVsWnyZF697a5qHqAdx3BYErtlbGcDRI20bEMqVt3PNt2UEsno
1DjYgXmmxsu9K/yKxYpdrpBAVPclAeoGaTeW+lMq8BuwW0Qvv7NpDtvp74x3KVJW/lsdHIgKy1a0
k/+QbKFB467J/h+t5m/gRD5hjhQRlOD2OgXhDeq53RNFvR0p9SGlrc+y+SRyJMcSVJHtzO9wgivB
8kkRp4mJNGOqKoKd9hCvfrBe91nDBbTlbW4evOqPzDc9WIfn0z8ObNJ2mRJiS0sPBe/u5C+NbuDD
nJ0viHo/YGwqDeUVQRt5T6H2WTC1rABp3aQGFv6flJvvA6teJ6Qsae3YC89v9cdRO81ot2MyyuoO
lWXB02nVCpf5NfDTbrBebkEQyrK0AZ7QX2UsjscWc6480POZsl9rNA0J6soCtnlztk7xA4ljfk0J
fryQKr5sEsxOkF69CTSFQaTGNQHkejMuYLG3n0QOqqu3Zo7zxhVEw7438f0/g7S7DlDpqeQkeebQ
9g8joYuMJmrkKv3OMLU+QzRQPzDsZ4F794WFb7l8JSpAe1VEsiml+CP9r9tJg71cDHnihV6TRtsk
21FCH82QySTKoNYDGkYW8PC940SOxv6YX9SLo+Hnwi5RKWLUuu45a5GAqS0ebHdDR6dUGI/jzC9O
OQMwVMk7PlUy5gxz+0nWrlgXHaPsCtHy0bdAyl55KvL8w+eioj4DMw0cnUM2/LQWskvrejyFHquo
wW9MRoBlfcFRHj2xb2+KpHa9yoQbO6sxhAcYyMi384Dcry6hX/6rflnNBwxcd/XGTX9o699SMK/V
/yUjuEN97DUQtoqsYwQdW3Axa6Dchf1nngaPvjcc6l01EjnobK/epH0veeOS/KQ28YLUhY42RmWE
uIIQBNBZdZ+MHeTrbETDykAkSCrrtCX3kGrtjoFzVtOCzWcr3979flhHiy2rkyh5O8wfkrzjd1C7
xlncFPV8CTKOLvBHgx8KSidhQrb3kLlV5OovIUdxfbJMPjA/H8Ris0zUECAGndO/254ltcGOnS+G
oKvedTOejhClP7aqTspxfcB2npnxQ+yiwUeAHmrbwfrFtGPICxNQtE8QzawWqaAXeFa3t2rr5+46
i11M2IsidaJ37r8dTwnKZ2KbetGdfRCbuObDnfMQ2HqbGTh8pvk6uv3uDmTs7Q58OrKlFGMG/3KL
FxpjWM5prhkT4vDcL3czWSgXzaAeM6mXQqLqNwT7lYpIRSFiQk7MjXgYvm1LxMWKOGHBFyBPW1Y/
oAOqRdFxYyV/kLFf2LCQU5P3E+oe6MV8+IIgkFjlpRX923aNXMA1Zjx3bZpsr4+/2KnpnWxrpeEl
ae7TzyyDeYEghL0QYPDkubxH1zbY9eeYTAiRoq4ctfrdYCWYqQ3IvIQ7G/ZuVoty1/p79JdGkQlF
bEj+8n5ZuyNsdjygdxh1gtsSFBLDgAaQV9NllyNOx0ajWptKAhEqAIN1M10KYLqtadLKXKRDSoFz
IpkwlLxBiuDWNb76aAJK+vwhmBKbUkb35W/DOOlSdENyatBi/Q5nZuTCz/QlxZ4ShRxHL9TWQc0N
VdjYLRP+I/1PvlAcs1+0t0RSjGJXHUu7hB+9NxKwXEV5PQ/Vs9HYLSq1zgsvefobexsrVAH3OU7j
PaYp+FupK+RKp1BlPvx4unYy7ZEUYCF4LbBFdQ21Wjs2G5b7CkqdkxOCnCjI16vbtYoXYgMF1R5G
XSPfraQIeS7Zsvd8/PljLprAkFD/5n+PZiHf7OHIzFPLhiEiJ/+yoHJcIvCZmJJQHuHZHTGrr0+j
iY0Msp8obnYk0vNm16nKjUsvbYWJ7iLG5yBwdhhOaTpmvtR5fUc8wJtOfGcjUqUUcQpn0KXHGPMs
qRiNJXqNToQ0QxXfDJl95giqnwNFXgEmURTDKC27oSp8q0DWr4PgRfeWqKVcIzsrIgOlpdpg52Uh
I9uh6RuZXpK4BFXTQeyHMOaOpJlInrkna7KodZS2CjIPnsCtiEmisxuW2UX/gpE94Mafu406qvLR
BrUaG4kmyZ0gS9smTo5zT1wo4MDmEZUlqQkc3aA4rF/RKEfJk+U1G/xn2LIbztz1enNs6EgVFVf6
Ux6DgMXDAPBPeu6CgbwCK3FkvhHtVArUpWPoUZ5CusFVS/LEPd8AyH2hH35QLJLe8JY+2dMrGuHa
7LI8tyfBdIH3omrwKn0NM4udIjhx8nZKXf0LNLXoFWiHG4ZIgOLNn9DbdXpgwve1E8/1OJgdhzUx
ceXlf4qrDfq6wR6y25Qdz4+K3co6s/T+G/6pd0hQnVAxWdEUVGFoGXIHJ0lQumgudmIr524XdRmB
zW0vY5b879IUpGw/BmlJgIJEDLlcX4oY+c4ugVRkc9le6QqAIS++ZryAlGIOYrJAA3HChwGjRK1O
+aQhKXWz26GQozV1dsf1rzbXMnwVowmJr1Eozw/1Nb2kiOc1NX77JlCwTrdtssMb7dvGeojaXoDe
Q8LvGmeP5/3sOfRi3ourJW9NkKPtTY+QtEMCUhtKEMvCBqVOnj2LZVLHyde1QwQlDO0aPyPUFxBT
xMM78OH4PaAT9tw3urK3t82lDQjagzcH4BuZtpcuNqDC0MIyALWKgvQcUv1N/ecZygIhQd/av9cL
9zl+iilw711JwP+sCQ6Z/uFPEJm4i32iFZXgWGbVsq25XxZB5I4XgK8EOtwZNAHFFbSInVwy1AKZ
GH2/LUAKDSE8QOwbUa/1kk91VMTPnt4jjo5jw76wG32lDdU1ciLBtb9UTSKQqlcLXQLUAm2VWvYz
CTK2R7OwIzhBHcQOMgDZUbX8IlqkjQbcJD487Nv/4gvUgXumaQb8CmUEDDya+7MuLmZ+PdBSKGyE
wglfnOCRSKsRJuKK9yXdNI6dGHSQ7IOcAI8epAriS4earUjYN6f2XzYKcCI6gN6QFLPy5KP6rWhZ
790UbHv1H3MCJvq5AtN6Ap6dv+pSo87vzcIK6JkVEFGFvrERKpjelcnxRENoL2+Rm4wOXvZ7uJO5
UgoIVig4FVMcl3OByTkq5xfkMe+0nVGeimDokAyzOfGZmxCWmMSix34AUu19vZ39yRs5MnyX/9oC
9dL9h5JAw9XsAUHjRKaMxgrO52xf875Osqd+m2TSgLGnezxWyzUd9ndLFqh4iEMDwhUi0rSwFaTf
Auet5ecjJMqL6d7N8YMfrmISscq1gz1aZH9a08gzhNmZDvQXWjrmO/v58myHJtFRCIhfXp4hyXme
QN3jIb/4IM80XuL7IDan2lGHjOl9KQQkBjn3gl/sayvdAo81bBG9CvphtH5Ot2ENSZH8NwyCz9uV
jSJHGQ2OuFa1dYaPLdP7gIT5LNoYkk0BGJd8y17MomG7K+yTB+Rxtr95nxXhE1otw5tN6dnBdzQF
jaiMbd7NZU4BFgy58AZi/jybaBkKIK5uY2ZI/DfTcvKuGRh4KAl0p+yNE/O/Gmt0UD24a+Bj+IEB
hinKyKBScfoe+E5ErY5gfZMPHpsXBVDiwPV6MJha24fXWJOL/ktl1QbA3FU7RzbM/lT8nr7LjPJ5
9iZ5mOoU9TlZR/r8AX4HzN7aJJADEuvwMgticDrrtJ7R5nXYc5QbcIqv7qfs/xSehiGFV9zD5ghJ
YmEbDL0q97v6L5QCD4lUz5reoXBNvLVN9KpkAyYlxZfhlV5scCJHayAMMcOypYQbE/Nic9v7ND+w
Mr3gtS+6ibT5CLw+kIhU4fVswPBlgiFerwnFPu5tgstOIwdAlzLCe6lO2yhnB6lZrkEdsEveBoa+
pLCLcK+7atPQKTauPQauEpFJtsyUjFpkUqlpO0pe/mLg+eYhY+0d591GDBJQCrxLnYKbaWBBHaBK
o9EnjGXOmNdfKGYbD4pdVs29hQpxqZpa8/CjzTI8T4u+xHgECoqc99fADD63WDZnqdOULW+2JanO
5xJ1gR830bm+XKXZ4oNqSGof6GFAjgu1qo8NObadR/cx5E16WKU1aLBSj59MpZVI1FnbyvUYhGDL
C3Vr6WSFR1agPnyVvViBXQKtvF+vAairG56FEzw+t2v1MLEPUKsTvYWEY81fPj327AoN7ptlecfL
XeyITbB4cwl3aQAjo2PLjdvfhHUXdv4aJP5PzmEfzWgefkJyUgzxnUwoLQX8RnimkNwGjr/6cpvc
lcYmNCMJ2heVr6nC1b4ccrdUUafVHiEUBFqDPRq7nd2SSZKigU+tjFH4ieNd7q8hHMxagPI7qKeG
fwkvEqySV36fQWuq2hJfHhkOhFYKQw4QMqf8PihL/ZAs1wamK2n7rkPPtRN9pGTWMyB7nbqUqRWo
l9/3OO4s3V0ZSE85sfrdUoSH9v/iemE5kfrkun6Oy3PfccMR7WtAvGAI5yxLlSUKAjLT7do6V+6s
dcOjv3sVjBZfZk7p6lOTA8FmjEGRqzT+I9bB6V+bBiijT/fY/sqMMCcvQ3hsM6kt9V8Fl/k5CXOE
QqnRygdUnrTlIM7yuKW+92UFqPDMmYPXP4LUbnG7qVevuJGhfBMQaAnB0tchgTNmXIk1yXjmcEw+
Luj/79EhrKR4MhEJTui6VgQ6eFIlYL45b/is0q5q9pVTj2NwxDSUK9cNuB0TKfyC1N/w8YnldgsN
BIsh3UOX4EBdOZH8SrmziaqQupdqUjGd4iXQ8MRqVuzZ55VfzFEQWA5Lx5SYKfKLLLzIH6x7EC5P
bdfR/pRB7OIwD29UIVonLRHYLi7QjXTZKXzLB1YQYKie1jLyZ/ibkKaDZekZl2hsJKicDA5C4Wbo
eqDwIhjaFoZUYfareO+Qon+OD/LV282zDxAYLzAnRyqzn3t4nyitUru4oynq+dzAefp4dA9CcXiJ
e3lXw6F94ZNkS4aKxRWTh5UPWd8lMPN/iTyGcI6qR/ovh3M8Stv6+4DfQYJZVdm5gUeuBP63TIwM
ZcD1bqYrspsoN9eHB8NdJ/GJpwzVr0cQy+dDCH0RP7sSWKggx2Uozj6dshTWeGWzhuQ3aeXw1Bmd
umpD5+a1h5IsrzQ7pOtmYdoh67bPvC5BB8igBGcJrlSMNEU5srnxl49d1ysO47e9Ezbp7zv0t7BJ
zzm+YhX25mCdwdtBOK4RRJQGkGeszDQqBIYA2lX3douhhQxtRNqwsUPXR76Li35YpJXaz9lEQA72
OwQm2Pa0s5W28ZK0j83ULxpWtSF6qsiO7KW452O9/iUH25PfbT4TvfSx2NL28LUlqVUuewEHUh3b
Q+PgljkWfv+ZBpkfKcH4R+0Kt5xikDjBM/jU9p2L5QoPVbJAMjDj0sYUDqHBGqt6me4wcCw7fZme
j651HiVLtuyNOJj0fWzVnkrry/ZexgqCiLw85grVquOXAwnE3sImfUjuETl8PHvqynBWxekyx2Py
tNhQXgzj2J1rOnyAkb5Mq/6IDCIYND10zvoIdEqjE9W8LRM9l3O766bhwgf6N+0F90w3xHhU7Lxp
jBwDFnksnzM6BLbJ5ZHUvUkugty/sh/rrHH12BCxBt/KL++vQX3h/UtnXpE1OW49Cka53GJELi+B
gNzXoK1oFKBJ3DnMRlgRQU2Lglqu9sq+TwmsjkRKHeGJERKrYcF9BaU6xaTTaDVAZ6hBXqXq2Uol
g1Mm7Ci52uEiPKhDFXgD8Qw0/WsiMMxKbErogJ5hGc4eU5p0rh7QCoZdjm4konQOiaHTOGq1eDJG
IWem8TlFHtcjwN7YoMFmoWgvaWBkW/zW9cD1z9XJfY4BrPzpXnPJ7F/CN4FjPFcc5KitslxNFlSz
Y8DfwHo85MnXFcSUtwrJfDNLfF9zU9n6XQEg1R4dZiWYrvl9vIJm12ivPLTabNcY0cwe/G9z0F3E
yHM50joy5i4C3OIcm4qQb4mV8dcYAO3e7YuW9SMmLaAO9AXIsq3NIPJY9CBpIdCHOldWP0Tp/u2p
AKKus6ZHuDFPwNWrun+3VbU/Cfp428VzCxlyCnk3DkflrzlooR9ILqK6qr/w4Sb9fES1W3FbC5LN
0HGIOMM8eVib6O5we0M/I5De8s/Nzkx6LliKa/kdbweHZAprQf6Zcg4gRz2LzjPJKhlaGDiD2DKg
vE6czyLrDZOytJUWELEEj78/YF27FqWINcdRGoWRtynIoF+EXyfhMZaBVz53kfR/gvjMHb+9VBW9
fyo8NRNZkF+a5j71SyrWwsn1F85dQJaS8kKoydSveqSQpsxX3Dm8UOv13pxV+kHAi7j5S6hvuqHd
WbvhyBvSnMRWMsHDOG5dhXaesMUA7WLr3SYWC/t4BOphe5VuyDmtkJNUbBaBpxRJK82xBhSLQBRa
NGVfWZIJDeaCLG7+yB47ZF1afcoygOLb5jj++CFGJwAelgehKZ4NIL/YrI7mG1wI1G4s4M6nhnTM
usfOeQQn9kAiJda5J/jAnkNRrAfxUwbPTjC9T/mO7jjcCAnMJEqB/uzC+vrpbyTrwW06oL/j6rai
cRb5DttV/exzMoYEQ5oAJkKLRTKbwTlqR00P9HfarzIiTA9EFWOJ+SNI00OjM4lkwi4LTXyhKtQg
gSOByFNYKhbqmeXtPjMYQTMJF2ZWfZ0ppdF5w23tQ2N5bvhmkDmVx08PQpPVXFuIKIW5WoZqfPFg
iAljCV6UcIuYMiPpazMAotF5Pk9uXwG/FtO2ZrKRtSoM+lEUL5bDXASPpFr9BVYngwOze3pSKfrt
pSEklbZnAn97qlG5kULQG35E9el4A5S0yUVeL3udW+pIJ8lKysof2+IkfPMdsNWCVi75bByZUDuJ
dlQgDw2SZLyVx1H4rjXIXXPNrrHqWcsnAyoxzSNmstWQ21CAB63SfTWn1TvW0lwxcLUSZq9AMLOn
cXJZTwsE2NaIyFgeRPSyoq4+lGnoc/Odtb7bzMINRUPog/qadHp9atrbFywCphRytWLZqsz1XECt
QvyMKtaaErEN8uRcZqZUXI6jl94ZKZ88aG7mwq1vhi15q3KrgKfM9t8yVl3wl8Q5FXOsu68SNW4p
1Zspm1rAsPIftn4DRQ4IgJ7G7Vq1Yow9+xCz9dovLTruqqf6iHwiF0DBy0kvRTSsl92mJauOyN5Q
/DkfC2eBVIZYd5syRNmlt43vJ+WOm8w89DvaS6+ZTmfY7o+je3LMBwhl4e0bUkXBMtAjWqrfZoch
UJYrJ1BpXOg45HQP0vgAX8da0zaim70RipT2LCOv8vvl7LanKMAXxorUY4G6dyWez0ZSj8WjS58g
sVpddFhebRZlfab0PTqhkjzmdHjlqbtSz3qOsn3ryyYzxlY+IKO6fsZYgoHCI3AoMsXmUpaKmWRz
zkWwPRJ/kqwhslT4eIV8nQmgOG0N9v0bpxtShv3JdG2veQVgDZy/nXsN8oSQWqiqOaYTh15N/bvw
7ECT3WkPtoOvv/k01iWLtgHyqDP4Ek1rGy6w+MpNKs3XAEEDI10s3y8vSI5jeJhh0unRamDEDBMz
XUBObppRhRJxB6OGa6iCazBGjtMlG2OeSlTQ9EKyCdP2QWWdBY4vT9uIaLv5gMUMcExvPhElmHC2
EbhNihodM5WnJrQsKL+PoLViRnFfM8xm+VC8UHE7P4wZBJ2DZgqwMfCTizkPweiGd6eSQQOiyK1m
ouwvBi//Q6bT5IQ071XW3fJ/EUxGA8pH3iAoeP8f2lXnO3JYarMP2usO9lvhqocyjfxc6bA88Fil
6C1EUdXyTI5xAZVuN1ccYdwlTCZ/2QM+YUOafxLi59Ke0CgQ/niG/D9GNNWDnHt2dKEcSWfqX/0k
hrIEFrnmF0Hf8ZUBVwSX8UN+OrrOD3NSlK465xWbMQNYteAnbJh0o/DxCs6uN+k0VFkzKvn8pEag
ic0Tr8wrPUUzU41Q0Y749hVh2rb2Wod5ZkzMiP2e1VdKbDzUG1Ji11bKDRQiJvi2lrK0LUhZqdJS
VbXCrwkfWssfhmcVcwzvshXrT6q/xWd9BJb4HjuG22jORs9r5JZPmZLi88wDKAAM+meS2H7hSHHx
nvwyT/3BligIK5yd9uCU/pYsmR9qJx20JrxJTz6Ry03eHq4m8hu5/vDl60U1YEEMeqfjMBuVIPqo
j8WT+HTN2f8bPWri8+04rTRyI9sY6so7JYvu7QbvJWkfveGcR5zE/D6Z9IRwmQT/rX69tct/nY4i
VQc6xfQ6w3m1yl9+0XV0L60Y/MXCuGpOpJ2yx8ZFyRK7slob/P7poLRYuaIPrKAeHDn6A9a2oWgc
yhUhIx8EwZ0Ctjfl2SlPjOThRpKgpPXJj/rVetUdQu3jq9VhKKYaRqDfNb/hQ8N9UB5NBJBAhHcF
TcI7J1okJvFV+LLJGWK2mZfnK6oQaPgtebIzd3KtqhGJ8NNr7IChkQbJE4Yh7Jo0sIpMY6x4AFqD
j8vLebqtsDCfHc9BwlsSkV8CKv4tw85lTNr0Ue06Z4KdMozZozLhwCLH7z6F8GopJi9qtklZoAPQ
F14nb1v7Iydnc5ukYstvHaBRuAgky4oJDvNlWjaQCtF0qaTz0Uk6I7G7H/164UDBP8TIR59qHFxW
j3ndkjisS1AZ8j84aLceIgidKnqkhWC7lSsl8VtwDzz/aTSr4tHQK44Otgb8CyEmpmX0ti0xmYDQ
FtLg0UT2Hl9f4xMwB2a6CZ1F58agjJ2ZJ9G5nEz0Cio5m9JfUzI54/hf9kYBAozVITWsmTOwfo5M
irDa4Rjc7Lh3/KHaG48+8mO/TMmxLQ8LrCw5TbgAJvWanCn5zlP33dueTq4bOUrtF6ZdaBcrhRx/
Alq1J14v207i/b3cmPV6rTz0GDOKyM0OyX/Rl8AGyTx7s5Y8Z2jfSge9BjKgXDlE/TQWsoadMBHl
1U5F+KlIGHp/bVshEPICaiQNR/uDSivnEPbUTs3CRUHvtYau1LK+QyIP/cm0BY7yJAuwhNJNqERs
661B8Oi7Mtzc5PnZr54MP8YzeGsATPUzodjSgGNaSfqJIKowEAQQvJWGAd8EHiX1+fZ91VEjYvu4
rg7UC1TKe0tfGRezdM5m52FKF8EbLTPw6gj5MfrMD+qRwbfOKexXsDqJEQL6myU+sUyirBKiaKcx
T7JhtgVJKI2i9kWwBOAgp1oDy0hUl7hr4n4UAjbTcDhL2TCpjKUAQfBcCsQrmAPJ39QA288Li/uC
/0pmut1/SyMmasnz7qusW/7QJcKY7pbi+gBYtiQWn3tB/QovUNNaLfac6AoOj1kF5XHMaooqnPOt
Lwhz6lZ74/P0EWesr3fh+jnxkGdEwNN0xTiw5yqGvmVtt++l2vW3JX8HqJW6VIqrSY5ChnyMKSI3
UVp+PgrzcKCloYDACT6qjjHzUypj+JWC9PsM/Kw5Fra0XKqMSNdfsYs9klxveKCkkzgk6gP8/fz3
+M3LIprq3LPldiRuX37xXQrHHsyV7aJU3WQu8mA67qbVJZlz96sfki7GpsDLMHHDLRBdnljIkUk9
lK84QinHJjylZgzL/m8h64lhY0qjWy9A3Fps0qk2FTF2SmicMl+nZezLV478lMN++SRdPp5QmE1q
EYovxXFsRc6mcJTVfVMefSyANqjFQFqUK7Xp5Kf3337lX/Ri8VUoJHQPkaxuyIslYP3bb/5Y5HjO
lm7cs+OizFwacvfydKyZRCWkwcX3k9s8/vLZi2kHBtDcj4kXhkgwawhcP2zWve0xDDmVYirVnsTX
6RtH422NeGuYoPR99vQ7RGPD5+ijDAwLX+gkusRdpPmAAEPOekUQO9DrTa1z0Ty5a6bD2xCmQBau
vycLLhTyVUHlGM2IbR6w779QhqxpKkKcU9Bgy/j/g/wOgyS0JAglRP+zCdX716uMZFgEWlfe2S+X
d1Wmj/YeH7KUhPycFY3OY1yBNIlYDNP2PaKGX3qcmv+f+hFXvzRVqSrIhX6+HZwpopqDp9p1I+IJ
RRETphZUCaDV4C76C5cd+2uLcd9dMnJB/E7ovxmSpVCFlF0HY7+b8XTlbXTfHT6n3yCR79UOrt7U
dxQADOsZ0kwopRQz4djNkX04/JWrrG2PR250p7TwGTE1DboVLfkn2Nsly5mmSWrBxAHTRGdOm0Ew
So9TEmLCFJpBgikbeCWybnr11/uZdtCyFYjzCfDcFaoec0GArZooTCro5gOhHJHO2VpQKUbFz6FO
uLsbDO/2knCt8sKE4BiUKmyhTP3igggoIZTOo8NjDEjQ6NgPDaNEGgQo6HF3QPVkicMkSlZMSJlL
OOGkYxx7lf0nUYxsujilhAFbAnGCDF5zPKRx8NPqZnuLj9ciQFjyitFLTK/Www6Rg9fWMa/+aBD2
aEMEba/YCSF93TcmpSDDYkTvi72YDsCkGw3iH/X78UGMlqJCnKz/8Wpg0Ufy/AOkBcQ5Tu+NNDvV
sXilzh9BV02LeJJeEIDPFKboufMwEAzjhGzdsuJ0lny9x8huCjhGexftbXoajIfxFMlt/cmBagZ0
lyKj3c3KQcK5PaykJmzky4XXin7PrfYuKJnhHN5VjqJAYO1KMALXsG6U3wuuIlNzKDHkm2IDiX9c
bUgQMWjXZIA5qY14O9QzBlAfgVsqJeWD16KkznrWF30b74QLj+lmfz1/1GDzcE6UgIohheYkO5E8
zIWJ8pwjr5nUd6eI8GIXfYKeOZgHGCZ/fPgO3NJg8LGGYI3gvUo6hsTCL7GHTuMLP77ZKvYdLroq
2Cz5S6f5zQuFIZwXBzuqeDfv0Q7WcjMSAQtBs/T7AgWa7N8ILa/n+BrmiIyJv8h7cEOWBBzZ3i/A
dvXm+NO5WLgQkXXUPnHcKqlnRwYt5vHRTVeR0puQiLbMe7MdR/8DYppruuyayoZP461E95vdrWOL
aq/A9HV3bEsaPBmb6bYMPEoYzMsCU0dZ+11CbAhtOZ2BMPaGiBv3sHh84J+9JCv/bqhwuOlNvL19
wCHstMzI6S7bIsdHYvQPS/eeu0at9Ufmk2bVHrvpN42k0MhWQk403chEf/71Vccr3HZcS0ONxdM2
gsWA943hhajq6NSu+ST+HgjQXc+5877XM4qpjBvQVqPyKHtIpV1VTEdZDaIKohV/IljG8hB+LGKw
+fQMYlPpABwWgQ5bhwMlZfYPepfK2MsWkD/ORf8o/7PEPSLgNiBxmbcNqUAbZnScMABR4RB35lAt
DxR4Mw18BpB7yii810pqpvdiI7GJ3MSpvrjl0395+cHx/1wHEHDo/FpGu5ctDlgLKwcOJCy2oObI
znjmdcEp3NyAhnNcFHl8qxbGKdW/X80HfhKp8Xe3JCl4OSqo99ZbK9J02FnkEOcoo5h49W4sYUf5
A5YhWdOmBe5p6NHBIY3CXLzJG+1nMs7+L3foiYXaVwiTkrtWhOg+wVWGdt/Id8Gl+ZXO20VsDSZd
zHEW0TEqz5HOwJugd0aNGmcgK3f7bgFoZSB6KmPsPOgkn9nxgUkleK7rICjP24HxryjcRa84Q52w
pVn0E3rTkqAKmnVyjwIQtQ8pXFND7I8YIKbgo+XytxFfeH3if6nQX2jqgaqc4Af2T17ZSRkXbXvx
YUCmWi3ZbamRDyPvUSR8acdDsBJyvbLANosS3sK3IZcxj5HR9kMaG27dY+GGXUVpsrBiPL+CiDsp
W4cjLpxV1pZ/3nD90FHITy4qGRSwVH8bbXgHqA9XSWD48ooXjv3JsYYxTcRnMDBS6vQmEOMLc36e
q1LUUuWbKIMBWtuCyn+hV/Mr9wPdx9c6LNdi7PkiOjo/5sIr3pvKNOCMUr9j3JmOiBnkdUk7wtfe
Y29ZlmVXoIiHwfozkyHw1ZTnNwrx23n0Lbok4daZWxCFKlExZf7mvKELqXpRSnttNYoiKHKi/nj4
V3NdvksiTiTOtsAwLUuNv2qB2hl9mzd3v8cKmPI7oYcoOMzJqzDxX9zEYnnnuosMYDubzWMgSXC4
+zvaRd3Zk+y95zd1aIQ+DxJ3tL+z+dGv3lDzLqdvlB6WfnujW1s+hJSWP3SyPHEJSahLIg0DFSuW
RIaKoLtw6B6M5HGB+KPNB2hNgFK3RYWjXvC5Ry0cS4vzrXEZ9oEo3/fyuUzklgJAwKBmoV/JK/qj
Z/ZAQH8iOSUVM45rFbYSmFM4o6SZXRRUuGnaTGkxdDEmPAv7zwPrz+NWIfUeMpRYKpYUmFl6012B
5hahARbIMcGOk5qrKWXP9njEyxrtT+dulnQDFR0ovsd5HaQKPZ8lT0HgcVpEQPHttk9rTgIAcCjQ
Q+TpINN78M3drLfgYOA0ULYkzI83IodYLapUusPbvaQ6eAeZKMRjmVurZrJpT0nvFpQStDPumg1E
EsrznSlBMDrf8QLXxwwKdfyzLkvw/DJYcCX5OgSb62Ky7eSCoxiDQ4sW3GpuOKpcKpO4C3EjxKVF
blg8kYhAnhsygr4LnhehK5h/fFaVwRMatQILKVIPsMfrbHS9HE/dqdYHIS6fylY0qHTgzFzSXV+M
EY9sTkFw5k/+HIlXnMAB71PP/olSZTqMV4HaAGr0ZwlDpGdFvzsWTRXT7TbIqlJycsgk9FP2wIpT
7xpXs8LWQG7RGQEtGPDdt5MSHvNykNRQd3Efm5bwOfcMIRatvAy8Kc05htbl5HYLExq3Dk+xV59k
wkfh4zbrOTTgC14rM7JGx2M/RLAA4NX5Nhx3tl/reCEzGcaZ14D9S0IGceWjiSoTBHK5b9YCnMRa
OpREjJ0T5aQHeFsJLj/ZwtrUWY9UKQMUVNZsoyVkcJgUtYLJfc1h8ZNQSZtdxDc7mRmH+/possYD
aIk1+tBo7SVTR7/Fx6B6iVBwQGXj9iD1+sIFBBmykI6BC9NHiQkEKskvEozRhWgxSI8dYpHWYha9
xiEkyYQMva8VZ17I4XpMM9l5NY+OEkFyjPv5nlYfaIOu7lEZDYO1xtq5042zydrErVF7Nrz5EsF4
3WxvJ+QmfP8xRoTGO3ypmIWXE8wCWzv/s4P6Qzwm20AHUnAQLJUSjGZ5VxLDPVgUxJc6ien94vqT
2NgigxG9/vftzZuWMgQijF2J7oWyR3mJ/xZWbiRVj0OlQROwQIkH/hK+eUIR4O9GOyResIMNDoH4
inp1ltcr1kX8MUrBhuXoTeMXmCzq/qPTh6i8kPfKLJ2bC0+3uOZZEr010Gy/SYgm9b48beMp3GxH
WxAc8UatcKTCRgSHd9RJYVneGEpJX/P4Fkms5+mOg8oKgBuT0cc3R37o+hxswgWXfo8tiieCaJCM
0EDuXWsF41muqE7MBpmIEDFoIH6yuQWWk1EOc1Crd5DVSM1aoZTLS8f+x3UyRWo6bwBDETuFtYPT
2Ia9rplcGJmYYLZWcy97RAyYHtppmoJakHU2/zjhEihhDxGjxVVzSGWaLQ5hPmgtYf3dVQeRcuvj
lomFpOvBrXg0yp9zxOAc21hQ2rr1jRgxfyyHr+zN2tMpFZiVwPhjGkhajzcJ4j65Hie13vnRxJ2N
wtXIEVrBoZ3udMm9C1nccjEs6WuOmPZ7zERLoHL+tFbVaCGbAVsIJ5eD/uJhQhUz13t60716JBe9
d8oU3GmB+yA/0ejNpmUCM6nrlxqaH0Gv1hA2gzQii+NIj+StCFj7wZ+pFpvI2JadYc/YNHp1pfMq
1qmJXIaY1a0OZZgCUmbK2MhCKWumrfpzgxcg611HcFS7mDuZBK53MBidn7ERMNKgr0Q9DyuJFOew
Am6cUG2OGJE7PJYDl1GN91fz0hp7y+rVT2Vi8N2KUw/EzixiATEMo3zQxlGDruZC/PEb/cTxEBa5
j3BAOZuDgvf7WXBukTRnL+ktEsdjKpLqPtct3Up+h07N1OIOX9P2qzyANwrGK4moAjrQgMXAqNjB
DpghLOrW1xwLGvM3dY6865QlYkHVfNIpBHGPbNk3R7f3lweqKrfQwzINNxYNZT//pfhiU7luOULX
DU12E0qEKxQZDjlJ/1/Px34kGjgX2fr+sUiPi3Ey9ZxEp71Vz4FHbJ/jjrBYuqdak9gPKEQmPy+w
HegXkF8Ynx1M7LkKdjnRi2S+oYez3m0y7hU4Kcduc242arEwfd4TAFH4oepgkjjB0aPWAp6S4Zmi
V05P8/SXyGgdrz9siEfnEe40GxnAvBZyjA1w+fe/NIlx2Ctvmclmx/LPg79b1zhQWmCFmzE5J1oG
MisNNdr1Zn/loc3gjez/mAIziPBFDSOPrnGX9J/BN0hP6mA1yKBUsbN3IgV34zMb0ozBk1aBTmiH
KCFklk/L+q20gKaurCHBxLA4TzgqBLLS/MRLAJRNoYwyVSovAQGHZGm1eP5D0klg8k8sgyZ/QBzE
dotYZzW4nKW+vWqLd30uJCp1Bg7qybwBOOZ0c6ualF8PJbrBOsT4qYhCu8Ut0bTGlNJezRa0bBTH
HzMf+JBmD1WU86f7gR6txnxcx5YK1yKuxCokQ1wpntAMCPIbq4S+KhdoZgJwEsGBZMFwP4RbBU1F
1u8yPDeeSdEsZqvjiibLIZRB7QyusJxmyJRgzfEZS4BLCK2b5BLBQ2p/xddQ3aJ/W97i1MnK41RR
ZuQJybD9cWcvQ6kBZilbO3lWD/VvCBAb9B6HmPcI1qxpOxI9edTc5eym70KTD+0YYANUzWpCRlKN
y46PBCrx+x54i/xN+0BFpMDA7BRsWnY+QWQc/plZtMSIQasMHrcRwEg0vS5oVL2UWb7ZgF6j4wjS
HfKtJYKREIBMbebhiKfjqRTdCgoCsvUb9JlZbs41ivB+IB5XKxWo6srWjgQUyxTTsQ83JOadftXr
O3PHtZarpANK/DuSnnzMritVMaz+3cP2LHoa4pRXAI7Oxvb9OF5x6G5Y8GFpinmJXZn0EVQAzP6b
WHWspvxO42K1YT+bIOej/qgG795I4Kc0A3DDogtEaua/5imkCevBI/xaG4P11kik8gJjPCdxzE6f
8GbUegclZZ6hUiqP16wFYCVxEtQKxLaTgLWK4BjNhaFq8oBumW/vjXZM2TE/kroi3Tj1YrhkeAeF
eyMyKJX+Uic9mONhlG8EkeSsP6jVk4dGbp5HY0P+vVhvO69NjrMNCEc1ZxVJx/V8pF+LZh4XDuZA
DNRI29CppP9XXZIblGRWDqpsAI2E/dNRw3j1b3prpsS7vCWrMVOUpvBKAdRVgxEZ6lcb7MGrGKDB
O8rv2wdaWkhVzi3xbdqYs0P9so0T3rRe+ILdPH+D3n0EywhYKcm3UJUnJsAYzBG42ldkzvG0f4DR
pAfQ2f7nyV1QzEW+UFvfwIzqSNe8cN7mhT8KK0ajcGn4xBb280BoRmTcrcQZ/4Q6rmAc4uU9QcZP
mwSEqAlcgUllGquBNb8pJ95/ZE2YPaHPV+8VBApKgi6oulkTC0Prk69Nd4Tz1PrDn5nuX8rbc+2m
GiZV08Y2wqva6ggFKK4OG+Q/kwFtMIlidp7hS2+k6Kef1/copcBixaqTVH1SMkvGAK1NgmfcMi13
AR+sjR9RslkSxArnXosd5JA1tADxV0mxEENRavtXklxfbbxp9EmnZT3n6i/cNXCK81bidUXmLbZm
o1cyHIDahA1qLiWMAgaSQdUvh/1qQW7X2ENiNEWfzInp3b/XXdxPkxGenf/OgK+J2fd5va6qY23E
U5gCAMs/ud8LKQ2R2LpqNAhMKOPuu9lNnhh/r52Otj0a9281Pavjjsu9+GXtc/zTYLePQaenkh1R
4X7kWUtljip/Zrn+o5I/jqKZN4YLErHd01GAViqEZaPcklk7vE05bZ+oSch65G/j4mJD/TOcrIcA
BRotaNuaYN6gxdjBwt8JiZtGrgDelbNHBJmhjOZa0itGIR8lrlbEVwLHhWTf8i2T2Ia2Lysu1vBi
B7oRh3lBXvDlEiGctLvXF+ukas8V1m7Dwcu9ywn7+zmOmhy+GKLJNPhG4STtPWrvKwOTK6yxTIMO
2MmqTMub97DACsE32GSydSJVZeB1f3UsLfWAd8NhycKPRbGzzNyD+2Pu081Ks+qU+YIMyNc1jbPu
lJskOpDOj0SfXIWHBGP9Ydh87j32EeVdbuFx6llvYleJ/3Z7P1AshcFPnwR6M7/QJlp5WLw87Xli
2/wtOSWYyFoWSm1m5fOY7pKEAjGLHzAr5/yQKFifGHm65qVoeiETF6k1xf6USTujz+rtuPDzchSU
kics0dllh1+Rd8EGugQN0wtEzIAYH5JB/ZWlhRx6xbrB3xF/K/fT9248Zcz5T8u847k+oueqFrdr
7wV7yR+9BSPKI46FVF+ZyFo97L5ndNzDjmpA4HSMwG4+d0MIKkzHx12nSizmTOw9XbID+5V8btJE
0ez395Y+Ah3Wc8LtmsUDIwWMxNNDLzgC0je6bbIkWHVzFpsHvysubqft5PaiDe3Poq+OIL+ZW5ph
8VKIxnkSvv5+AqKCAMDHXtTnTM6CZa2reZsHuQNKgqYyuRks93TQ3rmjXuBvNVuxuicTB34lwZPv
KhbeJ7ufrQvsxs9ryDtJKu4y//rJC2NPe+++/KOgbn4V7GDhXc8g6LAHHnxBp72nXT70sDzDMTuz
T4swVnOaAnJEY43Q6KZ9XvKLAXVzzr3Uzv3k5fo/IrB9v+f3Pr+DQQzTMbgYBFLAa0jaAUmBUX9n
iCoGiCEYlIF7u/4AL+JYOVJbqIZBiPAw3jL0z/ILsUW8+vsqzUX72ZNh0oVy4UvJCkMLNXUcU2Y4
8JHKfTY3gQCB4K9MlM+NknVTdie3FwUFdz0ztRKRJuSHUoaA2j9l4TxwzJ2YZ3SsSfKwf/QsEG7r
I7wBr4OlTihyUPaGL1Gq7XyIcuLT8wu2O0BkBc2FktelrCr/mGVuJZcodrx1W1zezk8IOJANEE0t
dlHsfpzg6QjzQL4XrCyB2soc/GxztdMVk4BxVO82lIB7iSPDqg/VLIjuYRrtDfRsITWlRY4FywiM
JBKxAfFAy32uw8NbBnipEoHupTM5Ytpi9i2cb3PzyDlhPQl0EuPKWPYw8tUWzG/JysSsLhqnP+Zm
ZhNteG27dDES0wAGAJo/voEihDNes3emJh7mi3dDIYENsKgoV8uIV+CpseJnsru9ctGzMW0Ayveg
YosGSepd0F2ZfnvLt7LJbjlmqaunF9bC4CGa8QXusW2qQMN5gzJz8kEMaAwwRTfPGJoCNg5uFfVz
xeambbdpbjcOB/8VVteu0puIKnzJkvQSNxiGcw0ULK67ikfYm/UHQ7lETeIJ+Yzv2FonFgB564Wi
N3Jro3psLF0wKbqlZyAemra3Tyh/Nk/3/8SpGSRGHxj7SJX6cwjzjxh8mf9Ahpj6/uALwzMNszfA
EovSXuaK5SriDZ40G/ab05NGASslSqbzVgbrD7kPu7oeXPpY95TB1ssLlPA/qSMepn+2J/Q6eGGA
okKCf8JgFroaP638lkqVEqflZ2T6/X3ppbSQy67kfdDg0YOVtWoeTCMa6vP2Axqn7BITTG/fUAOZ
Itj/24+Fzsr5+Oyf6MpVag1nIUWI8ptt/9GB0qEafER4DEoz8ytJOgsXQfCK8DOek5ez9A3VLlsk
C7NSUgEHHvXz8/yrgGW+ifZBtRUHPKGlNQsvaVIY5VrWHFmEIE9c06i/Lk9WVOvNOMBWLVzCldpw
YJYPe6MnXzej9r+7yfntCWu01IDyIxzS7HHtIP7Uf/g7uEL2xNNxwVkg4N59jVZv4RhkhW+v2itm
8SlCt/yR+WUiy6cCEn2KXltr4FLkxJiisTJZWh+dRjqCA3ZMxUGA5MBLnbUEvns3F8QqvUdVWji3
LS3WT0b/m5+Ij64AwPhi+1TaB8f8CLrJs9Y2xckV80M0mhLeP5n0iPnjaI/AHwZkRrOrybftxwHs
gbyTe82UW6aySNd+4cC/W5CijrxmgzQDFIOts0lOoz8jCvRdRLORneXbNSNRxhR6McjHS06S32fR
N43paMqRVdmGRF57TmEART0eWEdsCQIpWcyZBBrsfuTdR9u7ENUq54jG6qqH3/c46Se39fJ2qJn1
NOfzyMfd31kOnPfbVkXlvk8llX5zUTnyaabKIboxkWodLKepWNoL69SagprRsCL8PlIQqXnVWNjZ
k+suCzA4Ur2y/S5g2zoO9HK2uz/9IddXXsF1ZfsdjH03YAjWyHlt/YJCDwPsL2+B9fVJBEFNTBPO
5DVKc34JUR/Rb+e2guFrGH+ZOGhZGkcgoKa9QLyp84TsmeyZnyLs6Q+BXE1qLCH2mRH4e/1/3Psb
AtWDxMrYPkyD0x4tl0JhsAjrVHPTWFe7HGDWAq6VarAxGgR91qO41UNQzoZq0whzLWiB3ojlPxDw
taRMPjpK1Vt75/A47DRuokErstiYqMtCi6Toxn7ecmvgRSw8PlH8ISAbLtNU0oDw9e9y4luo6YXD
HJ36UhvdK17phPQAGCAWsVOpDgElXnXatEVISOdyCB45hKEeUUZIN8G58md7wm1uuKzE/dQ9QU6C
ZyDvyPVPuAgZ/BBtJzSPkjuo9VJdxCOXRdCiu81sTCKSB5ilzKBG/6e37nKBGykiT7b+LxoCXfyd
iB+avvouJZQksXUzp9sWyTmOfGgVfBMf1dPCczFfNWnSBJsIkRMH5jU8wn1BQQQuyKCL7k+FQpDd
vl/vo+byylptXMfvYHyJVa3jBAPtRJHJ1alx+dvR8dfJJ3vlilB0dOgjpTwLAr7umNLjL4Y4M7ep
3A8ElX4pkmHt9OEjmqZ75FazB2ga+XmOwrRPYgOAeU+7PsOFTlHpgpFRbFz52BQY22ZDrlR//GAe
nH1vnfOLYdz5eSfF2x/I7b7X32K6M3CRxjR/w6tj/t6ZdlzJACHkkCBsRjDq1ivm3SZf6bAZND7R
SZF5h8PELUhSv61B7rAOeTJGnSrL0UmEtWt2zHLob6wK1f78VXdPBuUhgcTm9ck0hmKKgM/iTJ3S
twg9SX7zLKYnUqO3bFazbA834A90ID2fzxbhc1oSi6SWgcttCNnJ1sHZXIZo6BMBoZtLeQgtms9w
SiHw8PVLPu0IItF7IhA3zOfhfOT6A7uQmD/9TB6g9/8kt3wqe1YWv19gomyr8aQJotMuqdlXVqFN
OjsA/32ODn61nlbHOva7C1dsFCQ2XZjekybkmSVmlUdZuMWZJEGvUcBueBps6Cv3Y/yZ3S1gAH4v
kP5zIUs9dnLwN4/GpJVi/tqRP5aSDsg/XDDfSWaTTB5QzPE1rwJNZKP9oYLQgQC6/B4rDRD6TWJE
THlOz2ocCneXMNyVYzzWXbn+YRp+7gPv/5RDOJiS6Cjdg9bOOYOogZMvQw9UT85XyKDabazUZFNC
gKrb92KYE/SFs1D39NbynNjWDsnlGbjCZlTtGSIlaVitboE4yf3h1q9JMLTfpW1JS3l/IfTWqygw
g/6KlNKnoiWy6eeKE4AWAclPsbBWeZHIKICXYQcQ5shxUd3kbstPhfilrImgPeJfjZDpm/IMdeqC
AKScCcD/RYoOxKX620julupr6XeSfXEKEboomPLSU2aOZRfXLSbnAYWfycuO5YWQ4Ej6IUnMSH03
h+xVJ6VXjYMZ4KMtvR8ssCdCdJb/KcLpFrfYRZKKXokhWhEBoZHcgp4JwWp08JqaWu/Sb80sF1Km
/vE5zocJ2s8Il9JUmOm8iftjN12OLXno9HWlKft63dmcgQWQMkpmZy2YB2uup3rzzby4nTvSsQvb
+W6u50y5VcAx6vVxWgec5Q0yWLWbupSKYQI9GAeiL82WAROZRTGczdWi78wfsoHFhMdUohjJWbQW
Vx1dGEhbjOgNeTTs6sMBa6xojnxZ9nSqmU33/1FsKiDL7DnqHtqdIjcLT7s0cb9jAV6Q/69qQasV
DkzUuQCJttpWYq2j4Sa/Q25LFcZvX7CVuyz4Jtv7aVTGOaZJi8NxkdKz8ko44HeI0ZFd1OUGy+Ow
X455L3rwpGZRJpIR9RaJey1SBQUk4cxxl3/teE7fU6/Ub9KjhGmfdTyXAxgTuxTBcuG1Em1lc8Fl
3Ngg3J8a6jCXLnjOgn7NSRc6d987JQwuKGNPnpnS/20gDBP5PnpjGrjc14fNPoSUuJ8JuBHEpIaB
BJ842jy37MCtSyM4ilq3Smq+L5kw3Xig9tSJdWiRDRSh5735k/denChQKQAUCfToPJch+yWgs8hd
zYRDrX26QON70ZuPS+eEN5W2tYAYRPlfqrAOv89dC5+K1np3RZuM2Vye8lbrdSEjjnV7prfs4Qig
5q3lAsbXxD+fdyGs27n9SgyLmUT2b7Z8+Quz0ICXhPGLUQxNnXUH3Tft9DK1OWmYigFdutqFdjQs
MCdP2SMhbXWwS7LEMkLB6aDyB5li0nWGcXwOrbjf2UfbTz1z2kj1exGI4V9v/QF3nvEez1yA/ZM/
2cz/2KlBu1cCtbf1vzOR8XXYFLv3ELgaTjUZ3pMgEjZZXrxW4wldLD89pwT2ug8M8+57vsS09pxk
FZ6k9mSYvBbg0FjWGl9z9wwwOyzcr6nvw6ig/2M+STnYwNBhPNZ2Jre2Bkpi/x+SU/ywDUbmHz/I
ItGRlipTWspHk8+lSi+sYcN2z44KarHWsKeg6NdBdMecE5MtahWS4YVGDCG0ceT6B3u7uqSCG9o/
VmGluKEUUd/lXSH/qsy0SymO3Vp/Y8WbLAo6BI5NOjf1QKNcqR9zGpDLhrrfiobVp3l6dirfdrI4
034KqEq6YFg+LL3V5XaVJiZT1BPo4R1TORrXJFTGnA/j2Pys0lpWR/E0wrXjAnH5NoDvVxNxYw9w
RlaWO5OjEjAwE/NZYUkZF4AcHesXs1gNS5SclSWBbG1/PvJZLxszc6C0czTVXtrRPm1yV1atpKh2
hT1eyJ6DRNmai0mGyDNg45JvelYsnpiAmDkfzpXtS9gmix7gjeZXu3S7xxSgbmoDbokf+Me639fe
CtfwHKFoNRfCqJrMSyfIGhQF8/5F5aZjoGNn/N7S0ICIBvyeLIiP1Er20Rv83jkffdhtS+hFHE0w
SEgeCjPA1i79DHT1wi+tFQSaTHd22nTyFcRwQoLLQFKC5c7Xihil9o5UcPA3nqZ2o9jS2Mv50swW
VXWZHOxwws2zL7GpaAma0keckFkzVYTqxSFH4EIsVArgMKEHu86ZRC50lMArGqLnbrM+djbYNUfJ
G2K9Q7LsSHdCZXPdKIab6vvM0jMIjKWOfHlkZdSS4/94w4xNO2DeHVVOni9dH2tQ6UUXKNr8Jq/L
vv0GUDHd/dN+ZmpIjgbriXZ+vzqm7RqrVAkOXmQCUlCJw5UnG7eN0ahj7czE7zhf7DPIkil6bRBs
7Me/eZa/rv3pnn29dPWHmoorpvOFSR2hrfShQ8xTRSHgUBxHkU7Xr4zpELXwEY61YjK6pqlDLeVY
qZ+PCK5cQHlp3OsnYCv+d3JFs0gzfpDqNmcrlWOq3/QDhGzyVmZLllmLdFBck9SKRLef3rOmEaES
z+SX0LxslSptLqsEvIEaAZQNPIPp85qqkr4e3vmZvRBs294FCKT3ipewsMt6AHpGrT3iqLndFJat
Zn9D7e9MC1HLJI4E0G4AXxbW/uk+YF4D77COp6WVZA5rH7jhoZXGV76WnVEz5UY2kQ78rwf9/HgK
1TMCPJiAgx3B9i3+ODBVqmyiAVtxJMZ3ytGo+5oTuE+Qwa1vZxRGFXmW72XcaKZdbKm+rm5Mx0CP
Kwx0W78nsrw2UPlZBZXH4AGQpBRHH2rf0phZ86OsQwTQy9g/wqOhK3gH1zAwrMh5NOP7AgT0WLiy
fLYOGdgR1JyPEvr7M+uIAfKR7iCtpYRG9Ce2Dcv1s9IOdjwqoSGT+gLTRY7/ysr9gaLWnMpSZ4Hl
TwWa6dVDil2CeoSRS2XhIIQfMt5m1x9AM69WOsiGpSnh/KdD6k5TlxRt2usgwZFJlRf7YMtSZy2M
x4QcbNNFpnwGkNG9EHSlhIfIW3CrvTG52D9Df4HLTttDKatovItkjLXDRsR7nvq1QWNxceoOB080
J14ZjvZOEg9Ekf5rk++uWvHGwUMU1dNgAuSHIl/53Mt2HqML2GrFDca/dDN9of+RO1fHFsC2/AXQ
vensOZLEcWGutU08nJAZiQFH/xaSIC5PSo8gtdVMACRC3ZrqHJBNj/KkKXU51RE8oFfPDqRHgtTr
MER8mKILZn5KFMQj6XiIiSKpUDDIGWCgpmR/U3h90W9CML2EDTYXKLC74BCdC4e+HoymHmxx2wvz
FshI8VattP7mUNGwhbg+FlaE0xbiPoV6c2soMzyOx6GsAQlomgavcdj2+lnM64Y8A4KKd3tnWb3+
4ELOTZV+CftuUqaD3QZTlD8Ps0xwgpO2YC2qhC3GuxasvWm1zXjiu4pYKpPZzgomJ45E0G7Mwlh/
4fB4E9yy32lnyTkPfV4cnkJOPbFrLwzMAX/wXTpZqyfyJ9jILMQNPGmQqg2aWwQg7KXqt4VEz8pt
5OxYvpxysEfMHtX4bgTAdN/MfmyP0mmHbGtiIL/cq34ETb4nUDCvOgVRlLYgHtFc6DqwBRjFKaW1
BXgRYbiFzKzD0DHBWWChFMRDYuWAcdvE1YtfLHXtLk1o8Yih4ra0UsAJ2D+isQ4ZHnnmPIaWPRE1
LwcWhoE8R4/eVrs6M4Tbt0UcbuN02EU2ZYukgXjydRHE8N0+aJ1BNPYHW/tsXV7WZPkFaJ/9b08l
ILpwaoyo1wvyylqyKUhnNiHKh0u+EzBVQPOLgsRe8D1CSCnbUL60Xsm4hwwuQ3EM/wBSfgKOWmv7
GhdLj23qa4bE0xUiX859IAST33GMFpNXSkO70hQUL5RJnStZDEldmX2bMWYFv4NkthnSHs340aip
85v2WKxcILnJVwG5GZ6hbSIjHIRvBVC3atfBZGEL2iRCNWaLeCX+FARweIQj+f6LUnZXpkDPzK8/
+ew7wPCGyJ2gNdkKhnMXMhPyymvaKLncWy4xWHVuMmKUUF5BDBtB67wawvSXA78baDstsgjXvoyb
+UASinHToOBvKfDSK0gK9+OAFI9FKsf1ES5iL/tPFAUWZMrHeiL1pE7GoKoJuLNDu3rlae/gco8B
iW6EcLi5gKNWGztJ2fWOaqHgGaaFDzn3x980nwEPqlbUUFOAGDmAB53rPqA/su5y7vbVH17DcwSr
y0RMdkw6sJ4z92ks7fbwMVbP2foSPWFD6X2H01l49UjHEl4c76i87vc2Sr/XJ7cDEc4gOuJ9eXq+
VKmiJuw43NNTVIbKkuwksEWllJjCZqF9xhbSQ/Pe3677lxEOwSSw47y5AVAObmGi5G89ITSpzezQ
NzOT2lz+z8eqXY5q+HT0+VVEAk6ZfaOnzhZuZ4a0TpVRkbJzqUjcuaHvbhbyLTDuhPB7Hcbb75SN
EM4q3zfFisNr/zc7/ln+98Dm4GhSghtj2wcEsePLQDjaZXRudzfQWzZ+aYgslzmW7Xg0u5+yh0GM
cHFzhG5cXbDjnw0UrcKGeZwzri+w8NZAk03Jc6mffwb87AeIH/yuaWgIcxJz8Kx6066Nl3iuO0UQ
rUbV+Uh5wzLr/vTjtXyJymuhVCsyeo00d5XyiVTX7lDr/x30lOdKWaTfR4/REh2BtHnOOcqkSE6Y
bEuCLxB6B/LBZFROwPSgrjeyHFQhUazAbaqzkSSaMjoogachVCess47pIr+Ng+xZg5HPAubfA7zr
Yy/zrzH2Qhl9kew0ampFza8W0IIHayRd3VRdIQ+Q406VpJnP06ySufYzLrCt5rB0XwdSPZbv0GqD
owxpYUqr4cw7l4idIrx1bCzaswgQzVIr/SoyB8SN2EuQTX/X86zsVUSlWKLJhFhG5zkRmPnp04XW
VvTv7H7yGcavEU+0IePj592OVuufvQA8IFR3tzMwKEfuOIMgkRX2rrWUUnRxIUdinWkzGfTsTpNF
bSZa+5hUlQ7yq+6eBfdidLH8jdEN+9CxKzUgsky2l0h4it6rsDcQGnylCMQDn075+G/bCLBWnxYm
HeGLOhpueHngZ/weA8Uyfn+tcJKjQ0tISI7DEQ3tbO23NNU4AptQ37J2jDg+wIWbCsDaSyyvpMNV
qQaMiL1nrK0h+uwTY31MKgJBdvON8oKCXhX33Ynw9mwbDmW/iiuxytkWTVmgGfdDl1e/Eefdm24i
86QDi/dU4Kt/HEgWBgQBwZTfB0YMV96gfXJfuoIxmjy9lPXesOyuI9iMGCe6AMjpmTcBeCiA+aaV
1b7XdjEtSOcDzSAhIuqsHowxHGCHCgjE5qjdCrC9G5flQ9q+37dJJWJbKZ1w1w6nmtgc4k5pK2fB
5WO8Rb/QywoVWczp5rU+6fV+fJDMv86v+PMrtNJiZ6YqHxm9DGTLIkgHrMe+bBOXcgwcNXhw8qn2
JFaYpQ1sz7+aDuNLOqphr6xI9GN/nQME0sRROb8agDSXOIjQ8Cl5JP7HHEJQvEiIDGzpRzRLcXpP
1xlC5/7aaurHfWJiGdcb0gZTO5KXvqP8B5dF+aVHfbNK7XlAZ8MBVegdD90Q6gCL1YRBDOp9d+Ap
ZLlJwAaXTwoHYs1R0ifHh//Lu2M35gsuF6V6xTiuxGJMFcsv8D4XCOGlbhzDzbF/pXT94l2PG1T6
BfBQDR+GwXeNb3befbZhOyew9ynA+b0tAp4MsZdPpXnmg9CO2j3xi6zJnLoQ2UN2mobktlXJLknn
tnPZkAHM3cFp27zz+Y8xhi+fXzaBWKAnQvIBHnuTI6w47nhnA4YjQAJjMCaR2ypHB01f15uRRQyX
g3/Xv2+tMIxTpKCb4n12vnLi0LzVvHLmimKp3iMngidPue1LJfklDjgIu45VxuP5MRj/W7WwbYJs
uZM1O3I37nQztiBodAu+tIRmt8dhQvvNQk6fxYeGwEAgWUQ7mxqiRkybANGObL+uh+om7ayn7xV4
0TGFx5UtzbS2qqc4gIb/dF6vqSpUZDug7gAuXdH+XGcXw6Mggb+cm26OBtaLwDSoeGCmfiN1vBwY
H6hkUKzMKmFc8J6mybJtXn897uCcMg5LAsAqQ3IA15viXznB+IHUF7MEf0OFnT0BM55VaLBXBs06
m9WyOwWaCnQOz0gwyzvsvgj3Xv3wt162oDvfnWEAPc3zkP9NlQoqMdagTiv5gC+brNty83ViA9KO
l9m/JrwUZYO89Oe6mabcwQune9GFRtsEkyknX65z2w6KJs1mdyFZnuXgaVhXWY63Ho6gCfSOeSH8
BIU93fSorsRW/Cy1+4z65tdJ0nBVX5xU8aHhLk2uSIVsNj7EBbqCBnGKjd5s/RdV01gvr7rPXseC
ByDP1bj0asAgHI8K5s2Tp1GKajvCY7hWfWnmGmEstmX6/SVP34/L5XDzdocXSqKbGhj8TKZK5c35
vRlVgX3L4fCfBIP4wCB9pGSuO/w/+6RJq1ft458VlhbjFiXvZ03+50tC0ippTImBCC87pi2tATuu
W8SsMJdp4WCKk3W3f/RIUhBQW1ExJw15SRiQJixn7R4tkrTOfTJKDYKAkUfH+BV2pTy3ja0Ps/eB
utqQR3BWgSLPhQWYt/gAvJMhcV/SMYFy/tnOI7Xo5HSSYjBCw5MeF9xYiKywE8bkr0x8cC7N2uk/
i5IIFgIGnLd0+oPD7MCEpj9/OfQg6OkcwLC4/zt2teAx5vdRZyG/0CHhsH0P75/dQYhxCL8jv2Y7
VHwatMA2BMtDRkl41BDJGtopBg8VJCy2X4g5+0b1t35K6fZIXXf571eyntPm+4vmXJ0Zg+CYMcpu
7K7i3WAh42yW8wsJN8NN8CnfE6VXI4eVbRwlWbhk7QNlASqwbXz2Q4JKruIwN0SqHOg+LOElqdBR
5RvTVetxgxa5/AxLKM1t25jlQgisp+S7EnLauN7XETehwTVWZ9oqfTxHntYeTRdvfpyNMllD5zoU
S+ankUdqNgZdnzJnLB9RiV64tyARXZvNwBPZ3VhCYgBa9uii7nHhZByqw98mtThku0FY3rjyWY/g
T2KbVmNpd63whTYhjFWcFyOIPZ0LonNIeygTB+ylal500m+oLakHz4I0SRJV2BcIkUEVvqK/MlNp
CRM44vM4QP6/35nJ8gBXJUY4+jQfcRX5kZLQ+44xVwmcuusquhbTWI3RI05x3dh4V61wcBTetJuX
v5y3FAOs/6gBb8FtBCmGo2zdE+kdOFo6aulsZLBU07Zit9jjHTskpMSUhbl+jJ1w2216qVka+U8p
DEUv+/LRqutia75q2ctBTQI1mggc4WJkHYzFBPMI/qUIU0z65wYdxTii2hAeFLB58Hcujqv+bPzL
82Htmn1FEMT4jyc3xtFd7DQ8oMbSz9fvSw/cmT1+Ogk/iYi2spNIxo3LFGSvIDjXlzGHZGaWU4Zo
na82HUmZLIyk+txtF8rg+/p5hg6qX59GkLXSijVGR80NByeQGnb+5BPNsIrXrc+zza+p3cX6OzHU
4dQ/JxGbtMG0YixlYK7RktRXHe7xg9HKbog1IChq30hCE7ur/KIPqh7jut9cvV9I72fUXWbcuwV1
yKwk9LQ8MH80yitVIfBGu36LZVLQzcSG1exTzZM+2x6rZyOIkEbwHlVApuA/MlhOzzmqfVp1CoDv
y7uJFmN48gVm5olcE8J5+bZ6c+V3NuAEGaOSL5RbgmJ803yLvpxKIxUtcVbJyvIrLUWNfJxFSuna
fx5aiVdP9QiIDW/eo6gEuWXX0hyhxv7n4Mw93H907YSj6NVnmF+COoCiOOv+FbTyNYKY+h5HPzkm
sAkaXXC111TfH1WLtiRxhDcx/XAwoGT8eZd17Tgn4oEfQW4W/bW78XrFmOlhjuchn8Mp47rL2WCb
9ndkc9KUQ3l3HI8TVAZt8+pnAAi0Cq2VM7irRR7XbILXf3dOd0UVE1cHoc7AnXlCpWtYsSnUboSP
QHmizp+wge35oWJY/7Q2nrKs5CaHpjaEtaDvbmEklCynnim8R+6ncz/M5GCbviw6w63ZRYEC4E5b
wswhs9CPQLp2ondF36VQTwxxnImDQ+y9Z4rMfOvlrdqzkgahVDJNi3QXwBnf6saSXLRDYGCYdxTT
sBeFF9P+YyHay5VFYrlzOM9p9Sd5riNntgeYhVBh8iaJ1GS2Pc26z486KOneyDVK/jqglbjLe1iO
VlSKlsUMICrKxsvPAQM5TG6iNNUaLKpJrYsAZ6qJ79TRb/6QROzy9LkUD79C/4i2vHeSqH0lCjUF
FUih69UgFJuwlMqPWhc9ChYrluBrInSsIlGPsyRxsYXXztD5XxqO/W2PJmCNLUzeQ4fa2QMvQBTj
dKnHHbETSqYYSXarZ5a3NskeJMGIAqPU8zINGHPQN4IXDORwTtVWLUhsr8rViEjO64QckEsdV6N/
gE+w8do0UOHcA8NFgF+UyeLLIYqNXa4P2LCdd179owV/V0VSJCyJgmjUSZbq9EVXMzP0OMh95xzk
ELwxkKswXDLFid93FgumEMWagu2VVondUU98SEYXxBq24Lt0QcaY5P0/Jti3csO+vte9r1gLWtM+
lcB9OSoo7UFidk8ehaZwc7FLQum3R0xk1ICYy76gFA4f3SGzd7odcyApwv4y/IeH2R/s8KRD34OZ
O0hnZsuR2/pT/a5CS0BZVMYdw2NUUoD2V++B7mf7wTWlP28ggp6pS8Jm994462RetjLSNT+8FY1k
ugbDkNwF3dcP3klTdhQokcheqzHCkyO0t2/6z23Dqb4h5rYhn/sohEZsX+7UWXof3Okg1EQdkiiX
WKeFMO6M7qptdH41Zd8WrqLlaUh4EvZG5cIAsWHN4vnactzjfiHzjfuW22heRrwto322iILiUav+
RPNR2cyZBDyunkJkdfEcuXx1pSSYORT8inHELyjuSgaTW442uYhX4LFNp/OGjT+PZ5klzwwoVDMF
RtcqL2dSaAQ869k+4H4RvBky6WQ8kWLOKbBXEnbJq0fVQ2rncfr6cMvCS8jG3/lgqYqNI5rnvPZM
76+Uw19wqk+TnoKWgIUIU/zlq+JRS0raJt8cY6L7uBY9C2Rqc7OuD9PACbEL8+hLtkSGs3r9yyO+
EfARwr1RDgI3U4GVN7uEEGKo0jieGQlkVisO4fvt6CLJzMNcZf1i8L3/plIMqOjOIXB/TuhYlE/g
3MOEdF53XD2A9YP/Hf3+L36LpnWcFLOCJVbxnlAFW+zVw3j/7qPoFlJvQH+MECWh5b4+baWB4dJm
U8cGo4V5zpzKMranF1K+kAZn/isL/879x2O6Mr81C40tQUQFyKWb24uROxlQqxg0tYNDise/yR02
Tc71NfCC9KamEJvw6ClkKO66LJN9/BK5H71pJqBciqxd0w0BcPQgbnCagb0Xr+lCagF0IlH5xkWJ
dwYPHH6bEyNnXbUz5MZcJJ1iZxkI+M5vyyTQSQcqCe9Y4Tx2zcHxc71NnTrp5wezkWwvPzcAeTS9
AjJ4jeoiUMIgk2w9us3B79Y+67kKmMDRCKFf/bzAxA45mwXgJh9Zet8YkKiGsphI7nXPMKVcxaDA
JlZQt3R/M2v3O/d1VDfTRepyd/Jo/Q5UwKtLE8wFMRoISnCHXA4C6V5yDOV4Bo48NeUvG8mofLOp
TI/I9poPsGpx0ZjoieoC7CtR1qO1+ReB6Z4eZccI+TCKK4V2V+2A2qsgG7/l3KoRQ1pKiHVD9IZP
CVu3L9h9w3WoSekYvQU+O7DgDu/VhSAC7ossBF8B5n8AJNpMQCVUIobkZCpeXHPgw778ITxR0/Bu
+SkujeNRspcqU1777+p0gMUhXUvltU010ud6ckv/Sgqzww8aaTTWCOIY44nKgOvFb8NaWmZGaOCy
s1veN3K+GXOUXN58w5zx3YZrW5MOAm+K/YSvJWpo6jpcjOCFHCLEm/wF9y97arLKy1dIs/ysHrkc
JgvQJtX07TQTXresbCzGqnpPnmw0qaFn7PqA/M9v3OSv36RoxLhDZ4EnQCNaOIV3KQq1fu7CcySD
Ug8Z5cCsZYkLtWAn46y+kJaKqLnioFv2YfgZzoVzhxrOMSetZnLO1Hdgd+AGGTI7sGSx5+xbtAJ4
C51OaIqP4NwimWdWlFBsyT0Z8DgAZReWSd0LCaATkifautjszjdzt7K/ybBmETKVyuHViSKacm9m
aWNrJbtA5fySLyK80l1wE0yuDrFxjYhFbcMdFmMIKvo+o0RYH6j0h1qKEYxMzJ1yBmiEPr22e9Nz
aLDRYohpZ7J5AuBXL62FhH6eLJAZ0Oyqhj8+C7w7rO8+MP8LurzZS/LPku7oJe7LV96je0KzDCQB
RfFPupEZQl0SM314XBF5Zyy2KHPYGjUt+2Ysxjg/9fXvvVRwIBYzMucM3GH/t0QidgeyEd3PdtdU
XznAWz4KGAHD3h+dl36o7EFGrphyd3RQELNaY00NVleY6Qyp/TcVxHuMiAX1VtcjjSFjNY1Spivz
mztxqTwvGZ8Ekp0n2KJ0mXilv0IXQiTed4VK2YEtXTsbihfuO9sdPCwDHWk5Pgi6XMHx4JpooJT6
zNiStnRWzkY2AaLTl9++oSiO6yk6+b5lBaHI0WQd+obQbvrA9VStCKPAgAl3kcxfcW9iEEA3iJxA
49b/Mat+R7pR7/z+LCUHTJ9/rMR0LRhZBU+rZLUhfegmU6uHi1nDXGkQAricopisuhWgo8Sg8X5R
X3iCFwHAOzlFKx48OpOekixlCU85lMJohzx58Qoj+91EpkldDQ702SLv0OohhREoXYI18VRomP1O
ctQWZtV/pC5zvq3cISFyS0vEIRLF/E6/cZ5blmhKbHm/nG7GmLt4pVORJ68E1BaYW9AW4MC7FLIu
1BiXsJha1boG8kMqIetGZrnox7zf6V1QKHjWsulU3C9+K7sCYDe4lnqvfyg+amwvErim/Qu39thx
YgmShGzkJKBNzMVpmk9k+q9u7CRejao5mDAeJXPAohub4hIHrB6KXBQiNRbn4+DiVu+BMYSeXFCi
12CJOJ414JoEntQVviVEcE6Z+1puAQNQUuYvnsVCY0wHIuHAx7EwZiWOpAlJXylp0ZlO1wPjMseC
w5Ux7ZiXNzRloz1Grhyh1Msnyk6dO3n87/DF1SxFRKn0t1HzZ29Tf0GelT8Tjpsbs/gKoTQGcozD
bT8AOc0j6/IACGjf8ISVoF4T8gMjNEjInQ36NwRANV9+NPVKLarLQwBF5UTv7KXb+VJXjHkgxvCE
Fm+z/VJw/ehfp7sqL7Je/smEK7qmlRgo7QNPko7RNJmsf/BkwxEcQxkCwasOS8nw3KyKWP6MPBBX
dZs3sseA6/H5G++okMoq5UGSm8Tl5OomkETGJ+S/94T9WsrIyWJUlVFgs0Q+5X94ZfGRk0yoaabb
VEPLT7ylWVOicnmO5ff4BAAE2PzGbEpz3x224t5Cy4/P6yIC3tnbGsMr61st4ls+CYaFXsVXBbIF
TosD00TfGYz3H0o/TvZImaUGQSVKh9XDkE97LRRTmqb8zDXq0/GjhO3J2lUqAFJ7zvA7srIYu9b/
qTQ311lIlnjQL40gdGVEOZouZkhBTQ9BhBhNrFKDD5q/humSnaX6jYYAXBKVDSXicGbbWoYg7K4v
eD08qgFEa/b+/pAOLAoFqr/H5rXngM90riVike5SUZXxaQR0lK3Z7n28AiI9Vrj11DQ/criGAsS1
nYBeXLGiqbsVI8SFVAeM9FK/8Zg/XoEsiWIeAFSd/RjcSFKywpb43R/Um+ELI+GRlvbnRGAO0oEA
WtzpnzTKAEgH4k+ZIJgot+zaS/shhcQhw07yNWAKzKmJhVc9s7Y0exRjml6fAp9nxmGgKE68iUC1
7jz+CpkO+j1ew8l8H6S3M9KEWXFqnLXcs5SxSfQm/4s7rf43IXQ8JMDjdsX76FWjYm1m1QFEjpvy
nLbAgDnHibwR70HE9OSnEZhEaTD2cxvxiIF/jqv3dWIcbaPqUGf+SNgpiO8xKRxN2cPydhpt1SyN
FvqPxMxVq+iNNUtMeddb5Yo3PL0Igs0HVUDPZO8uMGkvqdNRR5omZqP0Z84fbPTRr+9VQJ29iSWf
bqacSpGiocoEEBft12I/c9/GbR9172XU+QYUDJ17NscHU3l3N021Dis+iolNZpIRhzcp8mWxAlXe
9QWorUDdEdsvObMDm98YD07fcknQi+50xyHAoLbAkcMawtVrh6F2xK4U9z03TmdjFvJFEWG1TQLl
MIDdkFeqKkVg1nEj65djaz2/WA1HAiD1NWVagCC5J5hN/d3biVwadJWNF830eHATrovVH1fckUyN
19qwk36u7QRMhiivArTUBy3zc10fRrl8vJ0jzjqxi9ur1rP1ZAJLfWdoSbsNKIcc4fQQZA9HVtE1
zdH/xJ8OxS9WwvjecvvuhjvNPocvUmS8uAdvocN9cvWeZlcgkSvzSCHkUKE2s0+/CV777uTdjJ+F
mMpiIuGuviJlLHvABA95E6lcFKezgVSpYMbJj8946seSgjI9eWnSo2doT7u8s7MoIIHUZ4PmFSZa
t8tFI9yCxYK0IzoPP/ccdwMXxr83uJlbxoEHRgH3SNuT4sGyvG5uvA/Bwg+oL4j+oAY+xZlkJXWg
kHqtJn6mPE/g21QO3tvl+dsHjEB4EueqhD9QwgpoC46B8yJUcnFk01w5FvJQgo/C8VWv7dDI1EGI
FeMgs7wPKdsaQoABz+hnh/NGXMSY7zN2rxnF+4Unp9O2H9LyLwiWGZtHRouU/fzRhk1PH5IXchwc
oAFmOWX6vakH66BF7XP+1rKejWrhe8gSVbtzWjS4Mc7oJiNuRsHaD8pApy8bGzFjRVy3vL5Qx2Uo
HLHidBKssQAfzHLVkN2iMzbpOfLt2HJy9Vai7SmloXthwT5w8eGcEqvAcMEYtXyy/oJw6W8cT7Y4
vmA8HSPslwcZptp6IZ8xAav334H+V9Q8rFZT/VWoFJFHSk+1Uvi/icGF/+IrRWwaWzj9TcSuCpuk
V103Zbw34AU/qArHVIwgAonXL2f2wZ90LxMyWXhAyJSIlcFhrH413ASOvHb/2KYWmZMjz0BkL+DM
MD5AymK+sMPY4oFXlk8MfClmWytyL0cUb20q3F/Od+71XEwshaWvAdkOoHfzNgGmxWmABEgT++wr
+Q61tOqvj1kTaoqx4HKi15LcET7Q2B8Py2xtyhJxX1FU9RnmNEmW3qD0sGOskq/PN+NAtTLkPiDn
DJsVx4r0ZTLe0wOZhVpDYwRNz0MjC3XtXpfHg1TzfzXTKVQ8CA/R/UXXc5TA/vKayYsuZAVv1FcW
hwTX9RkJdvS3p849+KFJSRFZw6ajjD8ornpwH6ddhwJtlmmOk5KJYb3BwWlYdj+sKysVWxBjd92P
sVoXpSLWmxA6s9tA+hJvFQ9qJ3dK7Zu2/scvDzEUT3gcT/5qlv4SDyk2X8TIKplRq2MEnBO7TCqr
2IN9A0CveOZ73NV0xiXzHsXmO11RYCNkjXvk5HIbODrZPjGp+rkGD88CihQBwx/cYc07pfV4Wj8E
K5YuV2v6rhKbKGw8FQZZrBzPJbrZ6kmEzGPTZEUNhmjGTLgZvXAskAspxH52LhhNgIV9/acu2A6l
B2Q9cJpnaOi8g8T6eZEBnjHmtXttkII3CJjYRYMMCnxcqTuVZ1COlH7qYGxnQxUg8sfsRHTG8OVy
xecMxcUTGX53p3eDmtQZoFY0KLlvdzxRWsfVQ2wMrO2jNKr5CpqOVYvjPD4/r9Tt5GV2CUdF+Ug0
H/3rNlnMiD5RxlbwdUTLCfUQBQuK/PSSh2FlHbxRPdIbgrQVtDGmn2RO2EywgWS9D2shisKE6xJs
RczGu7QkwNpgApRMK2cVvJZo9r7mqvg8TpeFdVtxKegRiK8G/dxRlk//vNjG7SiOx8kay5lNghVd
FHgKG+QckL3bQHAEc/Ed+BCBQLfF94AjjZDWyWk4O7/DSI45fRn6ZlSZgQdHS7AVeswtDdX1sExq
nULzQ4rI3qdiEuxIbe5KPC847BU3wmrwGdbGqEZFmOnRiRs6DKmw5GIL9nfmdHydKrXAhOpLkx8L
sKRza9wXfadqwcBgOIdqzLVgEzjbVxI6BeR3tkKgIkP2+44Ig6LiWyhgRLnCizcfNBOY9DU5htiI
4HeIk+lGXNOTb1PaS8yF4ZKBrpavPhgm/VFFAMcRhbdrjEny0dDDcuGkbp0dtwu3KBb/PgWzf8Nj
T5VXF3EUJQzktsqvGpEmWxHqEDm0niPT98vOju3SE/wHjtq69EiWiexvEnEXuVXpyqAmDpVGFdi2
8RJXek+HiQOa+Yn/QlWPTNuE0iyiZE6Q4u5lxH755uR4+lvBteLNi4xSg8BH335zjoa7hRWHR8Uh
gGT6vglElaUOHMBEtoBS7B8LtY5jTuRKYnHlefT+2lTMg94xRkE/blvNWcvRKsmWSs7YW7QrHYqi
9tOgv1/+X+lPBUW7nhoNvkYgTKyD+J9eS6H/18qekUcsb+3B/vapzMp3HB21VjY6kbD5KGWxYfSt
H/KIPT15JaN+GwFVua6HQ8HcrfeLnxvz6tcmRl7PTXxSf1/7vuAuqf1X/X3oqSRgqBGR9xqf2Hc+
nye2XcgInW2RQRBj4k6DIo/jNWPRRiurBzRHSHxnsgSMihqqJphvymIsN7kOCuRp0eySCMvgHWWq
2BibXmsFxhmWoC49LQN+5RDv7PhmDjdzi1uXxu2V5klcFZwiTeP0qq0Ef5BEMjHvAWdUGEY1bs8T
PjEIOv7eLay1yQWe+VYG+dRIYa66COFTU/UY32j87cfm/zoGjauow5/eskri4gNCPOgN4vX6VQGk
AeIY5FUHh9suQqp/636eRfawQPAy1bJxNzqp5hTt/xPjYZYA5C3sEZH/XYTLMOYjeamjQ7EJIpRE
BfG0yc8ZSKfuZZgLRG1TOC9ExWUHZHaSOYXbpW/MWgcMS4fa3W7xW/YhSydqw4P+81H/CuplZ6QP
N1Rq22/706ciLNpdlP0iSVujsglp7fBvgbxQhPQcPbXtb30oDlO7VHRF1w4XDv/0yypE+wniVCIw
R60JOaddO+ydF3cWwbZCiWbllSLAHHBBvUCldJrNsQsKN8lP86gkEjgFhCImd2/61qBp556FkqzL
GfWQPWg5BptLLr494a3gEyjye1lUCtuvnPNxIfxlguSlTcv1BmyZogITG3vSfKfJ/s7TLTZsD8Tg
141wKaIk+XF/tCwJVkTJKr7AztIGOqCIailS4XQXEg9m17b3jDI/9Oqay2J7KzL5HHhQEK573R9Q
jAWASW6VkgwonwxUCUhivpLQpmHiJXta1aI0KQCp2uT4OgDPT7gpOivRmTLCP0q1Gfd4fxvgMpLN
0HfoyMhutNSp+SOfAr53tPyjS+e/5UpBunB/SG8Pw3YR+g59lIMSF5hsqU8TmFSqTmi9++baT333
Csi6bcfku7EUUNGE/uWnOZohbdMRnW52F6FmqCFql9sngGTUvQAu3HL8Ex2uhKj1UESTY1nLImcQ
RbExixciJFMX1mzNPgE0zHMzC9H6MU2oQQdGu5H0cYsB+DXh6iyGF8oJxLFIKQ7N1BNu9HAh51UI
egLZj92cGOObaqvygQGMy2Rjy4fP8PLyXVJhA1r2AgtgzG3fbuW1mXJMSIFMhfTSd6b6rK5pHSQj
By4XGtAIaLWAdXj028BMTACwwfvVbmkj6GflmDFfxtSh54IT0SzPUHx5he18dcUQZI3SVHkCpA3o
6aH3Dp/EOYDr6anzNUR+9lUUvZnqLM/VfN5zMqiRFzEGZcAJL0Lq2pGARWST7630HZsyZLE+Sbyl
t/x4ZZLpcYvHfee3J4FIMCUxibKfuTpkmSjytov/EXPBopYgdiXRd4yV9+o1mCyLZFtTgufYH7Xe
qz8Tt01sGXQ35LfwfNlDze8RS+ijbqOemrwhZJtI2+Gphuw30MaDjzG+9oPhGTindJ4r1SWt4KCQ
4i5kdkinb1ZQljzaGu1JRLXGa6pCRuHVNPNQqDYB6SIit3msfB3XC7H88FKa4NJTIQf3h9A2Jtnu
VVMcbXCbGt0Svs+ewWqGj97il78tLngb1PPGnz5quCnFgagOgJoSVa1byvbna6bCpdQXIrP1rmSN
LFYLphV4Zj7Wiz/ODhlb8KvHwSwVSxc/y7hmN5rEY4VZ+XZyMhQgjtXPKKlWx0+MhSgrFuEDT2iw
R3z8rWEeFD3pDU4eI/qBM+YWRzKXojKp9WvLs8GwT0Ke2Z3/EzrWRur5DxItZ3XkcKz5WXxekIio
FOeNAAhjwmV8QsMHB8z78T88g5zPY6SjCenxv1l/JzOPPeqDVLZDdt0vu3o3xQfUpi/BhcgDRA1n
e4v3izhG5aaa5pmNwpFsadMiFiGHg6PRzeKCDZQ6dgDsK30wqVCcSxsSKDEGlnBcDw8BcYhc5VBs
rcGoH6qyh6JJ70Xkyyy+zQ4JdJehMqmmfGyAvYE8zQcl9JDMwaUUch5i9+/PMuDOwtZSlwZXuJ+f
k1sxsx4t0mxR44P7zJupeXMPNSIpWeuCEERsW7F2HGUho2yXxzuJgduy/2KkoP2elRJhFfrUH75I
WSTw8jS0jN/WKm487Y0fUsZX+0kiSLk3w+akwtYBZsHaLR7PXL6fazgAIcER8M3dJ+gxNn8XCKBg
3jgqvN4nuXoKzvYTKW7jNhLKjMqE8bzBhb1tfytb4dAwK9Ubm+eJ+U0EW+AQVoy72PLgLQq6uQxj
hsE5YcXiHjOQDkaH1mClb8YAyx7zIwrFvwgYu/GQIIp1y9SMHwdtA61vEc5SWB2ImM/rDkCQBxeh
Nl2d+WeuirTsVBTUi+Bb2FLiLxPg49RnqgYEl+2T/1NXJTI9igZ6Fm201a+9G+L8Hlhs13rJDZ9r
h5rZXSF++zeP2XvNCBeeGifW7IH+aksPomt0v//+vn4RpqiBRaNtMhb+AlyZ+prBWpzj0ghuahju
n5gtK391TcixZEbpCEpzNaOxIVwJzLMdk2oIfQlU5lOqAP9J9eszlmr8htIXhZQxlpYWTaJ3RzU4
J/PC5THny6AFig+Bg1QUttzMTYknvFO/Xuhz7JlKToPOl8IcHD/0w2+c9rbUuc5K7eM5Rwqcre6f
rPboUqcAwPB/9570kcTEJJzj+H2/hKh1sZOApxNXFX/KEWApCd+SmsZMA0Cco87N6rF1KwMfAwXM
yp/w9Iv+C+dkNgVy99yeRG9WvXrXQHXmYQLpPWU/PxN/DnEXAc3yodF6upAlt7PsLgrhJhzU97O5
Pxk/Z1T8mefMYVkQ9vjdjBpVviBbH40TAwazQeW1IlPpHDkB20buROz3MLFC/O7AI95y36JYKATe
VAigWEtwlS0VI9102xECy+1jHPogGRD0UmsK+FCvaJ07MaRU7mFijWr0b0QIyIL9++r74nCIbVxh
xBHDnqAX2LQIZxtuzAcvF5FlQ7+Do23Sl2R2Y7GCEk15XDCal0Nx2LK2aiQU0MukYwH9w3+Vxo4V
kOfopOJCW4dUBmVgRfb5BmynmMXNMCf974XazKGrhj05hBl9ycLIo+Wir8QeWRAg4yXBdL8TSDom
HuYHme4f2rgac4kHK7iWfO2EXPMz2o2tL4sPkQAa5ufzrgTCyioF5VJWWAq6M/5/pythcXr/I3uB
SawwlMi3lNZw35NgX5+crtUTRSyvlznMMRlN4qE68WL5iLj94DrYcnPs+XcI1Wg2kFCXMYcahzrj
8WNm27QRncLPDY0HDH7Kn7AciJ7lkr2TyinorO2wH4Jy9UBStiGXvaW9CtiMXx4IvVn8Ec8gY+vp
6jjsKFSBh7B8HPsSOjJzbvezgVQsRpJxJjPAxX3iP7fww5t6uu/fIHAMjzNU0RwSNpjGfcQnwc/u
UlG6eCdLHgWwoKwwOJj5k+wdJ4IYUKDXmyU/9aKVDUOGGU1rO13AmjXQBhxRV8dErIORgg0/d3ac
2+Kgg1tyzD733xqWpCIBJzy4cx4hJyQB2CD/pdJ0l4+d6RlkJEeklE6MH29fpm2OxYCTRmY8xvYJ
Dv4iQWWsCKJo7RMlABN9UNSAbobB3gGT2o/GCDle5a98CFLT4Aq3DDVvnjPh3Go2qS40RnidUmJQ
AoOq9AvVj4BM1mE5CjK56jbhZly6Os3ZmiVQ1dIxbuhJG2d9X23QwC31KV1ZUXAXpL/eU88TwNlB
/xPPXBqwhSNUmIBnNNCYYLKql/7lCKB7ekLiu6o5BaKnVBQjFecKRUPoojRfS+NvbTy5Urn1PDJx
xRNIu82CNMJO+OIAKTA79VlyLYibXX7e6HarEvHHuCktffoYCx9DMniQe8fwzNpHi8rkEJCiEb/r
lN5cyoXYfOni+0w8MpHml/IsoRgqtkSWA4aXDRFdWQEQ47OdZ04TBtQBUWGWUg18EPfeImUvrC6s
sbDjbyVrW28GMGPTGMhubODEmQiYZ1Rqu2+xQ1osxvOU9p3rvIOs+Y563vD3AJv77PsR4PoW7Co4
vHV6Bhv1EpApyNa7jtW9f3iPOZyDAzrFcyhcWv16NU1MB1Zyhkf/8tLwtY7/jOmo6LLeoHax9Grv
LuTHL9gOZvHPauzLQWSBcrfz8m1K3Xp8b073O3fzbJcpBI9OiBHMjeYiTQ3tb/k1WE1ksQJdeBJh
TtDLcnWrG4af908CBcwnbjSB6wF+sdc+0tsis6WRQWVh4RZxmxhsu8mk7nZXomXb2cbpEzEMaj2u
kLnc5pNhq9gOhRAijPKPds+KalxQd6KbbYTLHiBAez+qZixP1J83CPkL5Ig5XHA5tuWXiN4wPqTq
1GlAg83+IbSoc67gqLsRzErTfAu7lwAWLQ5Uxp1fDCr/i8ctFH7qK+mzzU+Yh+K/Bjo2k5UF2dwy
d6LLZ5J0yjYd+rNvtTxgQTMr7/iIXGxXGk+ZTI7V9T54ZZTQvhYJ3uJmYPtGgvDLyCglDPdMXIes
xuG7IcynoWPS/GQoc792BkEtWEa2oBGsoxJK5cNPi2yK02XZfqz7DfSHU0n9kn6YF8DN9ltsu+Vg
OkuqdxYL+2Nt8LTdt4ux/RMfoaXK4/4Kt63AYy5hKIanVhzMRDXNLSzcRjuwFKvL8KDL/6Qfp3QU
M5hlA302AzzXo52vd+B7rBIcLJcichjnuY9nz/KHggaDcOvWJU+3Gv8M0ZvPcrmdxH+hmQtiu9T1
B9K/LFKbVcsz5L0xRtl6tbvlohwMqrWbJuGcBE7P6RirGy03J1Y8qlsQ0YQhHVV3ZKyOH4i+XVM7
ffmDY3+2TukOhvD5ciNbwGEybowllsotIF/MW2QgNSBV337xd8dibPs7TlPXAd2za3M0Qhy1/NUq
YZWBlZ/h7mqezzd6OC8UKDqflZ2JZIyXv7sasbzGlo7vMR7zSPx0BYwa3sOjwdE6xy5pO2mrH0sO
mPFZ0+TKEXe1WMEfrTDzV1bmhTdzh1MHEkrTEoLtEaiiv8vlnnEPKc892fcfCnnqJboj0JlhygKX
VvgwxMJJrA5j7DdcwpIvoCPC8aItSDaocp2YskRPOeHZlxB84z4GnQB8K4x/jYqOiArlc+U0jJ2O
GiidnFACjPzDc5LIja4R7Xyz1xSdW8+IktTwAZ/js+xXVncfAUO3CmsDK4gpf4QQM4snQKAfyktz
/0/++zK78A2t6gdkAjFzf3Mms8mD7vVC39+9xjKoDa7veGZSSUhD9uar44rjlCrMH0YIekM7XOea
LzzgAypwPWsOfdGcKhDDcg8gAEsbahM2jBv37IkiORzi8O2fb+sj7K+ort1eQnrmkwmKvDgyRGEA
J1XcI/8d99sKyc6qXPkKXqcKyhxs9UhVvpAesIT1EQoJ3YsjYbO4r57E9plADEsmEV5yGL0YNv0n
Y2InRpwwyNgh6zFOn4HGINOVQ5pIQxpURt6CTn3p6zd8hENeEN5IOPpL50jDWhh+XQGKlKZDObsS
RYvdmboQ3cMmVCHlMlrupUw+DyXEwCj9Q9loo4GOVdqEDHz2iAuEhjaKb6d51bl8qvOQxMeAkPHo
1b3Eh3cLWe2zVAEeRK8odMlyb20jj3/Ck+Rqmx56JGn99r0OUaqqENS9R5mmDmOo0vnYG3SXYXx7
ptzg/xcrxeWkLmKZf0qYm3/NzXPEYT92fba/a+H+kcKLF/TbWt99cW9tbXNfgjaVF4UkWZuvPokX
JUS/dovfdTHMqxzoe7/fv5gsjZeoH7PEzj5yndvcFsOWORmkc7KVo/WY68feqiklgcJZegJ2PQ/W
uPvFaP2Fs36BNUPzg158WJHFrx46WZqbnP1fwxLfL2sa+Ff+w7AoENX7Llponb6PG/TPWCiUBW7z
FcOheRv2FwQPot1Wx6Kd95BA2aCwIJEpXTvY01q3z7JejzHLr7tIFvv9fVUxzDXTzDeQ4EqzLTOZ
sqDeEP2ESTTP9yE5UzcD8a4cVyixfO5acrPyqRzLoy3fPjx1NyyigtapiPWCI/ys4gkfMs47CjuE
dFR37mIP4HV46DOhn8+vVNcXIwiUjoshqAddCvXcEQkdRwSwH1n35kmXuD0tl+Yy3NB84s+r6Ju2
/y6evbNaJ+JX9hY/xVMrwtBwUECsYvpMh9hiWys4zq8NCxEiGg9ZKpTEZ0rdFRkHgK2aH9g/K5M/
YivhJFrjD3/JW4o+TWDrEwCJwsZ2FJ2OKZCpHACY2/xIauVPN9wFpQqOCXTW/WdR97/a3Lj3d1nN
ErSePqR91r4mkBOqo8g0p9Rbb2ucpMT0P7FuqKtAxYULtY94OwXLqXZIdZ6FQAY4dQ29D5ZfywGH
vwOoAm3yMnMvdWOaYI8YMwHNF30IKeeQVQrZDszH/G5K6gCg3YIu9py7Lq9oHoYI6T/S5//apH+J
/20H8S2Oxve4nbVbAUYyVfGobijUZsQEU05LFN7sNzcw01TWzwYhS0+mK+mBv+v1QTYKHBXCm/lV
99+BPe3oaYLZdbhfgAPM6VlX3+EvnIJd0G1YnYHnbT72K7YJe7sURwwgJJH7avD46I2RXc/LU8T8
FE5H5SETnJT0c5HXqMCb4r4AsDi78N93bJb9Cyu4qG97EYKUEHr81xyDAjwDGPDNcxbpVpBRBy6A
+9FVFZxwS5DYDtMLQEnOyphlOjoZrX/x8Q3l18HLNBlHLdBMJOtq18biJ1iz1bT6bzvsd+5w/miN
XP1JUZvjREys6JwH3IEvsv9mXoRx8iej49MHAJPHV23O/cnWRdKFWieftsRhQZKojeUuventSv4d
azfb4b3oLJpd0xQ5RH0t9jnvwLoACqxoj0opwGQCnnw8eRbXhOBuKF7JlfbYXXbgiJPpCY8O9LP6
ycGKQ1Vda36VX+95iY2Vb6MhZbRzmKlN+soDLFoNqi+C3syQzw6YTH2ZmUip6SInw4T9d186tSte
YTFFcIjYyLWbo1VYckjMitZDexcOo9Olsv9cux4axHn5Mrp37KrnXlW65gMXtt3gS7QpmmVjjq3w
wNlQq8OylI3sj6TtvgFC0gSMsg1QaTjPoDQ+Qw1mw6CKVix33abggAy2dRNlkOcnknHUd0XAoIag
MgpPPQyJ38P/Nqg1Xl20L3SYACNBjsas3+x4w4ewEtRII9T/Nf89PwdTD5OAwHYDGJeAiYZJhCE6
6P0ysujrm/EN4ffT+S8FjElIdw1x3ZDOgChTEMX6wBdtKlta3MTLfJijKRYzB1FArUGBeeA2v4C8
J11tHoDhtk0U/dFw37li86fgSI9Nifda8r+mJkWpQVZntblpP+DlfcO2k8Evn9J0f84WwXSBSkS1
tSwLjd9LtR/I/Mns5UgW22tzg5OEXTCgmYVjn7uhFd2g+XJngrgHDfPH8p0pAmjsAsemcUfxwh5e
IWooODFzKHlvuXbZjacvZa/p2xxX34qf9TJ+V/GlfWkpRLMNHWf1s7AjEmBv1vUyBRFZA7jeFrU7
Hq7JxLknhLpC8j6jeBt/xRtoeswCsYyoXuQkM40TMCGNm7qAnr0uPucu2mHtmiYBAanl7xboukml
MirlghIZIsgsGdrPe8S2toZYFvVdj0b17a2+Wa8kJS52ilEjDbcf1Ej7J3sQyK1mRyRP9V8FPHY7
chJejeqCOKGCSz36xNSt0XoB1ti0tcPKtDfELUTDfrHSWKZxLObG46LcAv3nzQNXDw+hHQgRFSA/
NIU1Pka4fRNUheOT00QFK9lhlNqoKipg8oDuE7MjqOCRUil08JnrG+UvGrxMRsDT/CLNj2xMR+vU
EyHVhNXTCQoEogEAFEcoS95aiet7nMpPVSk9xIsx9tBF5m9ZK2YhFoCJJ5Zpb0AO7S1j+2R8dpWn
eKoOZZHWwEyUa+9Ni6kA6X5AFBLnC7ejtK32xFPj3J5lZ/lAgnjJO2CgCM3HHL4y2xhTU5TTjJGA
svR8gXH0QuO6tnRIOhsFoDWU31sdxspedq72tjq9Fx3OFDb+855Ba9nImZumwLuu2LFDcHiiQdNL
biHwqbMuMZfjRCjXBAt7j8416SVNPhdRYwq6LzpECoKoVl3dZfnOrBjOzRDkFUcmuISSBM/EzWgE
+oTZGISObsaPChiidnrc0xmzYI1HD3Wqhx8CuzNdEh7jh9Z6GKH2iGQDRU+y+oMicds1ssQC3jrE
OogSNnbPnGRB3nWsySY/b2tu4XKOehTMC4w7Tx+FSR/4Mqxzw4TI/WI50yjDbi8vIB+EZpkv0qw5
KxYTLGvrplofJrt1x2LF8KiyWwAVGdcjQ4ZPgNBUL2dV0v4EID/qlOkuwrhLiIsQuFfsILXNQ+0G
Er2DjI66fAJVTTNMmgEByiZ6uUUUr6J88/wcIZ/AYfq+Kucxj2Q2nTxNAxDvQ9C7lKbDSJNbz74s
Qx7qTzljWmZ9QDWshHUnoeC2+hkkvTeKaMdisMCBQ0KgIoLGQZhfXGtnV/NDrrgLGOECffWafPQu
nlalKdhll79gWNCneJp+yAJwfQjxZmrIoUT3tlInMH8x4NlIu/F8jGNPZxO0LSuP54H4UIz1HOBS
yFW6BwFM5rsWwAFJSbCtBrFUfBt9Jt/YK8Jpan2ZJ/BOe2x7qFGze6tl3KPd9GwGyldAG/U6GsIW
2bKEsbzhhTRaerOXO7PEx/J+OIbrQkp2nVjJXt5QxSpQwWukaklZLFdX550OGgBS8n756RIlHV4C
43U7R4AKQ8qMhZghTeNyYec5BQsYFcLmeC67ceMPBDcTVzaGsBcmGYgrzGfxhZBCW0vgWLwF2w5L
0T51xBtxkD0GSVbAJ6fuRslG8aQsw1jEmJtq8ilg8Gn8iq01KyV3Pfya1EnAH/F84+BNUSez6Ldg
fYeZgv1ci+ljU/DAcupASBoDXf9v23VdMf548oPexkjtEfq1Gw7EEginQECdVIGPinaw96QAQO5W
SOK79ennpzIq3+ylIggS5g1KKK5VmtEEQPtJYj5STM9zSnXscUJFXfNZoKrX7q8G5JgrDCN3x+U6
YCmkU9O6CL9W7JRTi8em9nLaWAvh18rGnp6FME0hh5o8pOGqt96hQ4w7ZcopePOKCG1vcXXXlw91
ibYzRuTbyl0dn6+nTO/59vow2aFqfNGwAaO35nfLhFJwJD6LemWnc9L8WYCVRqH1cUBQBJ88K1Jl
yVNY/rp20vNufXRYAZjXDaDw3QyWp0vDwD/C/7ZA8HwupcPOM/OXRBKZpgibiiLiIcbbAUUj7WmW
FE0GV3ZqZeV0YwVsj8BM8lM4ndOemIh/BIhanPdeYQy4oeBemUcnngh/oH1hDw3ctD16MgiUyyzZ
eqandQLYw4f8Z9AYFfo31UWIFoWy66qlM3p5MX0eukGwKXj+Rg9hjv8gFrOexsWX8uf/knYBcpDT
36LkoG30v8Lc+iIKsbcYnhvBHCW3KQk5tJsme3yIj4WeBr4YJ4Gc4DxqJ6nawLKBMXqA+RekMXqO
tPywdi5nl3AzympSYm1aHGV376y/NkXAgs2mlLrTloUmcXrFMLXfDpms9NAbTQncw5/FFxdBwN+w
2qO8ai34kJaMtPMzi40hwjpz3bvl6m/CB+hbN8icYZjYRWyB19WpDaGAfngIk+TTYgDTWJdMSC/L
nn0wffmGIo+85wfBH8QNodotdyQuD+bfW7K8lcm6PNycU6QsptQTyKPAuh1GWJXgXJKZCRyWG7/2
+69IgiZLtUkhjAO8sS7vo+dsdtX9MjGkXBSv+3mhqjTTIo8VwD3v4mW5PTmJwuiIEwX1t3CNBShq
yD2odTxXFiBb+HDex2HyaV+7AxHk4Lu/YVAZF+Wf7ueJANtW2UdICWDIyrpSzDszjWhBq94yqVwf
Ghb8Ir4AQgnOQsbLtl6pPfwceQYO3Ie4T/qlFZ/BePuis/K4Eb5FV7Z+IRATQVhnSaqvZ9gPYH8W
xg682/i+N26wdYij971HY+PGLJgNMCwIar887oqmRBDnlZ0+V6HbTn8tcFqJCxN/O8YaDEuXLZOy
lg2AYfLY/N0rrXEXLZZZrpVJmSLDVa4hzBT9c9mZeGEFZlSR5xB+1gUMnbewHRWmLE7efuRmM2RH
dsnt63FN+OlZTu49J3GKhAelDLyhHmJ5wkpJNS3aDgMrU/cNL/+bHe7CGR4ZL2Yo+sVFe/A/F3Fc
OoWyIafe8coOUJMpTtDpwXEB6M0E2oEZFTsD3egFko2NxJCet4Z6+LSLTGPq13ch8/ZJ3hFQSu9H
iU8E4SbzhUE9u54iZCpuOj7TOf03oRNwpofuUfWevve6cdsqt2ryAFt9oTLl91BgfxmjSekA7//p
bB5pMtOO20fkJFwy8HGhei+wbBlbQmyWOjUClYrVv/GMt2s7a3LpyU8k4nuHN7qxxYSQIEKXs+cP
PjOnNxZzU9/QPn29TZgy/mYxF4GiFzvTufGk0+IqKhlIMZh0V8CWUoDvyQtd8+v4UtRlmXU0QgST
wrumtokttMTNwOLgQ3cP7/ZjWYwZxoi9al+tt2CTkrd1LYU3SK3FUVwCS6khoLqGs8p2NuowxmcZ
Wnlrg8TkfQo6LS1ssKG48+n/zGrQowh27EXxugLlkbGSpJFke+b5XQDYGJw+9htzIOUKjANQp3sb
S8EXJe4nOPwhKfhaknbWeMmcMoxHiqdKY31FVoQfwFy8H9hj6c+qw9UusEHbDq4kya82E95VT/pc
cM6ReYRSNVykdN+gZ2iRE5m/qTXHU3lESWUFWVIc6iDE4ANMLdQhdU/Kp/hHjgrCu0N/xQV2dWj3
4agOj+q+8iG/Pvqzb7IhhMljeHM9/i0SKrClefumkgoEjN/5V5qA0bYzm2lTl0mSoVabcqRFhISZ
bl2qiLZ3+gcyY1IE0DyRJ0jJ12irrH6c5TWJjlwCRbMN6vyd+b6aVNOIzYDvexBhF/MU78G/xRxA
mzEF+k7Zdk/f5Vm2C2hyB07lGhRKeUm+1wh7NdWRqepEtxpcJ4R5gV5HMpaElZrnGof2WAVqMkee
zx6zUX6pUGv6/bxdoK+8N6vT2gyWZkVvQDtvttjlHCWA+TyhrRue6i4S3YbGI0j04yYzN/JAFBvr
7+z+QYbJ5mAAkryx5F7xpIgBFVymb8mKaG98gQYo5zCNG8wzAbJhSfoFhmgIeiodVYxADznTJRwg
76M1ZU7zJVEzq4+WbsvBmBE4BEK9m0u0EiLS3rsr3hWJZf0mW6Dn7hdOiwjglEdAOiQkW0ytOYoC
o90/ESJ8Yla/KdxrJwupDg576J6Yp4q/gQQgbPXOzxOUL8QamA64qdDN5UV9na2kBQZ0ztesK31r
LSvfoe7u8PeJihNP9WBdJml/wywSiSkP+jQ08/GH5XViu6wI+0lGoLaPzVS9bUzAkQecIqRyf2pe
RSIPDY6N2I+XmhzdtxfS6wGgUZPR+uy5Rm4OooyztYLE29IaCflJ8sbX+Mvz4Lv2TaBmvxrsrprE
IVdkcx4a9MxO1UHnFbmWHe4iA+ozZbvLxeBdSnYDdvaEeUUoE35CRb4ar49ebJjJHpvXl579YafM
+DU6yXSErSJtfZbYNYwGdqBXGa1mVRp2QZSHNsWF02WsjM7sy3nIIUmnyU2MZhtEAx7M3RLX8F5K
Ba6KzAOnkJtWYki2a9qGD0GQQCryRRTIgzuKlNIQ80g4PCcnlwa6Ihd2vJ9JjlC1iSaKcZKJluJW
g3ZXbykaY9w9GMJ7Jk1FZ97EPTgzneRKvAzlghR4qSotzLa35r+QM0eGpDYJSqyNaGHn+F/AgZVv
u7xEZcAaPhJgQZeXG8PRfzq70FGyMCYlJouFmCV/fO/i7Na8Si8YajtB7tJnaEnhriK5FWRipWyI
BW37+DfQk0B2YiJ+S9DHu3bEYP0tuG8URH+HVmmir+O9Bwa5Nr7r2ddoWGSOVtHypBf5Osfhf2sP
uC4IIj1Lru+efzTz0eFgsvl+ZjHmnxpkr7dOj8UMq5t5uZDDjD4ZM2WbrXI1jJbVsqz7K4RcgzLB
wmrSjelDoHRQKRvcvTpvIfHuJjoXpj7bCABJdkB0Wm33nFP/E87ifcAVUIaCCiHY2WNtvjVdwCbY
87maW3/BViIXKO/JjcA2fahoTM4MNi+MQ4HKPXx9e1JkA6wQ/kaD0oWNjGbrRG0QmgDZuVOnOkaQ
1vRsp++fzFwQnqP+LMu43uwomoBOEK5KteAxgow7PLd6gLJix388gEpHMueF5bdKJp21ewBWz0Z6
ra6I9ZwAeGhZ5OijlpIkLFKtvh5531HFuIs1rL1jnbgt/CkXB0BWoAqJUl+55DReXK4NY13DndN0
0aOlTXrtDigGMmzfdEwFdFcxMy5atZ213wcSCOXg1HSQ5Sfs2t8jRtA2/E/j6X5ZxEpl/coY7WA3
yNQKJf0BZ68T/o35HxH/NFcvsI8ytERHyhkdXNKTh37pLSa8XhzPGylAmOQuGOTrdre+UVl8Yt2K
V2KPPLKC3XZ77tzsRnVFiBvc0iS+grfkj5wmcQhVc1BFDEIV7aRnmujAGiqP6EhIZgDtbpo3cbLD
K5WfaZFGaIIv7hMHwilccDSGF31UHROoVCzNEg90zcpoxq5zBgdPgewxZXB9adPqQHusvVudL5VM
QlWh2GVzIA478NKMJbi6Hfan4QULTiS1CTKVJBN/XTCsbNPtHAYVuVMZtlvWzlBd+Q6zlyolAU+H
T5olkC1czUcjhAZtAtE55rR2l72s5PjXpQGar6CBOLBJjOIeKrTBc45wxm64OVXZpzVKTv8J8+Nq
oC3XA8PXH8Hwh78ePjf0JgAxG8Ei8DbgZnOR6+7dmw9/AchRnbrJCtrpG+ZT4Jz64PziEJCRJEcK
NuRMa2DK3RQ5Fx8hXy4ZH/wQxO3JZTGCpnYFGrtTl+bSY7IfRjBXsammB0m/et0EoA05N/Nlc8Aa
3qon5yUMs7tYf6oMjm52hRbJA5I/nmQGOwibXVgVO5WIfUqX7nkcDzcej1kOLlFzdtDR8/NFyrmL
QWucQqfVZfrKIqVqwcbYsq3WR+J6zKFV4ceTRVQyTRHry8qbt9S1NspFiRlu/d9X1jcL/oQZUPIZ
MYIwAbTaA/CgymNZ1/K2jMHXK7A8KT1OhMUFrxAdz+U/DvPJeO4FjjPuXFnyItsr/XtU6LS2Nm7B
44wNWari2Whc87ta8t+3h5GZcFmpzkZ90SN27vsW0LN3ugNVBct8MmOXSzLLi0a5HjAvi7KQw4Un
AkTCafUSpwuJsaHOgV18OrYcKUsYn0qhUGhobJ+QDyfmOYk7wToGOxVF0OHvIiUgv7eUE6mX71YO
uYcupko8xFkj+msxa7RoyUrFxO7j/74F3zbr4W9SAcyozN38CiVloCVdYhowC1KjJ8fMP59aEdox
FUbo1IEBwuCYle2DBSBcITYWXDaCikMeYFb0Zd3WGLUh4fZIcaaHNrwT8KXJB1TtBkrRaT3kA8sm
Wdw551T/Ob9QXca9375u7Ok6s3EYNVatDVScIShU1Fi11gVAKAVNS76r92aHlEo8Ftuip5BzB9cy
sT/+P9mRPWhB10NILZ6mzNjPdlW0Fu1ByEzsVXZ2Jy2EQ9p6I09Q2KxzvOwyQ7b9YI57LLNcTUB2
/FBXRLNCb096AvhwVLW9meJAG97QWq1Hz1ZxCnBpwPxn+C8OhgMZUeMOoJn2ysZgWaokQ10yAnX1
YQ9UrgmF1YHomUT7LRuP32FMWOq87aW4B0oTuYuGAe7gFzBnlPe1I/u8ELtjakZ4SJzZ4OWlO/b6
LJMdIsZm25uWYh/wLWGgfGmz1Ssv/IXgv+jrIFNMPCg0JKcudkh7Vn83DE3rdyn29LHbZt97HCMO
sCCjtiCTGc8aysHj1nB1JjUde4V/cGcBGfC3qWQ21cULTu5bsM3sRplsdWsUs6TpYDXN+9wtRbJ9
3HvV1N2G6DYSO2YLvlH4WNl8gA9UNitWbFSCw84d9F83XmHgpQur3mPbeQcmVraoAxTcZqy4DTds
NleaQvM38+P8bFvRLU/GN2zbkUbYxeMtVkOpYtkfJd8pbtgJDxrq0MvudNzxck86duJJAdHqetC0
3O2j+Iaj2vgEjRak4lcmFdzoe8xHMUpqIKQ8jsBWmI8dCdvePVUtNvopLn/xCkGv2VfKm+wx+8qd
UMe0hL1D0ek9X7cI4HbG6PAvEnYfcB3Nuz+Mn4MwJyPOZ51sUdeJbPRAoSztihHHbs6cf3y9EWfQ
HjYStysHJFFqIBLoAjMqfEQKwjRvI7Ca1taw2ZYnpQ4A1zD19hbDP11JiOiJ9K6qg7eeY1QFe+C3
xD5UKqpFotDCCZ/ysN+7v8fYCkuNmFAgP6jYMdmqRJoRQeggayYPkd+aX3VzKDwQtUsazqHKZ1AN
yLABBacyJvv0uuc0l0/L/qUs3bivMrJy/QnYzZhFF5tHH8puf2PDHEli8w10LxGikUjMkQTZW9Oa
9JGxvemO6yB1VwtdJtDc326s1c7uXKVipOGzeOnUt3qF0I9yhdhR11AaLqwjtez67Fn8o11MOOED
eVZ73n+jraxDkgALdEb1Cg0I5fftegTnnplhYMoOUtAY2poJIZn4Y7BzGrwqcS+ORQs13uIwCbgn
E6luwJjtRs3OYLK5eLY6plmxNdH4RTVUNpGW6jyiorDOSwUvAxC8ObnBZWXpL3yvjM+nTvnP+yWl
AWQTl+Zwx5/1Uch6mAm26iUVI9u3Ma1DSLWNxvinlYw6YNA4N4SBsMH/YoGvM2HynN0ndMsQjEu7
mgoQ5JRp6rtu3fq3oCB7+KYi09J/+xjt2StHTG+J6lx2WTfmA+3H+XfcoVgHeO6hHr3vtqMpWyrt
Stb3a+UTlcFmPmwASg47fbuio3Ha3D65YTJrhDCzRHtSyCWEfmYySa2Ww4WFLfs4Kr3uJUyweqwi
BoZkSo/a/xAxQU/fTnmeIGPVzty3ntiVj1Zm30OeJpwUwbl3FI0vO5Hl6Eimmy4DHzoeQF3C14Fv
+pkWRQpwsrbH4YmNx1HaGQZdM7eGFzgqvzrp7eH5mKypPP64kRNWKXNspmnjDstKFiE8j41rv7QW
9K9hYKudrDzZmsfxEoVZDl4FOp0CSyL2kfIWf/MUNgoG59NeWsz/tJfP2pnWcvn1m/m0k4hxA9gv
qg91QKJ/D2XMY7PRS+qGvlpcmJPNWtzc10FMGKoSHOdWTqUyWygLJtY9jGDlJmXa6y5LtHs2R3ox
t1wR3kkw4FZvwXh+U+Ww/5BwX7yl4lxGaDrBgYqKymTuHvVSZD42L7sLmQPDj9q7bIL1uYqV0FFN
Roro7cIhcKHqhJcm/gGp9D1UZlncUVv3n6hkAfbkV+8vLD1VHyXxNIw2BQP4+gvvdPvRMk+c6zcW
vY/Qw0Kyd/oXmMwswYcIO3c+e769yDdswIXFV5afDRLOod45qxFq/lF6t57R5UlTq4enfnWvKkQt
drySXCTUTpDhqiJEaL6h89bV3H4Cxm1HYmstyINwmjOfuyIMP0AmScsabhaX9bt41AtCAZF70Bcz
SIE/VkLP/ZPHdO43FXeuXwi9NsvviQkMDNYwXmDWapDs+4uy0CSKm1aPgvbUpH1Nt07B33l8KBTB
K18mE1Ymq0SmeAau22VMM2MPLCshCO7xqdzBvQK184KJ0RLJuhTkDhWAjYQHZvB72tfeazMxVITc
c2kzP24zXVBSK32pRpkDY0zGEtVX0/S6z+CocXM77z5tcFB8woPKGECVCl9sMm4ZSnB1UVBti0F/
WfugNdBhUHabQiZdGSp2D1fWEzCmtkQiYMPc0YtwBkrxL5JR0eaTjx/e94JN9pMKdt4u9VQ0I9+W
ao4ALfMorYJmQnrzjjQHVkfdNpCIv/HxxqbF9wu/aC8eL+gJp2lbcgIJ+eA821+UUIkloLEk6nPA
94ON99EW02EakchLQx+FOjv78ftmaBViU7HDnC8POWa+TV42vop9wITe/5u5S5z04mMZoqtY4ybk
5MvVmR8N6c2vxvYbU4TEAtdsbU93GJtDsl6yEesPu+b0Pvjtja+d0rIfo7jtFcBpblLeEg155tP9
NMpLW10ZC8blKbGgUyLnZpm4gPhohdBpR7hWYxVIjn7+9ZCULQiuXbF8f1U6ih47joplJzgGu4Rb
80nBZqrLMCxIY+CgOZONT4Wt9jRM7B13ARioqVnZSt9gkVH8e6V4cGkLYUALeMjYeSBBvuI1pYS4
Rq1GFaMCwDxZSnFMbnrtKnGMMaYOyCg3T+F3rugev41RGjnBycSBy2MgWCXs2Spryx7PJnrhVtii
1joE0TQP49PBAv9Us7ImVeynahy696040v2/wUqSXniDPoEji9nE8UPL5DiaxjL87Hhu8Ozc8toN
zks2ouIPy0KIPqhZxQTkn68an271lSwJ6wxhKS7Slk4wAIeISqoEgHVANcwHl5M5UpgZ93BZbLEM
eQtpmIXTNI6i9gSftJXNgUSaRq28G2Mv6hFrIC49fQ+BHnX0+ywB8C10xUbVLn5JisBVgjfdyUSe
8Bvr+2BGNT5He9FInQa8H+5iQyEkHGf/j7CK2nepuNvAenvgc77x8OvN1iDCuqYWVFSamGqCX1Fp
toiyOsIaMQOZpVJLZMb1DU1t9jbQhIV/uAAIpDmf+UBLwRURn+znCzQ4mpJW+Gd1iLLVi0oHzQyn
/psU0hEXXWmx+r1JyWK19yJwOfubA2Yd/Pr0nLE9kFzKUO/4ebhok77FqsMypSBAcDvyBQZra3ra
xHkuUZu4wl/VUXvlVR5RmCT1lWZXXXqNPuAOocIgbmt21wAlA3FZucScDJ9fJwCHNsVWlnVCeGmU
RtfVwCN/UF5esiB+qIKui6ZKIm1y3kADfwvRqGFU8qiRksp2CGJBlnTyoSLtmKdxW3a1No55oEs1
YzlbqISD2y19IA0NZzGXEE8OgACJN5TrlnDMJbKgXTHYgXKmonrht7KogqllCTHDlw9u+661Fuem
C1fVxFTlixoP1wAmb8mi1JxqdM87Z9b29jUjWUwowvWwGUgzjIMXcZ19coI31Hn+lON+hxpQlnWC
cgFnUaTjkYn3BJyVDDdORHyvddrQbQ0r9nQ5YWzjy5p95uMeYgeT8kOkme2y9LYLBYs+SEkk9G/R
AbpaZWDsNnGSaxXoviMHT/MRlzxH95KsbrYJEvcuTjLluTEQhhRv+KhdU1M049zxeOxW1LPVNfhh
q6yS8FrU8p8Vmbb0ztxYGD3RUdYo7pHlALQCP2/E8S1lWNjm+cKmHezbSIo4s3WgoO8dMqYBSaQj
Rwx/zRzJw73I6+ul39H2OKxRUedMl/+479DNkCKfdP5Tmve699xl5q6ekshq2DgVuQgxAOeLUCEd
wLDiWfVMvIFAUdtUj5wxIRkiG0JumL4ESWaY0+D/imT3H1ZN8eBJXXY7z36QYIVEjodLH7K/Q4j2
5aQisj6Y6d4u3uJM9gwn4J6gKHBdcVFdEs9sFq4IdP9aXqnF/Jl455Q/vQpE95Mahip4K7BSYdxb
yxixurEkjPcHgdORpykM8LOBQJUeFLGHtFbiOtPdq0rynqCt9sgVGRlD+2TYGQ0/837dEthXo3Pz
m3t6/cOQ4EgLbO0k9sOYBoU1D7fEhVkkyJq4O+DUDvqgEnAcrQmYBH9B7B+WhJ003nqdKFFfPA13
yBScjdDBL1zqF5JV5oCfOW49QEhge6YrqcMcw//tZBP89aGo/R90hP/TMO6G6owAWEAGJdeop8+v
Zw/jvBw0gdNK72OQVI2STD7JkewMIegzYrFAtpe2RnRn9J9uO86/B0PD0Mcxt0T6W3kORF0LRz4w
MAFMxYtWlrQBZTEzDfyMdMuTYFgtVAOTkcPJR2sltEq3YZibq2RaE+68hUQAk7d5eNnVexNyh9HL
zOFuEFYlrujf5MWNw8PINmNaphK3SNpsKzvtipNimNcJJ7Q2S69wTWbFJVyahN+/pBW8fVH/jj7T
wUUWpB7BOsLqAnsoDHvw8hEoCEe0z1hDARu7VfeQw4oI8N+TJ9vI6PwuId68ZoRIFeAK7eGI8uER
UiwFvvvK/svHArkKw042daVgT8l1whIKUwlgT08xebfU9Fna1Dheo/hCr9qWLeZd/jjVte+1qeSy
43zPfafumImDu/2fOMl8no2hSZ2ZvAmbh0J/fDjB2pPEsAd6lqXQ89FY2wbcEpQa/PmjrsQS3ScO
cZ1qCsyJ0zv2r39LpRY+T4FkktweDUk28jJzct5XwV0AvnByFLqfH9tBIH39ixiqw1MrR23mOPtH
/1jCztpsj3cow36NTTDIdF3Dp3UCihAwWzHUL4c+bnpOHHFr+SfGCX1ZSw1vT4uJ0JkFWqd/bqbo
V3deQi5d6o9KeLvmrEH06kCF/3lKYz6q7Kig86avLDdRkuLu3eQcFBw2aa5rAUT/XASoeyet01Dj
WqRaNalqA8t6l/6NL1B85D0NKrZMyiwCh0i5mXrEWqB0rILutmYW99GlpEjnArti7CQZkK+pvdZa
jDJjQWFNBWFAp1rxt/lNkwFtsLq6+kmS4oo2Eqt6bgKRGl18dPQUxpDTC83A8M2VU1d//2jbphPY
LMtwITIO+rQaprAPfm3vVFdLcOmiqJfmQUjHVcMLvcMI452ZskuoYyFOJoNjhGTp69eq6dHnmsx5
qyIXoxWJt6/Li2JpCgKjD2hYKinLvx8uOIzHz6mkxt0iCnE3j1wUbMWrm69v41mffUAD821xdW2c
b2zj4Tx3D5RKLZtkm7NTqXjCLhoZu17yr3jtk4KU8eALRVF9xxWjNlXLBI6R3dxALx8MsltMbTbI
AC8HnZegoYVocSPW4TnXEMidqCz++PwUQXOjanpfAzTExT/bqLoTSKjroC2i6gcn4I4hvuH5Etv3
UImsHtDY92JsSCdz4Tb7tvWWnBnd3rKN25V/n6QDI+5seKZuvF8snG4scptflWOD0zqNx/Mb5wC6
rrmGwAm8/qYxNBFHjXOWf2E0b/pgODaKnlThtUDfswu99sSz46xDAPBzVbVLejLVGOPDbehyx20n
D9qCLjmy7UAeWNldTCaWEuwwMNW5eh8TE6vqpG7a8ZOXWUBkm2+NGtRHxH7Os/lkL3yZG7BRzqhr
T/C+27RY30As2nJoIj3CW7e5OEsiqmXGpWbER0fg/+RyujzdhfQtQTdaYTnPkOvwDFUCxvctyVmd
c/vuyObq/+pBmAIa3c4vIqt0o37ZlWGB1iNRkzFVPqJt4KZn/WoKoFRJKwmR8WPao/mVDCLDUJ/l
scunYl4vwrOIlIWVkuY0XoLHPPYJIp7xSE5mW4Q/JKiSX5QPXA29hape2ps7Ia3q04QShaKzRvXW
qI4m8MzEuZF36uEP80p1UA3uAoMGw4uzgemppGJHL38PgZgrjYwUjWEBhnT/shJNGOqnz15JtffJ
NytmIZnXbmhp157CdIi3QWU8Uoa0kooaEIe+8CtQUt0iufBDrHZEMzk4VRioasqgXX5t4buElsqM
DIBIpReQro3mPrDszk7tSKGPpqRWCwD8Ku+wiBj4Fj/2VfaDkLWiGb1ulfT3OtSBR4BYjdMjMN3m
cDH9gpaBostNK2kRk+gcJB6zSxctLaYxWilzV+pTDaquCR4lnSx4BwAgedS3fsRO8L46vF48YoMu
B4NEVU5RAZnmWJNAlPycVwisc0ANc14HjPzA/LDWly4N9qc45MkQfHKgCTotDbuYazJsKMB5hL7p
lQophhNYdMvr4HHKeECU5vz85k6D79Qww9OZQiSYcq6/BNsvE/Cwn++6ihF1Izb2qTUU1yTn1FV8
4Khr7nZLpW9VJTz3+sEr4Qyc4L7NyasGOXyg/wdAS+qZHBMUchPjmvD9uSEOQo/gr2w6nUMEy8Xm
HHRffhjKtFjY8VzySVDcu/Z2cmKkHKnQCCqQOVHK55HfGdI9gy75BUClEDyOmZDC7Fpy6BA5H5N9
0YX461Z2nDqF6V7Lj4LPVDXylx8Jn6CkDJf9opVRk5SMxMlUgslIrKO92hg+e0HOiGAAPTV5weDt
bEUS1/xLHhwl7ejShrP1RIaiSF8r5Ci1wXNUoAPUzXDxvpm/HZE578u3p2k5eaJptmLYN3tWCPLZ
x3+MQR8YYoyyOk/QoCKuaBCjvMXr4SvoF1jjCp9Bn0fEUPrzogNRah300d93sbhx7+1lNv/XJ7LA
zqJZ1Ro+D0NkGqbyGbySP8lEf6PbmlruDORGc/bdrbIMbS/3lypA+t4+JssomLKfNl+eq5YqVPB5
jazTyOm03M219gcJYBRZAjLEV7VsYjXMWiuzMcHPZ5Jo9MDBsIQYaHNpdbe7Rqw5DPbdKEgrUMq7
G0Efh79dkJ7ZNZgMrXEWWIIsGp7+WJT1x14HrGy4cT8T1c31y7suRTT8ecAuPZvNMvY1AgV16jtr
3KqPiDrVoxVhz1GEALVOXeaHWF50b4r4Vm2mtnJuTRFCRdbZwdLdEGuUFEEJFlSimNGWUARyQ/X7
YMxPS4oU6CIQRF0AaN2hgtPMJeo/PvJ5y6/u/HYWBTAxCJEkbW6fUJMda9lwZ+3lRZI1B+RvNtV4
4e0NyhiymaLV7kcSytV6L6VMbL0Xd45vvpqR3aZnLpAOZRMbSJ+vCOeN7JZ43fFYkztKE2APHmZx
m4xLX4GC1E/xTDu5cF44eQHttYDlHxElxHGv9QdSm3gH6KgDxqrIOFg0wZg8IPw7muyNR9fgA9s5
M+sXB2ea6udK32td96/hHusQ3WaF2uoBOjrBfpZq18fpwbBw1zCRT7gAdkHRyzX7hMDjwTp3VAEr
Yzy3NMJwVVvCkZzljmcDsDAhVMub1hsuJKUlxCHkRhzlvy3/SGhYW2T7TDqU4gAnzlN9ysW91LEM
Q3F+KUymiAWgOjYkDfoIEqCnNHIKX9Y6tMnZxmzhTrlFLRMr8DRzy5Z4tpkMehsoV0wGnb5tVTp7
/RpaiTLYr2I5bQv8ZjTj1s6J/Yqt144BgoWMxjTwg3HpYrxWCVCV/zwoXFia4nx0kr7DPiwGeAQk
3glZ9xksp9XMWzBRDyzgXlf7ihYdjZfppRqz9kVAakJcEmyfBLvH+bd9EqSGd+qL7Zn5BKUwyHk2
T4a1tFsMQjVzhuanmvnrzov6sBviEMcKg8mK6+G1zEi3jD6hRPSdYxRVqTWgsoPR+31Bq+PN+kA6
5nkC15Ari/cw8ljKOIL30n9iMT9m0up9SaAGyxI7eXPDWxWE23DUKLiKFB1fCu9CNF3tW/NK/4od
B96CQfGoeDTTb4u6ikAOvELgPfw/aXAKdLqefAD8brJ++ynLi1jx4+vHXfyjCQteV3pHCVhEiE5u
zLHGfsAf1rEfkJqgWVEdqH/c/iNFbyyH24x9/23oj006LsnSsEco9Iief2uSMwOvtWtxd+pYmE5E
BRqCGa1DJfqRUGJYeVNwFmBrlrk6+cQOoqFwIJExa6pKincU8LZeDEbwPzSQcUOfVMAPEnc4K01O
655NiY+D2NtYHs1yP6LJ/33ksZwbp8XGy26LkcxVRjYlplzYmDJoUsleVV1ZkdnWtrKgXKQ6A5Dx
6n/aWVNGMGdn0IObctCXmMJ9MTNw/vGSCya9Uq5ONgSIPJdY76S55zl3AHWLIkn50IfvH04W1fLS
JPtLOwTcOCGpDpU3XFacmtjrDUEUDD6+qS33eck/viBKyatwPjKHQ+QPFtjEmf4rhJVuxeVrrDbE
s/l7F/AW44YHyDxq485X5IRHlVmOxcFOdTt4kwa+dLrUVTgh+CnAtkM4JmbSudG+ydLqnpRZnqlV
MkGNJNLHZFNIUNZ3gmGC2wCwv+mgmCzchoPoN6XYGutcJt76yjL3vao9Eo4hzutnOh9aOqRC8ifx
rNqVVcPR3Ie+pPlMwz8gMKeVdrpIP2jkqY0dFt2MWcKiqHpZicqfoSeMsC0rJBqlPhE9+4YHolF7
hXfKgu2QqUtjE9GorBoe2zS0BF++SzE3nO/7NqQyLOLKbjCqUgJVZdFfHOfx9OB8L/snG25mcNhr
hvoOcx5ykpvLnbtkUUMjjGNCvsz+dP6U7RLAHDm9djvB+1tXRdKX4G6kmln8xEyoQAPlMWlBRG7d
U5D4g98XLtb4niF7NmPv88GC5LVDX4HauNGguErOQ7+/EhswcLeqnnifaFQBXmh/jW6ByVZzLsJO
SkhTSdEoqRcA77cg9L29DjtPeCO4iPejmua4l7+P8MpUQVKCsuBvGGsvmhj3vxCb7gZE/SeGTWHU
9Id4f4G7ZeiOfuKpf0bcw99ta3rbLVVKfqLBDLViQfp3SO4Q5lsl+Juz2606PwI1g9Ji9dixF4AY
lOGB8EaM/2A3jhZy/I208JPZHNCnZux4Qurl6b5J5FLtRocwGOAswJ/DZ8uwrrq3RlXHtNhMFLLF
ztL8OMnHjKEbnWWtY54qDX/KbkrmEHbjDMzldEcK8Ze5Cfndm5Y3ArAKiJpB3+986GPAjBVGeIIX
mdr2BcPyXmajWbAANSZyeNzH+NI7jT+LoFqbZoPL2tgnDjifyP7kMMBzv205K3BooyapF3RSHP9y
Wa423W9eamEkP7p4RfInu8L6CsU6hHPnbw2f/ehCHknKtsey9LoBXZnDzj0PO9Qchg/h7jBLin7X
RdoIWQnvYZ8XhqUNSU3OA8Y2SHjO0Lf+1KKzZSCJtJuSF3yLuVFnnaNN4bxd/c5OR70WepL+dVFw
PpOhZ4yRHYzEq9OZZsUyErI2SUg5mC6NYpmjoD2jd5rRCy6mc3IOLzmhtsS0ENvURd4A3htr76fE
BBhYYK2bHM6S3qPpY8ikczIx1/tPW/I7Jhw40cMurcXtnVE8FDWDqGnYBMh28XnmvrnezSKz5MFm
rxTJkB1WG9TrT9GOsm2jt3aGSVPhli9HRt3oyrhf617ZwFzZ/rPZxhjDXFriHTjbya/qtHbPneBr
W1NGMZiep10j+F7O9DMlOjhP0osimfi4GurbTKOqDA6MFowEDK7SZ5uPcTAA5z/QcUpf7rNXKGvP
5raYmc2NjoIk6KOBWmY4U7uEXUMLk3T8jVHEq0rBaGB9eCR8oLz8SIVswbtSy2B7XwzlLW6bpEdw
iN684g2sH1a39525oGz55CiuSrrKRIHfK9u7TigItrnCMRABW39lwCIxQg4HcrXILKGDmX92JyGV
ApVOWwRpKcE9jWO/n4Kky3fDklotU2iLPP8kvmzyytDV9jmrfvVEr2Uq4XeLYMWNlH6k72/2nlST
InjGWF6bvdBu/wZ3mFfHbtiGGz9jQZ9PCdtiy6x+J8MBfrmzl+nWiWhbZ5W4A0xYV1nKXIbrc+EU
+Oii14Gqp4D0fIP7NJLVGhMkCrDVehk2QLlTSg70Q82/pJ6vZlpIHfninZ2hnmxPKXQDtyO3fmPB
PQtIFLaLipnysKnln80RiwBAoKAdw7rpFx2DsFKiZcNW6nU5LUgbI0zdyb+FVksq7712dktFIwAz
ycdiY7Oxzwr1PB4gtgMC9biMjB8Q2yHtKBg2Mr6PpMVDwX3m0p1wtjldrJinIlkcqfro+Ieyg4IY
IgDS7e18pIUR5R9fL41gjaAqcqiN1UlatIp420t4GkdQr/BjEScrhtJCDjVZVQxRKzkfPxpnOWqU
o+f3l7MEhDSvPcjavsCgXDN7MBz1Lmzd2drpuCB8gS3ccjXnsQaQfhzbKlxhn/5CbaBMhf5P9TP0
I0WHvDPzxwD6/a7FWQGEsiWn4Uq/YxDthU3EDoDdhB9G1dfABJoIo/gMX7jyPymCToUuLD80G42U
/yGYNNB1C5aF76O37WXch4zspMLoHkohXR6KgYqd5qq1rWmWIThy3t5PD8LCu74NeB0uJoB70fKU
kWxC3KdlSZIzief66il4lv58RnBFc+bWKvAOduwk7K4XO3hiABaVjiFrrY0waCfHaUCVJ5+GXp1B
vToEGL+vwGmibDTlsWQ4CZILWnxqHNRmce6KUBe9qJdSalBb4R4VLSdTZr0YF0aqKuRkoIKL2B+h
Ni7z6sU9RZ92KPUtbZyFF4O6XqtIQfqvEotriVRHm1ENqv91/qkft23eXVXoi6Nk1iPiexzc3N/6
FA342U79gwF05jRW2L2iCxxmUMLwzDg8V+R88U9v8etOwqnZMHJWCN/vn7q4Wlc3lpaUvz6v+AJU
SQ70wfnxdb7fRsIDbD5HAgBswomHOxdq3zn1KWUwmcB65A0Eo+0wAs8wJguiQBHAEXZmmrv9g4Y4
tYuEMIEtRZHaeBpUaof4W7p8kYhRcJm17FEFZBkDTD67Iun+xQygvMehztAtpMiOX8k5VIx7bODI
KLDXjj5+RXh3yTuQbuLNEtIi/JcfrkPuYpOz+QDfBf/SFwggfxoXvxsP1j2+0dNLHwE8P8szKh2G
x4Gjx0gZTXYzaBiIn2tRHYLjSSN3lOqB2WLei7i/SUMCvvEoVKPQtWezJ1SJQTB4x2xzY3PXVTp0
MZplmw06onbaSLbdZjvFXRuOAZAeWnnMiHwGxoL0e7VU3IFGLIZyI9VWbUAZrbJrBfer6fzZY2RK
gi7rUzYDUsF3tA0DbwVwvzbJLDOEHrPoDQqGLNkfjWdjUd/y+vY+TgujzBMUOx+ny6N8hrEZ1IBD
MaAckd9dlq5sCsBVUHhqz1LV+hxqSObpz0qr0L+OoVGfdrXqgFynbTOM1UNfeDry+w6RaVFqdho3
iUl4Vd6OQd8P5DwyOPOruu46kkktl8PQjf6BedKJ4xrlhSOTD92ZKxpvNdLyZ+x+pS6hPgZz4xVe
Nk6b6fxx51+FibsXHatvxjSgb5hI7dSVIvmIFDXAf1J3SBWVYaReMsDOJC2OyODclbeYhtE3ji9C
AfZ5FI+/YOpAkIa/85USR4oXy/wjiXWqJJSZRxI3lV0uDH6XEvwKiCLzrWPpVn/EFJX4ck195gyk
qXYh7YSj1fF0UW2P27ifma5jMHazYl/AYL2z669sY5i9grmDWT+4sHLiJ3wvNeQV1HMga3PZY042
SQqGxXqecTkCf171vhCspr3uQzo+tw0arspRcwV00n6rlgKq6Hen1zlagqXPbfG7Ybs9aIlvXxHc
SVOSDUuCQB0C5Hqs/V9PvmRDZ1ZLedt53FilPt8+YK7jTrabTy7Ls3GAUS4GnYpTlSmo0fHJyvcQ
AwJogW62xY5yAfHB8qqWxk3JLjv4UmO8iyD4B3s1ePkHGU5I6JESBoUBWVfLhml+iTgWjyFnkdsB
8r6G8bpywK0s+7JDDrbl+qioxdrBWT7+hLmXuj2aoyg2fJ5gcvsaRyxHBFfAgjCSZfEAsse48Qqn
/Qd14/JShz3tr1e397rWFHj61tz3wdcQiPgFS/82buOto4IU5ACCsYzbrrQqF6o9tDSOYuTCEJmF
vjasUC03tPVEPOjFLRHJuYEcWU2Q5Uy2HU5w8jHmG1MtDrKf46RbeHULrnhi/pRekmbuuKewFEq1
xpqjt2cFzqVy2fNcpfSY2PynM9uAf8cFxeiN3XtnwC3IIFA7Ei78EAXSBS2KMIX5a08C6SFLv2ex
QmR6SHuvtdzNqxgmxlHp20aWavyY4saPkK/m08F1DUn6s57Ml/ld1e35fBMoObTYQh2kbaOClijP
LDJBPkEQYXiKkL2wCgUc8qNT9k+9CEGTda+6T2Hl14B5X6Tf7hpATmm47ARnFDyvE2hSsRRCG3fm
JS1hlVtT+MGYAk/7tBTTPbsWuuMioP9NxLs4yeau0IU91PW88TBK1CsHJ4huxxolTGe3IZXw097v
m9PboEltQe/mL7cNLIC0bMtZ18GyQLAxqOhqdDMzA7zFoOC7eFBur/dUc1jUqgIeyhUx5idtoZ1y
RF3N0YbFZu9U4r0msFA2FnSd2Y6JQGZQIDt2iy+KMezLZvmDTmoGgexv5NX97BO+/Lfe88Yb0M23
TiDNSulq4nKTC1aUBsA5UhVQSVOVYy+JN5HUWmmIM+s4gLnDdu5dY1jZtvnVPxiUbGaweAnDQWwL
A+Rv4avJzS5kchwku0qEQCtD0QEUAYPZgSkD6IFEvIA3RUW45XxwGn/YTQW2UZI+thXiu5iCcBJH
Olr7OVP1QmFzR7kbWmLEWilFraxyhOcnCewsQgc2tCwyf71kl5FdfwVl8WFytkK8uj7Q0pdTxa9t
nlkaPRHdEgaXbRNRle04o/rOf1F+aM2ZLZk4zYLQmwBULtReJt/zH6CVZTY1n52iFV4FJZ3cMDhE
Wxxs2UID5Rmn6ohnDHLRwbXd6+iSU1P73yaqQXsJ+izbu5jg6vvH0vdUs/Ve4K+e/8Crvfmd6XmU
3Bvo+L7vm1h8JF3o4vJoWH7hH2EYgyX+fOV6YiwDcfdnIBinx791in1ASnMGZ1mUd3R7rTP3H3Ee
EFLOJpkoDau227Y4R1ZkHtxf0Etk7nCdmyGuzZCsXjGS/ZkPL1Zuvvr155HstOVPI3GRIdA/f2r2
EKL6ThxRnFTlbK99NaYV3PvCXntjMpblS2LkQwKgDtT97OGZ8fM5WiJPEurMr9HCfjv47xLMV+Xq
099sf24fc5oA/SezQF51ZgAcXj9PLnsIf5AQ6DDZC6DiGRePg4PjHyXjGw0tGNqcPS49Vgb1I1Kh
yV7RRvEAwvYDsOKnwIXV3gnuAQYVHrFfjw+7iihwf7/nyD2hFcceY/OlV+9IFs1THALj5ynMQm8G
MCy0nIQD4D0Iopw8LrWNM3VWM6EhLKdwTEKdN60vXZYyuRAVRHH4HDV1REFdZytYDUKQKFNilbf9
ovkTpjHuAj3QYfZT/wFYic6eSdYCwRNP7eRrFZQe9wOOugQp0Rt2wlDhzFUWirn8IHcGK1MskQJV
D9rwjpidMsFPuUkI/1zrOMF0dMPkoATiohWW06uUu5sSl3xLvCevFLMzREazL/rNitiCKcmfKcc0
yT03j3u0ji9ONICPXdnm/VFAkwxvx3LHqrd7Yev1mkmWqZoquv5dAP/ysikFH1C6WS0/8rDFG1z/
W2IYppQT0kjX6BHDcrIuPkZubVL2rIX6+5QV/T/MhYd7XzKfeQvIBgZ/AnPHV3cZuSGNeo087ip2
O4HAUxYfLyrQq0hmS/1R40wQmKOJtCqAEpP4ypGeLDxXmclVJM5hqKXJlKFiDEQ3Q8SAsa5zoo0w
Qai+iSeS+aOzyrriaGQK/k/hjYWp6glYie+toE4oNnAFrfFnsZhbPRfEq8DVnwdjycagCekPhMnR
sBW7fqnUAeP1dopiowE7Lz2XlNveCz24DvoKii/s0USyEzxxXaUNFQofgdOLWlQFvIUrHGRX8bTF
hlcYdijm/1r8UgwDsgzdbpRLDUvLm8txgRJbiqJTc6gcgys36Ls3iCXO+5IL7o27lSwKiAcaIrMo
PAtUJbCZ9mV/bxdXf0blF5kJ2r9Oya8qkK2U4PslGkEsLwx9i8iNuIz7d9csKE1yi+w6U6UBgMCZ
JMJZNi/MLMBXMLh3rmOwgJlKkRLU7d2uf0ciRX6eOgjMtDK571D9NKlBxXrzzjBcts+qzixuyGuX
YWkMgmeyVLprzWgRH4fbiyJ4Js7ihMG3WgNjwkwKQU6hmHBM+CG9gcVJOmiZ8PCXog7twLTfz4Db
k0dw7Cad3eVtWJ2s0Cx5lYzpgUzmG0fVIcpVw2OCblAv04q/j37AVpVPfoQsrXQv4LQveLnAGbnE
sCFwMES0adBRFcwyDhm34WFTUo5VOk3WxTE7WLjwXX+5YS9HTRqtinOWF7vcUB4rQ2DyQHlurBee
vpw8X3rLDx1DHAGQQP1skLspWRX+doXqpDILmMwFBfX1IaZxhZ3CARuWzFDq8UPrO21yoNv0Ir8P
jaGm5c6UptWAJOSvTmA51NINVFMfs9qOpJ/vrg+oCYzXxJXmuGDzdL2nZnLO9lXWWxi9GNyZaaN3
g6TowbS1YvVvESSwbCe5pY4CYymeJQSEKJW8Z/OR+u/KWW/SK9Iy3y3VvcqKY/6dHswSFWQGinvK
ODbAnD+C11bJEwd7eidvhGqMsI/+KxmbELb4bgH+PyhbDpVZ6br83CIEyjEezB17A8N77KRi417r
WK+MNu38nVC1KTzZNGcQhAiMg8W3d4AIRpLR/FZUEswOq8ByL2AG2+6IdTtUUS5z28aouAQCjl72
OrjOm1RzZQ1LgzG+jfcCsRc13m5TO9VU0TqXYTnhfQu51+b4LFAc6eXq4tj1fx8anb38lIOehJ3K
ac9hn0geFSiuFsmerGnN4qO/AIOCTjr5LZPEOdbRF8R2DTf9qn0DyWRfpsr7VWLMcSy1IgZ7Ctfi
2xThsY0m4mjhVMyLn+MuADy6L0FNDLMQ9XeN7JpW77SnimtacmrnqR71YN53bUmwG+1kb/AS8oMy
hOseZBBuE3BAFBTdeIxI0v+RLgvKkKDLCM8aMA6SiCjbzEgvf9xvqOXrIt6iC//QKmzx+J+lshgS
tXJkRmAGNLG8zs4BYLBjyMTmm4XhJY6JA2POEKSBfTEqtVgD3iSn0Vx/UDHlSZY9bK45AEKet/nO
Fy+B9GrUeT56jqeHJh0PmtoTScAzNCGdPYQFRPYYvZ/Yb/dBIsGI64p5BxLw6xpXkgpJpgvMjaeb
oDZzrTHCVpuRR0tdSo9dzgnlQxV3II+FQz02pA5pU+VEQbK3wxiif57PYy2SN9jhlkKfP8j82hMR
r2w+SPOgxQR/sQJztSpx8U7Vmo053nDnVSs8a+MY7iAh4YZ1lqjHRWCWjQDdSksXl8CrYF2m/D3k
T1BzjYZ+tYdpytu+/3QenN/WUrgvJNBNW+OkxL6MrTD29QxA87uvpk3aazNwQpBPnkLwIILs5dkT
KAQaeGRxp+Y1NbZBJFoWXqELWiu1kBiVRLZpK4kCd375FZ99JQf/PpH7GaL6sTYzx+lOPlgVOkFw
uUWdRnV4Alf0wTR1klCVCHkiZ0c3yoB9ZvwkHfwy+NCDGXNAfb5AbaOSKvDcrAX05Y8tI9FOzVJ5
Xs8nSmRU7aigj+DkjQoLmmxx8xYoWXY08gBfN9F+/9tGPUs1ySxj6mGvT/Idrbw+uHZ54KEQISbG
Eeuc+d98jrBZ0VlcHReIBDNPtaVUDSBsT56EplCOlbRdyxPFv9Pz+wUVI7c5DExOUns4+K9+kMU4
tr7Yu+J3t8/yFl331MEAh90DMP9piDa1VRugubv+io+thdSuZtWAjvTdm6io8m/xwtNjYTOLdFRF
xQY80KqQ5iw/5iNVCpKC5sDia9da0Jc7CpaQXMRFi766RExI6JYnwAmY6siJP/6GfYXwuhnBtrbW
qrLj4+b0UA0eljowaSoTxuse3inBe/VRJNsXvJZq10SJRVpKCQqyulhoGga5fy5i2/qyOWPpl0ys
NIU9wPlud3p721eaS2gyuvKC4jNUZMQe/KbevyvJMDDuMpWdOe5GpiJUNkiHuHqTGUNIZiip71gP
cFa8Kc0Sp89JpmcZ+5H+0A6rh1nXcQtMVPWhLv8Dnezc7s28lZIgDnaor6iCU271ABTlW7uHz/i1
ki7QmYyOAyrG+BrbUljQesNPAcOX+Pgups8v9JcUreHrNH+ZBxbE0+Ig07hcjr19CN/GlUclW9TX
dWtgEC3MBBN5VuqWgPDn/HkzxR4rrcrhUgm3ukhHnv3lWY6bAq9g7EGBlt/pNR7h6gF5DIg4e7zI
LToPezD8DUL9NDLC+LDvUWX/sI6VsRoQDzOFoN3cWgsFfOFy1l87jp+Ls6mgefdn8cKL/X9h1HXm
6C5m89hSDf5v4t0Gx9qoZ2Z4AdXqbkD2RXL5CMnCJyAUEhGkSF5V8+wvJBSK/q4/+9j8GYdV5dKW
V8NdtHriTvgpNwGyREmDWMSKHoJ5suqrV1NdtB6dJwxw1oGv9Vwn9kzJ5tH5udmz8npcjfPq+7Nw
weCrwjUUlCMAh4I5HNrGZgBuR2ulrzWgUwVLnTLxX1ZViyY+bY65s+ECgPzkw7DV2LE/Ghhay+ZT
Oiv9G/dLNbwLEsOcG43ztPds/yliKq0Xw5BuBIWOPdF4gzqGAqJyxUF02sF0IqXEw9On0hZOIfNH
HpEesfQX62QZScGXnVB8tWUwsbkSlTpmZq/acKL7QrJ+gFBZCwFy4Tf+Z1bRHpetRd294PhrsSuj
74a90DXS/QCZ6Kl5dLQW1cca0wR91yNP3K3dAY1iagRsn+fJ/wVCBvroxDx+mMeThFa3/m1byzDS
KFmGmhaaNibboAk5rsnD0PBvxGKATQzcV/vJ4CcBMbGwDoOPevCbte4xJNXFQT6VV9Y47OBYYQfW
bYWa2kwUR11mbq0aiz8XHqTVEnPmvUK5p9CyOZoo462PhL4H8bZFnZ7FcfCjSlQpqEDs55G/kuWU
+SCDk+sf0CT9TIXFP3J2+G0jwkOKMGr9YnX5A46ZSz5srNTsn6ji3KvQ2/B7XIeIMpHiNZPeSg4u
n4fe5PqasDdux117mcfOEoYZ52I/fFT2ynUIm7iVcntjCuUKZQkqtuQ9jM4NzHL0tWZpNljRiNBb
E9zljPdVZfg945L1n+ZxxdSBLfsDOnZh28wJGCfYo/7o/wGRqMe3bdltPZ5l6GFNSreRU7t80VOw
eAHP7aBTkQwxvQyJRxi/3ihBqxhA1RsjnCFzZx8Ns6w/QmpXN/Fx18O7OnhYQJUKl/6WpVftV3rJ
MPLpkjRtwVdtb3XzASJADmmRwPIC3NjSbgzoWs7bYDRmlfVtMK2wJhgHQSKe9iu/hgxvMA2l7jfy
3wZpFzzFYFnviWWiISfXhUCi8UJ7Iv1B/zcZhw/bQsL4XVZi20MAf46ASfGMv9f7030QLhy+HCTT
xwqwmxpf/RFgTtQkK56dnShcPea7cxnB3WR9njcMkPnYx24ibimL7teBxFlLEf2j+O/oCWHu2WfT
QeU0ql7emuKG0CEGB78iw1LyjsJAGMAOF9RWlykalW3xn+dm5/du0gnq2mrLM9lxYyKG2DWFGPwe
ItnX95qn3el+ACjpNsIjiqhB0MTrri/ZxqsNTWFnf5+oJ6N/M5R6yWeq5raVlsms88o6xLIs3o/a
AHYPIkkMnde9RzINnA2sZNK16kiXaUNv8KSMD8JJ25S1j5cBb6azEt4SXdpAkQSAkw8Yd8kKQaiW
RjQH/1/0vYq3fOQjKoApu2D2aPsMHeYnCYjg8N8DZLeO46A4Pjk0YiBsLRWE0OygtWXd3aRksC8K
nmGdcc9nsnJXgzkaLYZR4zgQnn+M2fUiATNLI0h+O6zgCG6cZ19CK4Mo0zaD25E7te+XTUPB1I1H
5ttUbz35faUkeJVftN+PQVdurNYsxr0cqGQ+GGDIUcNt2qnW2eACXXQCCNog+L+ZeZkqysXz3WRI
+FCBzRwzUkxYQ4ij7VWI9k2TCaj5X2xD0tABZuURNegoIWUm8dvwLbgv6TNsrNkEpSRfWafqXgOT
MyUbf+UEsPL41GucA9SbLP0Kt0xyHZomRK/kb/nfgLrNgQMkH21WQF9Zsu2fV7DlL6LkrHnfLBvU
urc3ZPpoNRw3XEstTIiv/xR2dPJL3zNYoRcuOUS/47TOOEumOMrPZOagG7SGu1fl0o3pFs6IDFh7
6mQlBkuGBJf6KviAfoBO2yP4qfINga07rLtESH51d0NNrbwQT9Yiryo5TYqqubCRUl5fXdTdZHhy
L8F3a9xmI1N43iutnQ9OBXHpieq7r6cxR62pWa7H2TMLSUjVD4vOYvoIBuycPG5p1a+rqUxRnv7l
AmbgwMf4GDSMQPny3N/Q2D0R6X3z9pX1rj+yihLlok+HzEJ1L/3ovs25aw9y6EdmcFIvqYmHF8rg
8WOhx0u1BkyhZH335Fa/2HOPF698h9QM01oDVx1fEc3tje2yKAe3htgIIDKGKUWmiUSGHsrsowYN
nAPTblssPXQuX5tYx6SB+vZdQDGMW7qied7tmcoUCnfqL9+LIuSKhRjdaacpJWTKjEnO+0Haqwu6
/1AUdblEuc5G8BHuCP+6xpDUckPwWG/rMjDEF0JQ6Gg0JAeX+j0Y5s+DgKjhxSmXbZqcE/KL2thg
T2340k43sTSDPmNI0DnlfKI/vsqHCxo3ku8yiArRVOa/IJwsbtztib4f+q251IrWi28HcohNlHxa
jtfRGkE2Z2GhqspXJdQKcIFCWV75zyrcUMO5criCWUt75fp4FtIe7Y7KdwwXJdZConfQe/hZaWbe
Kf7Bu/YeAdIST6PNCLEoOEvYiTtLZ3Y4AXWHM1Hy1LjV3JKbXMv1CFm+L2w6DdMrPfAoukYkgXQM
X2d9Y4DcaQRAWOrCVak7bmFAFkKdr2CijiDFiMUNfgnxS+5FKtFbqQHk2JavsXeDHqHZbXm0KJ/u
uel4rlBXOd7ohXW8do185vTneM7J9p3KsAbHvmn5p1zNq1aNfL6GQmBNnt33FszNseh3ys6alTCl
m0ngltRSdq4s+4f9kRlIafLNaYfo3kpC50JpbJDOACCNTCO2GXb1mEc6/XpfVs9owCYr3YMKf3Xu
iyLzG/AgfYpaeeKOufndPcXuqeHrS/FnozR+jNiK0m8PWrgeROiHn/Wg/awfqzvtalCReYCkWlpO
D2aUdbPmpVL5IjXH3yENypEL9BOFqIYzII9BBn08O54kCnsIHEOTReml4S8riFs2rLhNVFvbVN3d
6YBaFtwOi6kb5yfLsOgsk1Tp9rOkRutV8BkiQZnliX62YL27fP1NzxJhP9sxFWmc4jtEfpBxY7i5
vqRU93oAPIt5cse0HY7NwBRIsVX+8zeBe9v8hb2MTUnxbVF17D3KeIsJB1s8MEaYPttEN9AaJGdP
+UFkSbD2SJnFh4gFM0QSzEhqLJI/vS35aBhPtd8ITFq2T/p0jDR4Kc5uVr2PPrPh3LK1XyYNdurS
eeceRhmTKGM1e1C0f7C41TTW538AvnL4kc5O9WzqTvRwkQ2QfYJq/GuRAT4Q2LF+ygEj/sEOGjAE
ABG6iHj54CvuzOf/3v9HTtHl+xy3rLpJgGB6pLUWxfNCsAZ//HMUkYVd0UzMs4/oKCjC+kp3YgGH
IblPY6eUmvJpN0N7qAfb7dPoJagMAYUtpiuhK6WbCeWKk6oRQ4jmWX4WkmR6EwrYktw1VPINbk12
gPf61F1rabrNv3scyLbdHA+tkqUmI0yBJHUtObzXxouRJRyzaRZb5mlMS8CgYg3Zd7SfRI6vQRkW
zZAauFl+rChzKQMy6l2JMHWcmgmnzSRDFTojMyOEq0C++UrtrpT0nT+H1uu+neG/Yyw+MbAg2nVJ
+XCA57BXnsAtHwhvlautZ3xdksmlPz5yF5DbgaDgwgPEqIRlqeI88KeBKKvkTnXklCrk33Nj1BK9
y4miuK/PEICrhW0kzmy5/HTzp458i0rXUPUIdZXnL/DJvpBEHb4UrMl+oxq7cpFlgIXYdnneMm0m
2Y4NNv6oG86IwJaojJfR6Vv2JmnxTHX1Z5EfMVwAaKPnq6bM+xVHZo/7uHGCRc1zqRYQMdEpBtvc
bgh7aVA+c+7r08o4wQn18qans5b5AspvbisWCTG8OePsZ5o1DD+u/U6ew4kcLpzGFtuhxS4EbzMu
GsYuwpUo8KFOI6bU8Hior3+6P/+PID45q88IgcjTxvqeY2zOqhJWQsbwTCiIi0lWguTATb577WEy
JCvbSA3dPBIJbC/kqzA1fhTtDtfi3uJkWZJBPqlFecCVWXVNlppGZO9WyVJnrlR59y+tgrpYOnVP
Al49adqmUXnouUtw9FdQmghXoEL3ogrDGkxlL5eQSaQdP3wCKzRi86BaSfGeghiBcCorpR8Efs68
fzo5jzAHk44Pid/wyK8pFP6suFyiYPG7EfJExW/zxwk4gGutLjIoAFHc5foerdOdMAeEIcr528ru
MeqM+3c/pZVH6cZ6fzaaeKqINWySOXMVF5gCON+I3d+7PmFcCgX2x1zkrYDfSVR6PpsIH4Qo22Fr
4Rdmy6hc//+dSe2LltxTvSZgTpI3C6VnlcrlSPGvbP6AIbhtwN1s/PgcnpA5NEcY6eecDjJnXqMt
KUbLlVuLJtCxxOfB7btakcJKfB3ikVykMKkqmoCJcfuPGm6J2P8UFSdEr7wn0sHdP4hhMX9KZsGf
WgzL3FHsO/ShyXv13Pbk6bvW8y7xwKbKRWgq7jfrpQI9LUsARZOV43IxtU0FJ5Sg7pZWEZuDuG9I
llcWr9yFjiGZsUo3CG4N7gjEuQ0PMP/QQyLlDed5W0UOMT6k64dTb2b2EPNLiRprhOwM6sCzNKwW
LzsdOVaWZ/WU8HWg9OB6y0zQHJQ1F1C4pBiaRc8rk51jS+NXLo5UgCOjrA9wS0fF6sRQf/Cis0fe
7KQS2n1lEsttRspFF62qRfwugOA3WOsc0KsozE5ajIvvYml+O9cidRrq0Iir5IL634rX8qZpK5ce
cNnAI3+k7JrRSeaf3hnWxPFLzYOIgwDKmEuCDhlaBrjzphFYh7v0NXl+TOWbACQi8kJf+W8FeBsb
MXM5fEv9ljxNf6m1jENRWSlZd5pdusaSfU21MS0G6GWcixY6pGMHnx50h8Xd+hn5E1rzp198DkIQ
gSpHlGn10Myi++bFhcPDwVGU7SmT4PEmRGpeiWLwZZtnkZWBPFNjciOfHQwfjsE3kztHhCb1/B0n
JJc8z+Iw8kIa8QTcs6+SZZRR0KrZvdUwJ1A0DOravfN780MglYy8r5kuYpEE99g+r7yXiELmBUNo
HmXnqxu3MwNgeC6FTArFba6xFx3Gb+n2C+fj1R6V27MrgPbOYQS3FWO+SGe5PX5qlJWADJbGzJQT
R35enTYM08a8bsN7dUVE2nrpDJNQ8RmndBh1yugEmkHjB84Q8tyQUdN1PSL8Nj40jGBZjK0CZhce
/xGdEpTsFrDq+Kw0bDtxxAMhip7G+VWvwvnNTnoz1PDOz8IBEebGXd/VtC4SCeN3wVbNdnGm9XPM
0KnL1a9cc7bNutwe3b33226JPjnYoJ7Izd2knE20DSSZKYGMsil5fhyLTMWaSqVtRQJJ28BrcQFX
Gm51fRiXmJSQlviFS2ylEFBJdHBKDSHW0MmJWfmDqP1LyoZymgzXTGnoGo8sAVJqW4XVG3bRiETh
C/FgSB6jTpIBRfzeOlfw8arveAQZaC0uaLlEptAxJEXeKZQxa74y31wYy06BNxgIyXX4uXFwur0c
I/m1w+zORNnDOhNSi5IjcLfA8NXI9DmsqlRIemdySF7vUApBoeqKx3yXJG0LePyhV7xt3yy+KwcQ
rbrXSxJZZAQ+fJsy1hkoRaGllaxJtQXXuVyl/5gluX/cPfIv8GkS60ln9Ffe1ig6h5reXECuP8eK
fFWFyUVVLyKuncrMEzdtWS1Zmt2MGvacSmVNbTX+GrygFIOId6YwtfNXZiXHctfBMcSC3WoQzjvn
mE3CzJa7geKVDdJym/sH3Ka2JUIqS5DOP5wJRN29EZcISz4rmUTssG4w3HBuu1pADHD+H3k2IbGz
bYmLrJeeFZ4VXtR7yKNHX5i8XGowg95Xgsby5h/VcteO4F594jj0sfP63PUavKZVqobY/YU9gODy
jaeFLzygjuFw+IL0+N1C5X8ikERQ0o6Lj9U/yTMXDgfUjEAyIID/4j15C+gHEuffD6FRj8auQPnf
3IpR7C//RcnvM5jjPp1NZdnx72+GzHN7axK5dhcTuf34Ulyq6s9M54a1haEfZFxqk5Goe1z/S+hS
ulzUTU1+dET9z6vw9OlFJJTe9iG6HMOZ3MrpJnCBv1LlVEW76wlzFHjm3iAHYq0t3mykSY+QwvzL
Qh/slL8uAsnNudd7sUAAjf6N/sEhCsbmpghCDRsn0Aboix+L6km6wzKB3CECS4yRNmeWjTVD9Z9O
xm4btYgWvf9mbD5nGwq95ocQKnKwQTshrF2+yIjULsHfwggO2bBTXkfUh0+dbhyIpfWaVHZW8nZ6
x65jR8LSDIIdbEoHVnIqqzBJJNJ+6nMDbX3BEPWSdlrscn9SO+vALkYTUpPrRUIxdTveqic8mC4K
TPGbhjPIaj67W4rk1pF4o88ItB8fhIay8DlbcRZ/20Senqjm7P5D8hWHjuVoefegMtEbTNH0/WCX
UaOztDbrS2+Nk89nY/qEKPkd+W6BpITlRwzRX3lsRSq+fzSwniQnILxHtHubG0Vd9gqvTbVWBuJO
2Wu+Tr7JN3fhhv1A3OyvnKyFPs9XCnI6s2DxjBsacuZAKzjwS5RkWWNE/ItBQiWNVdlkxbiXMEjd
TuZnLpZ/P+0bfUiGYKYCjQKSP7lFQ2t84wNmjAuj+eMm6CFpkXDSS9p8BSkrsouHe4Ydf0nK177H
PYFfqGDIU75gHC8AE3HWNwPDNwpqNL0f47NGNox10scgTF0JRBRxyGeJPR4W8XdWpdJvMWoAc0iz
veRtNElGjPDHLYU3EuonKmBko3n3TRKBkJXgylroOxGkjh9H8xmK8PGfbeLq1sv1qds2UH2wrk0s
xOdvBMh100iqDLi1p9VmlWstT/YmHHqsKy5ZJlOLwtrAX+fZs53teVwojjzfJbtlD+4K3LW8p3hW
i3/cUU0b3gPOdXjMVKIFUJQYbQLr+nxxIjBlOFCHpKzwatiGVGxTmowC6+9paZCPPYXpuB/yiWqv
avTf+sVn0rNmLxKx6ady9JO7H79iUw4SRdDPLfTGsW5/wMzwyGA8epWnBi6LUrRIuiIATzj0rkuG
rKhp+qeoIg1Es5dPkkJjG+tFlStdlUdXEsPmMGUhTQyB4F1clzbiuNBW7yI5UqkR1DkB9Y2SppgI
0Z/jIoa8DpwNWf53bspdwPkTBRBGdyMd+U1viIWJXJZ8kYLM10vl7scyEanIqR2V96DbpR9RPhjq
nCbfzyiAuUbeyHor96ugZiN6rYFK7PRrmd45c56+JO6Hgim9JP/8keqOB1N2rUnbvzPai7laV3tY
RB5DYf73toMyOwVw/RGxJrGA01plDS00eUu7IslxErCiAc7EjmZzccL0WsYyWUELtV90wUWWZKe5
D5EqWIrZh0e9T8i2sKBcSYOVH6gBJPU5Gu/TDSlPrI6IEJ6kTGUGBnuAol1BjQlJ3Xg0U/48Habm
O7tiIGUsXqntc6BZXMSGPhp94631/10EFXgu6ziq6f2Y90go17afcySSrl7180Dxf34Iz5kvwudc
w4ZZiX2l35sDCgX0Okh6gkWJBHQc6aS1sQPdKAidhxSpYfOlccU8JdJDvEKjn9zRoXQFkYTLzGCB
w6I+TrucxQhBNpfbqv4jSyzMC9BXlJvloFtuMujcGgJ+qr7JZyzxB0zHVCuhoWwWHoAu0V6djnyF
kwBG//3GHC/QzlZ4fAZkT0oDpO54oG38Xn5ErlP/TxD9LNUma/prNRkoT3F2SJeqNRldxeeYMQA8
H/r8bnLs+5bcrfR+FxPMXtCmg4UTpPD3PzEj2t09EH68XHJfKjGPjgMsY28pwxizf1AUYHw2KlVs
tUYkeYhgqXRD0yHRb7I1o+5iXxKG4aWNWnenWxwYoCuvqr0ZnvPyvJqP88WqmmhRJyP3OxY2LY87
lqw7ncUQOzrnsEZd5vUbNQDqhMNOETOiU5Yr2jb9yrLQMfuPRdBJxolyMI0JyBj9E4mUwPWS+gkG
8t74HxZIyT8tfe1YMBm1Ilhh+e0inFY9ZxXC1lSjaDX0tFDbPkdHFT31MkIsJP4o2VAbel//5DKJ
Bjd8DVtQ7PDShxv8zv44sCU2ww16LWkRQfMEIWiCTBFTbpmKSN8runBdlD5yHG3gOY84TDO9iycz
BOslag46/m3A24bJldTNKvmOX9Y8lhHeZQliIvmcs3ASn6UPJUbCGuycDQhnRIC50BUDOpnVFnXP
E1H+uEem2oZrErKt0oD6/ytLKDZHuIIEnT1pVEvIDGfCStWZqmWmjQwsQF/oIxwJQ+Q4eWoCVaV2
bXSVISmrPfjNEjV8IjTNw6tILcm0PCzYQHXIxlXC6+xzUXDwSAzSvPm1b4svJ/YqLyzxEf2kx8lz
AQsRCrTaBStdcj0XpP2evKo0v4O3/5bLjYKh9slsxQt1dAJU5pj8ZkMSTa4rIpVMICQsO5Nbs/bn
t1Vh29jYOPKK9QKnfTN3idfVkcmul97d9E6aN/kIRKymPR4BEU4MsZoZNH/F0UExPpzCzzwGq2I+
AS7eoskV1ggJijFJGsMcIo0bnK6sgbxAjx1/t4K/ceSOosN92OnTGjELZVqWheFrVKj6nt2QiNKm
bljjxg/5VGDOfRLhfChcpric9oVKG9zlhi0q/5ihlOjPZrTpkAP5gSpTHtmULeVNIdOS0qMxr0oR
X9KVjsADQ/gfpMhVqQ+o5QQgI/XhLI5dO5DLG0O1NcfMCQuS2rVchgKEHRjrSsvN7VUWKs5xFBSt
wwkbHzPrQ5v/yWQT680nvol7XfzCovbBsWfmUbUofgOwEnxUb594wEQTZ+20XhQANERYCxhjqjHJ
MWmgPhgrGdaLbLkD5hIBRoG9VUJlfD2Zv5th4J/Kf5mldk0WFxUzZW5si9ngke+QEIIacQLO10Ji
/K7NXKuzORaFb4pOG//u8hGbx5nDAs2a+YgTqYjLTMQJmwVYdo8TXGD78BHrNxRfgufxoJ63dMkv
VPHPizgEbuF8qE5sosybuqPYZ/yQ06yD1K523z7nUW5tYMXtxkzEb882I0ETvSCeA0Owqt+sxiOW
HHokfNuYtzrRHsKmUV6eukF1s0u4BSzawx4SpskcG12sGVNoMtAclCYx1mo909haMy2Aah0GTCMv
XRCQFi3WjHBeDqkKBvZEfNHfGMCszNzjyaC9AoqaDoMPOg988WJvCDS7eh9nceqY312QpPaJKU99
vmFmDXLPZK0ldxYPiPW8+kRvclFCMx7UT1rwRIdSQD5ZPiwBQ7P0I0qT8P6LinixaNJXDVpGfQrQ
qXKyPzA/p7ThWEyYYqebZWcwZxEhjEf/yC03ebmFyh01w9E+MuQBVes/s8GKHyCPYljtacBmGEdd
3nGdQZUXOqPBtNp1mP+iIIHu21KJmF1/Rl8BjVk3YVFk0dL8hOkc5P2lXIdwusk79GDH5mTcSpwQ
+ycpPEcVQvZ+roGl/EbvIhE2MMH9llUYf8OUTLhfYWSLKHd+r8Wtyx7qt3uEp2NauMapSUqlriyk
KzfmUYMn1XcX7ngvg8an3VJtoONdw1aJlb5kxwbASoZul+N9DweRaAOdlbci4hQh0zj5cVcN9cyQ
naEozW50IjkdF7WLkKF7DKRMDcn7J8h9MO45LF5Hng6dHJ7RAYMWLcd++VzkbXjhXC3p870nkKvl
nMBTedMPhd8DzOeBYMecQiR9ttDv6amgjY9sw74HsIQxsiaDVG6tCOirO0i4oX+6iFL+6a7cML4+
WkJ8PIRFKiZQb/8Othwlg2YnhEJRLvu437GMAZA7QW8Wfo2PwcNicDK8H3D28tLgZe20UTTFEcW9
uwaehozOPtAxm1HVEL1uPD3MFDyrb2ADr6HlGQKCDMHiJKNX40YwDwarILkmlHRBP94GG3sbqif5
7vjxAb/HHypGlwsrmVc/ytwRsvmWpCGJhCmfsOahv74yX+jNK/4ke8Vsb7yPT7SU32hRmi5H3rAz
2vECFtOCFQUH25XRBjLSiAXZLKgMf8HjCly+GRTUHqfedXzrzscJ9+6Jz0jF2eJ1EnB+rwbQ/S5d
Q0dnHjuMjILgJOdKiXqMmwPd5qv90TXYUhyrTGz8alYoTnOFdnscyQJ2ne4Ew8oevByo0ZELIN5R
I6xbPvZiwasl7cPOOcGyzr8vWcYPNcRzplZxDF2jLPKnaE8p+y1SHjq4LRyYXsgARPDDB4T7QVpZ
vm3FYX12CDtVagzFuEEwJDBPfrG5P6ECRJAYcxH9j4ZdBczuZKh/X9eDkDN6jZEM1EG466QuEQge
ro/5ZdLdSjr45QZOZfd0D8qpvj7tARkD5WMW6aX5N4VpDYBgVA8ZQ8KJokvfWH6jt/2anq5V6vXp
YsStKIW0PWOSJ1W2fDDZwwlwwchOY/pWj2A0XXn0KFRQPbaW68iKmTA1o/t87xpnfqEl/uwb1RAl
c0QopMSVcsKGExWAbtKqQ87rD8bFkrdSEPAFIyYUQzqbf3oDtu2peu9kK+9VzGRl4i1EdLr1drj9
8nsUYJO872kaDXByCKqjgVMJIUyWu28G5GqUrZCXnyS7xijrYHGSllTUk6/TOoxYtY7GZ6HBJZaC
hHHWttXyaEEjxW2yU+BSsKObzg4G2EDNM9TTehj7xWVKJiYCFYbsoU4dyrg4/pyo+zhpaTV5VRXL
jrglVeP6nb7sNtzJDEE65naond7b8HyPpxd2bcH2HmchMUtH14JxGsdv0LgzSBrSxbD9t0AT0WKn
36ePQkFpRxKFJuBs3v/gbeA9L/Drl+AlLr6hphF+atoGYDbqC//1jKLBEwbpr8fT9e6b02NPs7G+
gaXsE/4Crpx5hhn9c2jtAyMepBqV6rFNyHEAKHGVATJklu9CaqFIZJ8BzG1Fj0Bz7weop1xcDWW4
7Ibd2Geyz6Ddn+o1Qt0h50NUfDHoIUa4q9VOcvnp7HmpHLTbjg87aqj29mktgzQvD9BhBpEl4TFO
QnIk55hCl9d7Kueppd4tE/RZDAn9JpuvN26wZznmWVUOYjGG30he0wKKIQew+fRGLkASYDBU8ziE
RdAZETbGYbLBwViYGQsTE5oQVsvrBTfrbMZQqmZxAbab+xRZ/4BjFt3Gt0F+4DkruHvr5XpA5/7/
9pENqfe/AQNRgFu+krPkhXSGXRkoKy74iaYFj96iOjBdaCPa1SK8vJMePzv+9lta2CrqB/ugP9RL
J4CP7zzXhvS5y9evwkSOOOUs+zU8PbYMCQqhIGLaYQ5cRimw1+p3vvqVaNIW/kgwfGRb+UX6BOZF
nKIVEYSaQvhdd4FgF28/R/h6VVWhDioYh3koCE5tSnYoQM+LjrjMJbM0rmYBayw9CBVv4jPkyG81
sUihq+6BM3bVHkY//H/yqetkgYbBl8jHGpkUWejS1lRa1d+8DC8IHwfIiRfR11+NbGQpWnjytGrV
Izl4bJrvmbO9p9jSuyyD1CsLIjOAARRc93F/3G5Ixbxaqo9tKvYexFcfc5VDlb8Jd5qmuudxWZWl
I4etnqPEc7R9pOyWVoqglD3HkoasW8pWFoIQXVJlZ9fm4SxXDl8y+F289TOf21KXIBUCa3ZkQZQY
cbr84SUu1psibMIsUFrs4NaCD2bRqFbIeHBr7ErZBd+PkAZZAPPkqlohAFrr4K5v7Vr9Y8HHQMYq
eG0r50o27jyONJATwP+bNj0pGqHN30rdAO5sNlTHZap6eyeZ8ANXEZyYumJyidsL/z3gNNYGiCHH
wzFam83T/eQpden5zFjLd6up4TQXkZORHM1aXDaDOExHztHwW7d0fTSf2MCfANSx2nr1riEGkGR4
0Hd7P7J/DlnjwQUTPFbFTS0PPJ+xMQphV0PbR/pTzkhPbApvLRqp6e7CFxudzbdmRwDO4QkRXn+v
U36cblGoq7eMnmBZr6C9Qx7evl14RWKxocwsoAiapcturJjB9NqDeA6Rk7Ged7rwb9X42ULSE7ch
IJo5Dwdwb6ROqYjUbzgfW5WtxpXf9N+XlloslZOb2O3354GKWKzY3QQUhwc7ZjZcZHxp2vR2vBpk
vkuerrIZ+dlYgwXkWmWfD2SU6PF1+Z8AdCm/C5RL28Pc8VBxcVYRiwhpohQ0OQXp+YHQL+T0cJDf
1OpfQXKgr/J5tWZbMfS08fAc11MXMVqUFjJxFfUZQu7npKLufiL/UFMDNuv2j99L6Dholj4EYcGv
GeakGFPmCzjcp0mAlroFr5n9vOgs2PH+3H1/TfCVqIpSIcWflXuaTjXgXQVxNEkk0+RRxdhuKKUo
jx3/rh9xjguU4pyi1/B2kfdO4eAqHD7Txi6CBJUOwjwHKQQ9AE7FAJTzdx67g4jf/Ef3TBINQnWk
g3xsLpJLlGeMPI++HJEw6UTx+j0QAMTJty8spRYiOXXddUjKnj2JLMIxCqCL5kmoNUisP3AAOMGL
rileKv4SvefnOVWGEwK27o+9kY5xS7A++xC98U/3AYDb16e+VoLQH69BxlH9CsZsfchgMxnqrfTM
RWGbmVG4K1F9AQ6uWcze6ZQy1CC6EYA653uuohhJnT1Fef5/ykF0jzqDyO3cIfydRuQ85J9v9Ulm
9m5jfY44zc1toWVIFHtBxctnhwLwLy0K/I+0Gy/+RNKKVzV7OqIHByYxaDMPIqxLU9/OsGlOr26M
bUrIfXr8nCcdp4iKGdx+VlKiVJ8VDJ+mDdd9VsGpVJ4alinM0PYAldjCgDP0RQNJe0zT1dX3ivsx
huHZO1Q+0tt6mkuzlTmVlYNhpwK9VhIil8E0g/SZe5vUIp4jGqBeiFpJDwLCmPfRMwueMZAlXXWn
9WTWdaDGFdTBC2nbwVhVt6zcqtiiaC457ZwjyYNeroyG+H5J80bPLW321nLNl2EIiv8uPXqKxPnD
JM17yphYoaOUDN4l2qpDmJZT8TxmOeqkW6+vCP6k08OEST0GgDlVpStZbKEx1T/AoaD4/HBmCzk0
00W5E8kr1/SHwSp69rdiBWYPLoYKKND39Cpsuc9YZr9i66/rafU38WlCrv53vHPUwSPDUMvr6FpP
UQkF3G8p8qPiuV5JPDgwsX+Dn9n1S8atXSQSkgYF4WkHZn7nc3fvRtXKzoxXQ7zuIknkOlCrdP+c
Mf+pLNHOxWU8ea9g7ubWbi4tM5iaKOWtmGuduMZYRWO7oqZPLk0f0uInOeYqnbB8aGWRE4VH1cmD
f5PCKP/dcu/XnpKoNr77YWFI9SaK/ZU9XWOPVtkjuV0cZESq8wqBwJYYYQcOKx6mbaSROjqFMca/
yw2BHyDZZ8rI2HEbNuFYIxAhvZ5QLDUIkCFPGHp0VFSM3lMj/twRb+WHAvX45R6U/hWr2s3tmEN+
xDzWh+b/QKOUL9U7jyl67DEmxnCBVaRzmP72MOXbcmsQUxahYwr1S0srcZWn59nzAnSfiOBiWTK4
ElHrEMKog+CnOmhZbhGeijl3KXfPVNAg6fX/82iBrjWMLx7BEVy9tA0nNu0MaWkV4O4bahZoW95R
AXxlY74w/Rjgdk2g/fU3yqz+wnIQ6ZXJ4PLNSyG/1foorjBYlK3Nwqkwg7Ehk2yiif14HwZrA0FA
hTiv/ptB4JPAVC0ouNzxDSIQF2ek2dnBy6X7GWC3f2Bb+lw3vDWo9HDPXLgsIGkJBAMJmcHYUgQI
In7xq+QNwpZ3R/bPKmwK1qt0vhP+86YAhs4LKGsbSsFbXbjtPMu2f5SuleQBvgBF5PGSdyf4rcjU
f1yBfha+ObapCyzQrYSCmWW5a9Y8fsZg6tREAYlMlcqI+oLpsLGPvvlCL0wiUnTNtAieKheEh6KK
ZAvP2YgpIeYLn/gwSyY9+gb+kUMvsxHPaMwteZ5n5xji9VfBrkVVkPgJlqMdolnZ1kFJ+FBzEFDW
gJn/6aXCf9bwmMxGXOs5rRzSImopsAK7dKwxmz3TLYUmRqUsMvqKYgmi3GDcRGqHdeJ/1TbOlWpa
hCYYSZ0KS7Swq9e4UAmGXU96/8RLYaTuF6i3YunhTz2F7gt06cn0gNwo2wH2zTwXC8ppTzsu5Tvt
7vbtG2ya6G4ilES8Q0mbFm8yuWBJ0zwYfDRmx+t/oJa8eKNHbZ7Qr8onE9ROpvJuHxokxSDqpTLT
ZaGu+pQYRkzDp1rx9USbnTSWyBCf/2qGgeFwQfGDel/AIemojPylXkAQEWMRWOpM75mx9jJtKwn7
lnzVz7S6WXMgfrPLPqq+kSCOMD2zM7RDIwsWwSdryfYEBfwW8bcjJA84coL/RRH7vYZ71+e5iF6v
3rM7cMHRv1zgkHPh/qqO+Z/mSXxeQb2TCPfbYsGedmlepAMyGKWCx5aehZeOx5byUT28P65+MIpW
8z3RQkwHPVVUdgY2W/MME0I/RvH8HLEiR9Xli+o0n/5xCbBdQcOL9n1FytC1tK6bvobLCmmKXWEd
AmPG8fGs6b25OoOobxRHOqdE9iODD9hRj/s5UQzFCapcYIbcPHEfSAfyrtaTGadHJ3hDrWwcGkkp
LnfQw46VvODUNteA/qB10vWx5//spYk1z44J0SZap+6ZOWi0xECUaFOuDzHCMcuwN640SYUHqKjR
IRDyL0aAk/jKUtFNsctYj5Divh9BPvU3Fxebx9/zj6w2bgfis6gmjWwcnpYDwfdmySomWfd2mCn7
kZbXIJtHuAAInC9YuF7PqKVJQ4SnmIjpgCqx3PJnv77EDh4yyuPEvC0wWiZKVCEG0GIYab4TLfcI
3ZxH3rP0FPG93i9GZJ7K1vgQ8HshtRtBJA4QWDhxXz8SU/w3AazHEIns/8y8DMBALW2b9BoyqcBH
313TPlvfVyeTm3n1fXSkJbQ8gS+HDGvNMK7wPb6+y8wYfC48FrIpOc2ac17Ir3aw5gUTqj/6IL8W
ZKsCCDsq9dc0u8hJihL7gm+tI3rbXyaFD+z9i2fby84MJbnyZuuakcmeKTSM046jw76acuP8PEGJ
flyI0PNS0G/WqZaqqQZc7my8bb/TOhhluBxsRJmw2bRz2yGUt9wICPB00DAdJeGm8g8eNsNT4aqU
+jzKm1l+9u6N7xkjh78mzqdrP9T4F6xbPEBYqlsAavLLHXi/oBG0m87RrO6pJfXPbNCyQvsVRmsV
Zjxmk7F9He5UsKN6UzIYEEhZfFSmahwCpRPcrH/K+MIMGZMB/QUl6W381CvCQ0s1wm+2RP+eNhPe
g5qP8C2O6ZgM3OQ/5KoeV4+QYGhrnFiQe0E+yJMGMJ2IVO6ysAlC5zClJxrBLGtGG1USmDknnOae
xJOz0zF6MZjcB+xZXOHAnV6donXbeBtTAfPFSBc+amkcCOt9Mc6iQxb4ZqYg+F/MQ5bDNvu257Pi
5ysR7jWeo4oi3+rNt5ZZ4faRZrPHler30H2KxhdhKT7yZSbtig1lRF+232Q3hYjH9Mu93sHnV4cr
Zx5VBGs5E1AjQ7e2X9PQW1rq6hgT5gtb+OkAecFnTsUT6cXYusRCMiT7E05JrP2pvVlcrVz+TomX
zvn3IoxtJV10TVVI0+zcrj+f3wDO+EOo8wCZTGPNaQQQvpPAQe1Rgf7MEYrpxp3n0oj7iNwvS+hA
4PlAQr/xUQhbGMzSUaiKBNsXKRLnEVT8HEFT1bXOABN3+9uRmkiTKA6R7d7KtsyC/HK39tMN62Uz
G0nxkCsjgkCPmbJn8NPzEWwQmhXWs8j/Tc+sDlj3KX0/6E/C4lAUrP5UD0JdpzOvAU1Wal4lFj8E
OGQU5agXm3McYagUIava5A5TDO+kTFjJWXmbfI2CqZHe8RcRObxb6jdm2t/4M8h7x7ysphKyQIBU
oyUmXLp3tX6cqzWKkjAYrBJbhJDYFs2EljdeYIBbB9itji/yDRraWrzQFAsWL0QNYse97ZMyQhlU
Rr4q5edt+LiRQZhoQeDhuyMTxcdAxVvfMkrqFSSEsPs6/zDsUa6QHSHtcwTZPQOcdF+nVfHf1tAW
hmjEBtVgftYAoUW/7/vXcOOomGVKsXaBC2PgpOU2aRU2U9wiItX/vzfiSaJIKFjan3ndobHy1ZMb
+QJPMh+oP0fr188aSb72kMeu/+EwHNQLPSxT/Q8mrawDRDNv/yiUwcsF4+0HVr++N1snTu2CExvj
eA8HYRvqhSpv5w/IDNT4KJfEmV2JHUEz87a2Y8anmXcRZCQk6cDhTfF2pXRTocP3q13dzi8VzQQa
1ZLbv2q+cu2wUlBcF8znG8Pa0U2fgiinwAvzSQ0mmY6IyslD8wbdR4WjAxc6mIXdglD/bkuYXFdo
nHQ0TgX31fhomfqozf/CJ01qNZTYcSBfFP0xL0Tboq3M3ObtEYZBwEmhxvDq7nl5/e1zc0/5FMdW
3VDjlKBQNL5el8IqipZv8infl19zXxu5cSqtaEzNJGkwlg3Bb68L77tyehsk4UeI0IWHC8JhSo5m
J/Mz1WQtykTleTF7EU1Sv0W19IuaoIDcsXy/ZsR03kN1BLDJxMHYxbbGdXymLluo6e7bIuyyEj9C
QHzq9H/dWhj4Z9JB7ry7a73w6gGydP2Ms9TWP3XFoF3HIMqPjqZb3A+SdigiRm+XRqwqeGnosyHN
ikqsTZMf5XZMeTLF+LRpWQsnKd22K8lnLyPD199PkiZlY4g1ZBxFaB/0fEJgS8MaxLygpMXqBZ6E
MChNAAVmK8lgPFQpWrp9rXQ2Oaha8dOrhx8YI4XxKQ08E9OfqUQGZUuNdUo7nQhM3jQA6kj5vO4I
KOVUjgnxTZTwcxrKI5rpm5LAK4JOWJiY6ykrMwYDseOzrUzm5aGSeigjxc1WX3phlfRIbXoRz2gl
+iCb87TR/JH7vXS3axxBE1260Eg1nmmZkRenbj5TEoOZfMiRI/495D/oOwtOVbgwOb2TJavY3E03
LhEWVBItF6VHtfjptHAYV18BFLOriFk/WZgux42JAb7fLUt86rWYtC/fjWK7LrmphGmAgc6yQ6yf
Vz1+BuRZvdPlOmiL6wf/Wdo2Z72mx8dZib2ubTlHJv7Ca5tqan7co+TdLQHVHPRuWxyx8TDkn5PZ
Mw7ry+ol8ODI8SB2qRjO4jIhbcTUjfu5lkI/T8gdRDQ24mQZzx6pk14nYC2raFHOkA7Yz0xiCaXV
tuAu8EJtyDMFLndpxciADN+uTTic+ZYtp4FrMIj9zEhB9y5hm0jiYBOiEPZ/GXHLzNCkdilnCY65
T+gvXpv6/THzvm8u7RAFsR4Q43+FLmjU40cS2YQCnh8En1Fg/2TKEJx255aZo22buKwSzaUIdMSL
FECqiZusftK18gZ42I9wzouxiHhIKW+R7tvXusfzHhDZmr/FxvnICBt2woWUSucQrEj3OoEksWMQ
DUApSUMGkfItoeqUn3mYKhIK73MEDeZHxSgnLlFKbpbbuxGWVEMRTxrHeawftbFAkvAQ9mBnG10R
lAHj5gAewvFhnP8dt3TfmkX9E0/6Bf4ifuru+hljvHZURyhfSE5jok/dswVBBi3XnE2SEqHuLP2q
hbmfrHA5ZEIibVOALJGtt2xk7EoZaHoJbDhQSUbXaee59mtTXNaYL0U6paJqXNwNRO7DgPbFrn8b
4Sauyy3CKJNCEmkhitYb5AhSJvh8Xuq/B+VliaKzqD90GQahtvHhk6xbP01wQYb6pxT2lPuw68Q6
R9C52kB1OzYAJEXQE1tVJaLbuyem1mO7NZfcxiQsZaMCmca9S41xvgO3XOs5uRR7NtqgwDAldw32
y6m81/ylv/GGEioKwV134ZLLU/uXtcp1Krouxioj62aIroh7xAf+iRMXqDj9+Q1Hk5HmOyf+ui4K
kGFVZnt/hjQxihWAAdKyMNNkmVjLUIkipXQ2V50AKyiMiv+vTwKjS8aSKB7C4AIPJwse2bnl2jd0
E4GwXD/0dI3c8WooL7HC69Z7++WTWfcReFbKRdV5SOIkSd16KZNwZU9/j0TmfVIOJVxqyuZcH5AR
XeSL0b/sEefZnpFP+aNlfclVtYdGbk9ZRTadmNj3srOZUY374+hbsc0v0Pc5LHgYGTQfpG4unjiC
g9pv/lljQwRR7Ilc0C+5QTBBLMTQotDkMybXBMMFySocQd7Oz8mYt9gJHmpGL0GFd8tqxUq3Q4mo
opjuJEqBxCmXXsGXRg6VYyVx9VoYUXxBiEzcTjVpv3KocGCCvUBNDMG1jcQOepu/zEUXWtknAThe
pNQjf8Dxn5R6+imTE6JgNHYjvxBBzADHax9XSNZ8vEvylwvN5PKaAyYs1xN3r+2yY2oZdHJzij1T
iRa/5OCG3Fkgm0cBJGGecKBgthRvlkWRdv2OUdEtRzpAzLPlyXaAcZGXi6dbjt3V4NvxbPhu3Osw
WrKRqsUZ7L+S8RyiKuS3tl7lIyNSnw+otNMVv//PmbxlCp4sCmMRa5gnvKUGPw4Ko050NljfpNDk
9vcHEQ4keDLOAbCnkbPepyYnTFVKVB/OZffMqYfcETMFTjR+XxI/f4UxYg4PFUwW2aC158tp/isw
57SMhfCos1JaFb2jui4m0bE8qjdPH7/5y4cmRfdvRjDuaKjVXytkjHKlRS8FJCbYcy6LKjyLBTJK
f5YCYoO3hFJh6pzNQV4Kjx0tlxFZlS74N+lShmnxwvVrn+StXpuBROL9tJshwSLdXzdgCOBwh9Jl
PkiZgl9KyFLnlAcMKjt3ci8NaOLNL1QFS2vILpgkGQrcXJRF92jHu73aO7Lf3Cmfix8yFOm0XkgG
mKQ6U62Qjlap8RlRfesq93N9+l5RoT2Zk+xWcnHJkXPXFv9FEp7pm54iSyr1tEw1zYX2PbUy86oK
UXVzs1W2SI6s3OkobB2abo5XTJsr6bAJbTid7h2QuzApcbkCKQyPZdrix7GaaMcAeZ6lalAaM0mR
WaHatdUUGsuD7f+VZ5ZouQlC0RqHNorh8eTKmz7ltFp4WaQhJ+JfThoc67CDqJJEAucVfC8rRo8w
JxUQa9oAqtg1H51/MunYLNVx7VjUYvsBnLzvPpi8aGVN3hxSzCjo7S8SJjFPlmN4/9W2jnqiw/4a
wEGBPNDjDuL8TfG3MKxLplnurNyBKoV4mA9DUDOSguyDr2TYby1dngjcqmdrmuM86gHMYihQ40/g
YdZolqo5Gw7uP7s1eEcpmZsank08Mt4at7hkzZkGUZ1VBEG9438XB2IlNxdYj/zsIbudPF4j4Lhm
8ymxevBzAituOn8Y+2DIPcx+Hqz9g3oMA2RQLscsl7ef9tY0Y4lLHVLBA0I7JyB8xkvaW7AgBMXq
XXpUvrCqCjGkGPG1G/O7gLogeejz4jIr6dcQLTn/pw0tkS54ldq4RH+sj5AeeIer7ixCQgagxriB
/rTStx1vMae+k6/z1mTb6RiTnQ7iJ4YomA70qZW+ZGRVs3OHVisVaVC0+NcKg3wZzVdnonbmtKwi
Bqk7xKc5CLCLk1OW3G+eERcGedCnA8dcluDvI9Dg7bu5c0c28RZNQS+xMRy6UZEK3tUZT98z0Y5i
kyeoAQH0kryojAK4uxFiOd/XAn2z9QvywnnoalB6HXASQzcreYFSMsAq8mF3Os1owihPuMcgwafq
HH+ia/V2YhN5qYdaSJsdzsoh/RFxmYH+zurr7Wlf0eMxfgNsPxy4IP8bI8VCwY/1gu2GZicRadTy
3bfi1sXGe8jgBN601nLoTBe3zDlrckZa+c7ky7C7XCaSla1Ol6TMsDfNsNlg8EutpSP6diL4AXoq
ogXEO0ziPjNWQiUKXOUDQP5gUh+C6/bg1Ltet6twDBcEz971OqF9PPZoWbS0oSfYMs0dbnE2WTla
a+VIdHOimp3zwZKBjfTDNt2ga4H8h4sXR8Sn09pxkx4Z7VSrM5AqJnKAy/U7TfG/zIzA1fqHw+8N
i1DcD7oBoqBZ1y3df4rJwKTOR+YayYaJADU6UqUP6BNBPJFn9uaEY50BqR/ik//rKQ7dMxXZ8PN1
+YOQvIJUlq6KR1ZDKqlS4OM0QcrQPUW5/w09d5trwMSPyDcKYdwdGeNAH2O8/bSKvaL9wEZmec0d
a1VG+oVnLoKH9qsVFd6+VTWng4kCkOmCF/m8/pK9dBxHVLifNF1yvooQ4MAFQa2UbS6qme/DFVrv
KInEz2YyhgW8qZcXJIzZaK/O4h/z4d2/8YFqzsluMMX39BbZ1guqarV/jo8xrYIgrhsj/lzXdMYQ
/wjsAiObJwAHCDqdY+j072U3BtA7aqSJ3PnRIWrvT8/ZgSJ0mWwiMpkTvJDYOQRE5L1tg/dVyzqx
AFVTGV7tf6u5O1IOiRVvsEHBgpZwzl/VYSVLzhnKZRyhtExIvt5iz95U4jFhPG/DI+N/ZEX0EFzL
PFnkRmyVAzirmGbPy2fFsE4TDZXXnoZxLMDlQXKgOKvKLdahBu6UEJJO7obt10uZLdF0vTSYEc95
8EqHy/scE28H+9C/TFkk52oiuztaQYl909GxZHnaKK4c6a1+ZFBlkAVDCPA+wuEkJw25zA5l8n0x
jMPgarkx7Cazl2/Rs06obomqFqePDm5OhSlXV4tZZBwscjPDA2O9cbWgNR6Y/vTbrFV4+LOeogA2
BDbpwCEzbSd/OZ/bUCT33ZiScrTGe9nNbRL1Zp0079s6My7iG8Nm6Q+KyRUPrR8IoCUafjNp93bY
kytAAYULKfKKMcsrym8cBcSTOW7Gs6OILHNXmaD5m3elgtgqnF2PmQXss6iG+7GbElpLTVWFyRWx
OCqtziinjsGKl5Fojbz9mViXjBbWA9EMdlxWWyVXm6ryxxcp5RFc7UWfcMe9JQtUt2W6dfVeESLV
y0MUm/FtpoYcvK5BByWXfHazfxBv6tfygA0kJeCCVhFlOT9ZRiHNyUEiBhCIylmmCKbyhs7xDXGo
jAmuF/KiSMyDQVZEb7WzqWX04UQKUz2x5tjj0Dd2M9MGGFFWx4m9jMZV4dJWR+GgoPbjI1GzNuDM
4xMNVu8+l+BiIqpxE+sNOJIsH8Q+CDg6cBYOBEinZAG5N/DXvsmc8dBljv3ibTxXpT/QmTrIyjTH
CaXdUTFha6S7XjVUjEQbCMWYzoxPJpyD1bsyrs/lm3fDtTXleAgVPDqvad7FdmoUkG/ukraq1gT2
RDS6yq7JfNKZQFVgvE25KHSbbbRzMXxufKOe1JbbrSEPU+6keLXSYv/Mqjerj85JfuoWPRatQKej
DMD4xywEGaXVh77hhz5XZtCo01K4vYexaLOlMETs6KTtQWGnYoZk3vaL8Pe9f4AGuqj+40NqEorr
1UJjKkap2XW4r5d2n62SA2Ya3J2J7jXF4WOYU2TSiqY4ggQfP3sGiyHWiZpkpR5YA/A7MTWEME8K
rAEt3SSaqIxfXbqLS9rVw48LouP6uNZO9IqZsI2TMKcD7VZFTuLgdt9BVZQgkGxAFqNmI77UJZ9u
xwA++2uz6J1MLeiecy3ujhQSnwceOAi4sMGvAFI6LrfdiignUfzLFUbxtaQZueJz54kQwjPsDT5N
xpQ8GkjL8hJ2kJg+SBJhntfezHtzCnZZ+PPHDCoxV4YZt+RAlv8clgsnIA8FuyAZyxEVoIiXoJcz
P6M/dZG0CUyQutvg+wFe8NCJv/6wfaIiFtHxSeI2gVnhMlyaTMNCVWFpE/OI5hpBZwcjdni/R10Z
Xkr4608tsSpFjDuypytF8BV8DSJqdOOrIy5s0TU0ZIg0m1u4HjgOpmQT6nevJnnwmbzHeolM+3Zx
icbrPCiVUvyKHFGl5qr8e0qI/p4FltVTgt5DvKvHbTRieUfX7+qhSRFZhFSS4wvkPVEbEIJFt8N/
xiF5hWoNUPCNZabV2EWo1xIi/9ABTeK591PfN20KdKF/ZBDr3J9VcemRp88f2UL6cdgZICRFvffT
pmRFOjjn1Q+a8PVu7Ckli2N+6BLNERPZ4+nYb8vObyu2AjgBSg5HaUMi2miZKRhRpzPZDkfY+AEB
fd2AiX9FF9+NXTYs64O2gW5K+Ax+jp+gCuWfaJ2KT2LE6+TLzPn9duHUJalF+icX0fyLC/mNN6xw
mtlMP/ylPsE9O7NmJ96sMUpnXVOEWlbW9pNL/rW47w30eZBNmW9QEQKdnbfX6OVisKNAeobXbmBy
xfbIisJaHtvLU7l2X51HMY3W7+L16+PJXKYoVJC9Atoo0cAT+xd3FYh4ovsWm3n5Hw/UfxCqrwcn
IV4ZbU11+OOqjwvfha+zombHOQJw56mhuN0ccroQaTzaqu+publFI6JBp40gcGb0ISkSBr7QB3wZ
rbSF4Ri5xhQeOS35CQV70Q5WdaGAVOOMsAb/4QUgoAY7ZXMdmInr/lbOY9b3o5JgUkQCKJSHJnmg
mzYXrCod3rQNI8ebCezkZRshM4/nGaQOWjzGRRISg+i53Tq+NGpOu5tE/HrdQPSgm+jTToWqPxaC
5t00tWcGIdjzJOzgL9lkgBN+752q5+IHYWMjCm9Qc0J4aXBsUdXs7KHLDf73aV9LN+kVVcmFnqvf
Dy1mjyC0diNpfphY9409q7xZubeKMbup9ofLpJgBWNCdBNjoAiR02g2/pxF7MtywJYnASLNlBO9w
QUd0DGW3hET5aCkCnKuYCgzS7P6i6ZNBYuOnW6F2JwVQnxPfbBEiQGZFyn+voPC9P6TtvhsX5zDd
+1rasilD9JkuYOO20P94mHfcjh9R6mNe0RVV0X8DTajxGTy7Z88BS8xlwZ7Mz/3+b5o6dGNdXVDJ
SFL6XauBmUJmgpu1JMbpEfoUiHEPCuRyAbTUzRzx7H17AJNBXXrtlRsxPTwxEjOVzN45D94M0dbT
A2x1jBzcfazWE/YOkm1MCgCdptweIE4JLUCdYoLN8JUhbqe/RN+wZTZhnMJVGqBXPbal5Dgbmukf
kyx619jrxR8uwAlqAJPortSjsiq4vHlFk8R4mvTi6rX0eNW+pXh96G/8kua35AQ2lI6ZPtME5vaD
dqPrEPKS1Q4caaMuqXUnHVicUXasgmRp7tksmfoZMk7HcYzR/py39fLH0w8fO5oF5H3Hnd8wABSS
7pSILJov35aQDeAfJH+RB7WGxk82JaZpnU7U5CaADJ5TlkZO4RtTHAV541UN4Q9c2h1ldJDx9N38
YHNzw4mY9QAtO3XsyMCnVcrBCyEPBkY1e2kBvbcxZ/oLkhNyiiB7f5FvY8ilXBH0Ih1/BMWVyEnn
iqkWCz6r0MRC8Sxem2b7YoiQ3fwbY5WKqfGXauzOR1AlBO1DHqA6ZKV3wL81czmSVSija93tlACb
5+ZCGeFJvqhxQmtku/AkQurOJhP1mcwLvCJNVQlxMmqF7p6bMTA/wLzmCMpS0TP5488F3ZqA28Xl
TWVN1WU6XfS310/K500cI0p/xIXA4BW1zF4YpRkhLcJfiNPSB01ZOQnQF8/jlsIvD5Rj6wh9KuSj
4wN73sxYEXVP+LvADISZHSTsKThYaaBSiBjeih2dBPb8wsP0o2ZNBmUYWHr2+jgfXHVERn6panaB
zXY+LnoMk+ykPwwenzn9uEfMP/tLq386Svlt9Kc1KC2hFO9v+ZOnedfYZnk42LJHPXjwodAmdztB
/PTOFE2aYkVOfzdddHtVIGNUuKrYuqScu3I76L7JyLTeLsvC+vwp7Yhk6EDrs5YWaL8W5DLwdVoy
ZqO2ndeJXsvrLJqGax2A6HULmG2FG+yvdc0SLVu/3ZpdyHw42L5WPsPpUxsZu9Gx4xe3L/8UolQV
SKLrJlKlRsz0FE0mf0rj/an6kcYyFK9DpCHIGR/UYAiq1fCGNBN0PcCOMHLXcLJrWgsLi+dUb668
vJSRj+1+TxMXTB8R36NxoCdLPCydwzJtoVpj49pz9YIlYRvSEJjsF8duUTZ+jpeIeHZ/f5XtjO55
gAZx5Yp/rpQUZneA8nJsFAl0GAyLgFr4WoM7PCgjbJzHo9F9BhUogSIVBQ/APOXy+MniNVvJ0g33
zVGtcupU1xQeVwxKddmmyleuKlLG+Ey9CFmg28REM5v+WrXRFTfkJr4ztFMQh4+G+RpdVIJJ2CM2
qJkDFUX497BidMfWmnWGJI/Df0/uP6IHuZIJ3k3tnCZitgALBy0igBj1y7sgsyBOe+Pv1d/Ai3/H
07HJoEkYDSkuE3POtyWAvPpE7h71dX1cmP1qZR0+fjXY0C0+5WEikg9t/PHgBxHNSfGijJzm8j/y
O284hhNZg5gqeKZNbRxOOzySHwmxJX2CBkkdn+EOeTkw+UoKs7BY6r/Wb/SNE/6jyfS1VugN87Fv
Qrh9v/dR/zHc+XkmyCWdb0umPxk7gOo9pD2sjV9tbsUcqPGxlVJ+55J9fNidNZbYPUbtHYFlKBAC
0f+uCwJgnVrUVvysqhX7P8sQq4G8LUHfmI39tA8Kdgb9kni5Rc4YPYCdr2MFlutXOvuvuJFN7bMK
70C3IxARwMrYqGyKuVnbQuAE9UIbbZ9ECfcZryJFhLNYnAXv4EHYhfWXeQpl79u/eQWP4n56K6+u
ETJ0GA652VlS2Z4xwntb6lbQl7SQ5OI9WVJceaxRQMRO5635cnDFvYx5OcA+bdRwFXExK1q0uJxp
KKas7NWXsheN9PBmtXmcFmqcu8zBnFNlOVWvrlhYuvazSyPC1D/oXZ1f2+MINHNWjqysE3R3MWrc
w/QXFSsg4AnlyTI7j8RqkxPcR+ivpD+S0Bf+UmeD3tdrI2C/8JTWk1/ZhEZgAeu7RYPR4mllBTSi
elshLMvXO9PXQ/gK2vynrjQr+5VUQ2hgausp3dlODYicR7MFAD1VUc9+Eboa88/BOc8ApbfNEIoF
wqvrAL799t+wrsvsl3LSnaOuiE0O+gXfPhyxbvQHPrugFzb+KW0VrgnMsB5Fr7u/grqavgTFs1jq
GByJ/b6BSj5OpQVRnFXIzAv074mRMA6/xO8dJlM8PHX3AlBiMP4x3T3W4vrJjY1FHQjsYIva/yFd
NBa3Rd8Db4Xiegr4oRxtQo8l1jS5p/jv3sH9i1emtowpkfMOJhVuO6ZZgOthKxdtyjRN7z8AIIuy
BdkkvEzoFANNxQT+7qRZjEgkWPxSVCjdU3j9VE+UAG+W/biZV+fxka3wBymWV+96vPqLahE7f4Ww
Pap6A7TJMYg+c/+WZVRmjP7BgCnp+b3GaZWi39INfNFC5S+u6pu4IHdmW++Q5yLhpGf0bcVnKxQF
wijjJaD7Au1mO30KwII0sFm172MtSJIKOWwi+NmU0gWy9IdDalrFbIytssjismoYjCiaRxvaUoAU
aykIaCHHdJ2EQpw8bmRPfhGvZSh56Bh9bosJoAPJX+DIxzRcO4pLBvB5L80jnrPolkIEDKsTaZzZ
NsiKGuQ1dI7hQqyu5F2otKzBp65JugrnHpxqSHDE+BzbSuYop6O9vPykGkFRHUT4IxIs3WRddT0h
cMC3ytaXIG8a6pqEB6jDGHu9DszZfuP0MgK7V/xMYVjr1SRYF//h8Rsz8AKXSiYO71HveYYP3md6
PJ1PM/cFhUTx00paP3IlPiyjiQGtANqa/EQfTm6UxHO3lwMBTKHDYH6tI3eQkQ2jcFmpwJw7a1H5
v9gxA+0fSY2lTPnwgDzHT3gspIDbBcr3ISF3ja4lRiY3xChgaloITCVaTCrzNQK5Y2hD5QtAu6VG
mGWwvpt6fuQIXjyIRcbKP+PmMf0TusqH/WbBOQ35El3d+69cED9egk3H+mBOX5cbqmhzjfiNO1ef
kdmutg8sOrh+BOkqH6hkAAY0JyAWVwAlKReqMvIYOz2Xc69rhA8V97vriL3UbCB0FoafvUa806sU
L8+IosbvSNp5tLV3Gt9hOZT6hpdGFWAtqc7HIa1Ec1Op2s1VP7qSxY8Cjv+H3LXJMvNmDOxZcghu
stoOHnluITKjIYV5r1DeVBiqAhwukX5Z/ePbdQLEMYw4J4WZgCOcmTpKTCBsRyTAZyQEgejrJK8h
AEiKZYOdp4izzMoH0pkH87fuxhtzrDHaRV9zKCl6i5tZ29mrozZ8SAjWE9VAOY7wWpC2nWbVTxsO
aCR7CjrRV3VwKTTTxM+UDanTSDX0w1dTj39BfpjDNrycH1h5eKThKZqQlxq5rrBr+ncgTrngkt2m
SIUuYGS0+/4ss6UJP9TK2DE3uk3p1Iscm2BGVGmQUjquGmGqewOUENUtdI7mLLsi2VJqxiUWNg8D
WJcoPspu77p3UhERR0dZpDrgMkRdI2vUQwCvq6X32JH+NTQRFF9sLUgvd/O4fdJ9mLBxLU64uBdo
ST5j3gQT6jPNzgvMmF8UkNdH/MHphL4UdFPesNw9Vkt4z1PUo65lUvU7rC3nHzS8Ayej8WwHt8s6
4GgNh55ol72bpiwFnGzc9eKfRZnD0CBivEIwavoxHI70Dqeu8rAv5nWVhA/Uobs9mnct07ZYHYG0
UqH3P3iuwqL63H0JT8RLyQquSCjUSBl4KR7TJF8cVR8ElbZ78FMnWpqQfZ7rZrOf5g9pBi36ZScy
qC0ZxUemn240E2LPb4JnvTvagSjGFeoqWfXor+6shwF8MOH1BEgknsmAd2hhQzn9rk6s0GB55tkl
jxDfFjg5hg6I7wzJsI70abfjSVj4eKGObR7CH8r/JcJvu8b86xwWLnjVYEBxnNTxuVBpyOuhjndF
l89XJursnmOlhf4aMjGRCdKTeMJpgaykNbnytOpVqgSFZ0e7+/h/av4eRYxmiWTbn59m605IfZgz
JkZLvKY86NN4Argvo6yIXk0vLdty6pX9m0tqlI7ycteK7k477Xel6PT64DpsSOc2M5fTWWk7el+i
TfkEfPZYJBjQ68WktN1ss7k3Gyfrq+fbDlHGSg3rTMapiL0i/vUQCfzQ7dwVLMo5rLMAxQJddJyl
0nzkMWtIePAnlYJQqKLCIAPjg9jn5cOk+PXdUoqFDL6rXKOwAti3y7dtPiN5l3N8Jqi3BUBuk1Jv
5Aqf1bq6Z6B+Ftm/m0I6Bd/GUylCx0LtEspYsiKFYBKsrn32dDc8wEwvREcmj56QruiQSnHS43bQ
FI/K8YGAY5uNC63B6p8saAVU1/xGtUSiCvKu0bHEPj73z5QnlvyZyqenY8AYlQE9GR2qnKUCL00t
cw7RJ0CtOjTzkcF3Hw0gchdur5TRNiRkuHqHfcA/IX0NpFpMS8Wf/vzvk+kEtMWqoKedO8+qU1hi
ZvjFqqNVlxajzxnjSPWW21yQ/Hw8SNAbVdeqQA8mFXmpyudtBdHwbUVSuoN2P+fr8+VLy9TnG0HO
SVBwpGh2+qx6aV/H8UqD48ckgsZh3LPGOqCJYX9ERBWA+h97WSaIIbDjgExvCS/L4bdOOf9bKuBn
0eblKPc3ohCWmcQw2Yor64HKojGC8HEMCEOOrw8ny2sz0Fg9K/aUHBVndsH1hSI/K2cAcLwdSKKA
USAeJpNVwMbAy3xLnD3+eT6Lm860Wndl7TZHHzLFa4RCuxbPVZ8vSuErChCy4JBTki3LXtWaWbHP
yh+fDcNIpfU/6hzo1jUY4+ifTKaHQj1NQX5ZXOlXWNcgJQACcio4tClNHq0axJ1VIIeC4qXYYdMX
q61Qn2I69xJcYU4qS7+t/LaPzoFPlbG06LX9t8gNQuvV4LwNjWcdIzDvstCV6Y9LG/Ii+VWEEWoK
D30L6SBSWUdW9xzT2bL1M7XlWqtIIUR81BbvShMeJeOGg5hUzrdyw2XJBpOLzZytSgAH5+uhM6B2
e4Yi/3NQSgwpGDfQwm+9rv6bznn9ZLdylLW4CCFSyua0nbNO/uM8InzCn+Lv+g8gofEn8PFn6pPk
ibnX/enQpnSa0Ur0Zpb6n5FlPvGh1QT/jLy2rHFEsPLqZ0+WtKuPoH0LG6asTCM+Ocaeeg5AZld/
U+m8Qlst/20wWkT/iHRLuDbXcOgTZaf4qz23Tb4aDTGW+w3Nnmtdc+TCTbrn/9hKKT1m9ZyEIefV
0HTlmEiqgejB4OpSVxZ+RdQom5ruzk0tWyCy2JATpBpgZjcmPSPf6v7zQXKXV0/cuc0IPeyaOswp
e/hfFVtL9QFkqyg/O3HnlqL8zMStuxuaVPxDmbfcIkNyg+n+bJcGostqATi9bv/Nc8yDw312Yi3E
TMp0DSIiVDFEiHhnpyKldsvYmk5qbqL3QSBReFGmC5zgGskxDmXa/XiZzy2fhSS/0EqiLl1k0X8c
XApCdXbJWMO0uUfa6r2Cr+IMOpmQgveXOPy1NCbrb0bXlmMAyw5E8Xsg53e6gPi6yZ7LnNkhHTiR
3FAJQlvlvpVWcMIrrNbQXCXCFnZgJZYqwhnnXWp8mR+yxcnQySHF4Emj/gS4DHVXZTbdlaKc/aSL
wyl0hB8JtNsRthl+IEBTeOvk/ZC7ay/7O2uFqVZdaOvaUPn4knX7o1K5uR8uSX/Gqy77+SeZzAka
wi0jgZeF10PCb3RI1Pjz+AVDAz3xy4JOjqYopy8HNboBk/KG+cWQoLUm1wzNM64mdwc+a8yVgmtR
8w6gX/UExE1Svnbg6QC5sCN7S9xIxLCnMQU/n6QvUJHPFDkdrS+a2Gbt5Owv7U6N0kvw6R2v+Z1F
L3DJAC8d8mmTPTbqOMbE4TJBCW2XO1CC924/pmC1SzSppOPliYiBtA7X8MySujkNc2IfkEg04Pfz
Ibv+q4bgukFmiLg1Up5fh7evNgJzO1HLPw6/EQKXUvQAVWgjRb1kH+H2QDjjKKkcoKVh4HjAoH0W
JF90//J/iOM0KKoPwtlIAY7UKjGS1z2UHBKk0usDiSkFIxeCvsb1a5nsNjnDvRx5DE8CD4gWo2w9
r91JhscDyyQm7/sZ1I9oKO4Ny5mPW+S/WHqx2LFqDI/D/McaVKd3hwbB5bRX1QhgdP08v/CQR7m/
DZapWan4uJiWOTumBt8cVJcJTi3Q916f8WPRHY3E9q8zMSJohbYonbiW7lSIZvAxssnBK10ScOUx
GlR+LWs2Dx8dYqxwZMN93Bm9Zw/YUd8nFzasu+rSkwbUJ8iv9i/a4ZWdYMjZx2hpv6SIFEI2+t8+
Aa0IqI9CFxOEV09emALq1S2wwElCo10NBex5jHthwsfidzLC9EiTcPu1tXePxL1OwTV3eLlqimIt
clZG0hq8W0xNJjI9LuvQIVSvI4rdqTDlLam+J4j5aIDXoPg4AXLuXCmKD3kaigDE2GLSwh0CvwkC
Iklf4Lih7N0VloKq7NUlWKAhH9vwyafOY3KWovbnNxIsM+o5yTcjKLBx6bKKf4977Oan2JZNwBxe
oiCJMVOKJwfM0OHG6eISanYolGiViJ5f0eytJupgPA6PV6qFbFpKmWLR3sDSvHYX/LEUUGzAcoV6
w+PJmKBeDhGlwtQkLVWd6mO9xcgYfFGRcMWrgTinQ1uQMgMvdplBkLSFSxOeB4GKHot4rQ2+A0QI
rdVY0Hk6M/nGDtWvQGK7mrKk05bFi5zP/ZlwzB+zuvi/Y/4m6boERbRGlibZiNKs7dtjMRGeE45R
mFQgeqkJ50ZmxX/JjyRTZnnSHwN7ud3tQTXgsddkbIR0WkaF3UIHweXNQooKZEEYq+JQ+4K6kcCP
PM4bNK2e+cNgD0oo0awrgS6qoAHoQKMCY5AOY2tE3antdV32Xa4VBj/wPCYoQV7Aem28jOKr94cv
g3HhecCZpbXeJf8KkG8VELq0wQB2kgMuoN7vWOnB/merz5U92Css5y7NrXsOzcgENn5irFbCjJ/l
bB166ZBiPR+qYlLg8abcranIioBN0sP6ddVG2VgeAKwHYPOvPprH45ValQGeE5bzi4EgBR1BPAju
uHZnuzMrgvk2L3TXQ+uwDyoEusAfT2qXYJpScj54WjMpYBoHiwNvCaVGyvPdkMOQ+gWQ9b4ekTHP
kTnkOiu5qaQAnBtSDEiSvRO3KPxt5MTYPUdwkggc9fkOgqRbJZV9RLGDGgR4x4LwY4d5qbAWz2GU
K3LcDk4XUdsZbjDBswUj6Vs2zJYxkfd+s4llQ3HqBc0JqErZnQpbOU7qfJFk4DkgtBf1OjN6vx3v
pjV8YXoYGtFOND6918+FOZPmLVU4wHeASLM7fBnfbwp53u4GC7bDriEctjG3XJbpx1y3bo2Dp4ho
GqwSKxzgaGZnIk2NiWCTP/Km4dt6tLpeVqHF7ppkgXKU5IjsxphVdLsycHtdsW55t4LKqp0NcrxY
Kl+fCNZ6z2XJGEYy0kiVEMkh/6UuNZZfO9I4XBMzZML2m8XyMt4vG69Y5krkWKRtaGdbSTsXYrSw
2JszYxnapFgppoceaqjrPNt9PggAasc40m8PkOfQOojIzeUDkC9M3LDkTFdMqHUh0f0Qk/KOdSyQ
1LHp2O1AJbz/HgQjeDMknn5gUhNHRWhRBJ6UsIebFUE6D0L0qPM8BzBjOxhiAHQ734klVPfX+USe
GFw/fkAOyOljxg8hlEE+yut644cprmR4EhVsTvKtfIa5DNfc4RSCSFknEIdggdJ7oAQ29f0olhlV
TMSZdOfvg7thnIjcMubYaRZMF7c91AG/sXw+t+8Gc8ARoTaItfHgmsfwEJW1nolYKBg14+zOaWKz
9MxSkEM+YVhA4ez6Wau+z8iWJztw7OrzQmjPDeBxcWkhUeCSw40H/OEXgvrAOWYZsSquRYefjPV2
op5aYNSUz+oQjS6dKtpSmTy0d1aJeIGWkmFBSLTKmYP3gziwQcZ8mhi3G8xLX0xHGWz2v+E5B7ip
bzVSEuUeH7K/0Xlo2tlnyYnwsX1tz9KIJgKEriUuQDQm5p+5il2OMW5r30CmJEbwt1RPIFm8yasp
x8N1J5/hF4Bn7KfxiySJ4jz37ZI2mGYAWtlW8dpj5lXF5AR32ilTLlCQilfu8QPXAViGEjXaT3zq
Gty6J7+GfTU1tZpj1oXJ/BDGGwpHIHqzNBPYCZGkmQYi7wjnu07yoDboDhLYvxmUOHexIyvhwKuO
NN6J+QUqdaQKqiYrLVuZET8sUHo1XTxnPqwgZlsukPA6ztQKDGFKCCQE9ZHV2q/0hiQKqMbyGzyv
vCoWCMZ9Ent+wIrZ1UIN0ErFTZImlGFVyZ3xLi8c3dI/HiCW+1ZH6nVEz+3K/VQLxDE+gixODAJt
fute95TQWfyiCkNUpT32iOuqY8Ix3K37tYB74/eF/6BJy7tb5MSnn9YBrQINaHAN/Z4gFi+/+pSR
v+CGvfmauGkVcwEVc2zTs31lWd0gV4B6Gb4ABKCmytXRbF9QoWGt11qSWVJdx9u+XTM6bvzelkwx
0J2kP0F6fYMB78lv6FarIpWvGvcrJ6/Ro+makmk4RWKk1br4/dB0QwurKVjGl/JRzPW65ZYdDeye
TcYjMiQT+sCqt06SekbyaRXvUI4GwTrGvUTA6ZSyT38HrImxmX8yc//wHbg47AnlW8yBbL+JTOQ2
BuQCcj5Mkds97HbxjSewuZdh8D5e4x9AgSjCFs1wR242f37iQBfFXYh0OBapqow71MHbvZmKrBpj
Z6LReVzcj1KqXTGoFFBMY9JA/8NV4GepTvBEkb+8kyuHkx1rFgq0WPiu/Ey7W27o0PBAkeAzp4oy
LUv+wEGsG6NBHtFUOrCN4cuI3Kr0Q5ohD/J7mPTLGjZAAvN5cYZ11KJGHdWJxBCy/yWhVytviXLb
DM0ffawrMPIyFGwR0t3DjnDFtWwN6JFzvjoyGxs5E/LqksIeXxOTXDg3IQG/57zp/HM2LFMRFPeZ
T78glc2K0HqqF76w5LdLhj83q51O94TOiy4oqYpcYpXut8eX1Fs42QNECw0f0tF2ceMVs/Sq5wog
pkreXUy4Vwdd07hK4LGHAfXKJj2Qt2OmHqWj28VHbQ8HO5GDxgh0dy/o4MvKW5vV6mxbj7os37wd
LwnTRuR1nxKT9J+b7meK1yTER/SNB8YaWkl5ibl5UYODlEjHQftT8bDQ1fx+4JfZGNJHCbrkS93l
rJ4bgtLHd4xz0mKRcqVWJNpwC3QxFTRTLHymMl+XmYQhW3cBUf9TfEwx9NbEFhlBz5/rEkzO82zD
D8B7XOm+oyN6s2hETTW0p+5wkNFpcpUYFTa8HHGdiRthbSkWuA/XGRGTNXv68iPSG7l6aZz2K8IG
LiXf2IR4OQ5bunSMh213axk50WVc7yCMid8oWcfnGYaWwgegL8qGRwSDBRAXj3RbS8gwYKeecDoN
nZtVI5LjWik/0QLWye9+1Y2DQrxPPQtvGS5Og2NUljvg+BQ00xmNArw7xjTGoulupi83rpRBRule
+0DyMtY8PN28/8UHctfgxMz3skov3j6pwjwke0G21LIZcO2pYzsRkYK4ojI+yeaJWjiPFtcGgqNd
j8v5rMC+XZWqI9Oc7IQnSiy+E/Phq8Gqdt6DWhAdk5ypzBbzN64DBoMErJIdKyxhHO+mP9WMIYds
96i28wzSo/+EjopUTokbq2VKG+zvwAZ3VeBsBCSx/8gml2tP5s1N0BH/ZOyjwbKuAF0XpPhrzkaH
RiRy7CL0dHhlzghI1bztQQhNqnpeSYoALLlKi6oXbSpBrm4enPSyLwt2v95WzWJH/PSk/XY9yzrw
dnpC+qFpEmia7oGUsdnSkLcjZPVgjz6JyjTCdEUw99aGkgikRyD0LvMVf+1OXJ8D17u42amvHA0w
vVZhQ0EgLhOtkVgZ9ygM0GflRR3OUCoY4AuRD8NNVOhJt6Ew2PMRp0KYP4MkC3A/lYKydZRUydEj
jTP/gR6b1GdcJPrLmpq/5bt/690R1SjuN5n4sYEAufLkePCJc1gm04ILAQbWu9mZcrtrYvsWRwHz
sCVcGI/PbiJk1JXeKg9F12Ku72h/K7r3hhNqkyw+unlDFVu1GVsEU+bqcaDJxpFBataFUUOBAed8
GHIPD6SBmR81wgCNaye8OiYYZpV8wrj6vLCfqSTs3ZGR6a8FvJMYUUnuUfBfaFIbCS0aU5/Vzzn9
F4teFX00j3d8PBD0zDfkF3atFFEDlwrO+8+5y4mplw1bNVg99atONmipM5RLE8B8uQqV2nj85X3J
ukOxfkd52yt/48zSdsiNflJvadMNxtxBTVmvpH3KbvugDoObw8iwLh6/CsY6LMsl+ENXqIyRjEQA
F2sYvl9YMNEs9FcM/DS8/0Bh2WT+OVZK96o9nYTFT2wv7J3I2waQ8tjFbBoYOKQh577N51k/10RA
a51NMVEmZWxbA76x63AvYFDua9W4UHkKmzK5hLO/CCyK5WLmbpSIkCsaPw8j6slmWmIae0/OPvyM
lcn5hb2JTQk9sUL9d5LTH6kIqSEVEvfqVKXVAJB7ntCEEcsvnE55ItwwvtG29VBfpa1Osm8QyM2a
9SmSiAEDrHRxt9dwwetxE5joRVSBLXS3OgVmnn+FAPghuK2aNJKN6qOofAazqVupHwREZKtuavMm
0dPgJnG9wXls6NUH5oOWBGSxMb1x3Mb2ernSM49NojvQd7T+Y/HMP8v2nwLdtM40k5TxbRM4ZncL
+k/oMzHxfdY5AEyXXXixqzFIZB/Sx9DLTxfjM+idWfxo0C2aSFjKYNhtWHMLjxbXqrc8P/IFIGbV
Yh6o17SQMrWGtEoW68hkPu0xGyy/GMfWh0zK/TJCsgp76DYt5U+8cueyxbAAn8jcfpGhkvlDg8dk
d3Zi3n6knfwFJ+3Hi+jtx1H8t8qOF0vBeNnDx0Wh34H54NzsTk3CwOUF0nnOjVXd3xhHToAlyN8I
HaJHnwVbrRjsvkxy21zq653djqukCr+hbKBVBOP2yFeZywWjmlNBhWE8gKI5IKs7AMxpzIcC8Fhd
HaZ48uS0QTdLXND2r5t3WKRM2xkmuLnnteMwKa9rLgCbO/6WdlJrhRwqq0Dl4PDINQAJsuMuohna
2lcG9QBrpRfWL5ZpjnDVnjX/GfvK9X9UBGN+3ENq6ZDWX2rKlVuaAst6k68VTNk86MwXbFGWsmNR
GNrbQpJsrwOYA5VE3LQ7z0f4PhL3wXaUHXDGkuug547y77VVWQHd8a+PDVgd1rNOpzM/GFJ+svZo
Wf1UHzQq19j+gT/4Mfm1LXtdwLPQzwpDgkcBj5ENOUNXWXk7B5kS2QKNsciATEtrhnd/Fzi5ILM7
9kRe2yERkeRfd33+WrW81/xNIRs/xRxVGNZd2k9XXXHBaAetb1ntpooZDL7KZ8FN666jfST/tnEi
WZezGzOJn6a8u473XVdeTnJZnDAow+uOIp/wgZgyXZ87hHhdu7mn0prtCAXezh30+tLVlGBXJryT
yqa2RkmPM0Q1g9WsLiL/ZdXDTY9mn/Qh67kP/RsGt3Feax5lrrwa+tkcKfapq6QS0iXcz2bKTsUd
hj5HbZffQZParDYRe16DN21vJCotgd8+cQipQ8My7kdNkh5lMp85h9ubv6QLi5ZidSH6bzmEs8Bn
GuKqJz2szF+WDab403GTUYTJ+501sh8EGQgiJX6DwLP/YFTmIYvKLiA6w89IYstHU+KnAHq6dSoh
e7lB7StMN77kT67t8rOlAi1rgeWmZX35y/H6dc86OTOL+cJ00vQC9PADyeBIwiPPwpgeEoFXey05
CSi0bPgtZTrteOndvYNCEBZgfE4kQ5vH4vMO13rBWyVnrfFm2wLQNlHY+oOLexbX1yx2EGPn6Oc/
3x7AIoYxcBQZAbX7tKrQm1qyf0rKxSHQIr7D1ddgEEkrQDN/zzK6JoKX0IEkJQxw7jsht0tPdewx
PneCZ1LZgWTDaEIHbYhYdSByoWI57nUkt8POImfdR0boUMo2tFk3rVMGLdsgNbJlrH6yKQ6UPNtr
aqR4MMZ3R7Ua5T3LGKev0uY5NAv4uOZJH48nCl6F+BfTdZMXGCHRm0itzSnFXPSYCH1tHPkF0kQc
TNHOnJY586CjfnPGc+d1JsqsHq4iCO+CsbHeQKZaDTb2m7SQwJs802C55xOOrknM9Z/c4ybYy5xr
lEaO1r8LKTfQqDlone3NndLEYnVZtK3IuwMVofl7R0GAi6ogWAcT4oWsNV/KiFlL79MCK7c9wgh5
iXnO6VkYMp78NMP0gF/MiEH/CEedTgwraR85lILZIdr4YU44YvoTqYINPKv+9Any6NMeiy7dLqzU
1Sb4t+IazYnGQ8f3D4EU9NTVRKSwx57r66k4dzYga69u312zYLCCnZBZjB3FbU4/7EsKFTfFxvf5
lDM7bczNCT1knIM7zXu90rCO9k//i1mv7Rs+hluDdm5tPvRikLwco7Kfy3oHbP+DRyrWGOVmOEsC
UuOcyuYlM4t4z2y9kkWTEvYs7iMoHwX/uLOoIZUnWRUj2MkjOpnzmIUOP8BSYAb3v5qvwbdu/MSw
oVngTZoJG/u/z6+3syrSnmxm2m1rkxAfCv9tWFijKCs3VZtZdjkX14Sf39hHbwiYYfSofA44F3OF
py6tfFrQeK+Gq6qM1La565xQiG/jWAONNJ8eeOle2AgOl6Run5k9WqS9v4qT+9Fw55SKPjC+9XOs
a+/MCeRGy1GAHp9tYYABuKI9ZQxkM1Ntfj0sm6pGZ0/EXlOVsldf0SfczYSNnj8ei+4XTLUhEB0I
UriRUxbsk4L6IB/501iVSEg/A/9qUHPI2IJtflu4Wg8OXpQq0ZX+MegDqybXqc62vt7lAukWtXVh
zFs2tBl6nmmOs4WnMKU4qNIQ3Dk7ep7be4Cpe0DC+eTahl0J5t/GqqRWGlLEe60sUFuZJadIUpQ5
IASo6S61B4IpEKljIqA28rbj3oXC1tD/MloIx5Pe4iL7vTi84RDsEmuR/vcCAHRgxCGrgnDsFr2a
oqVgMnpLDjfmWAZw823zFbhtecbG8NhdpaY7+QECB0ztswC3JyI1deqSRYksk18uK697sAEzTZPb
NT3LO/3DyN4j7yPj+17Fxm2WSuW+mFgJKIsGCsujgmwEcbRVTFmQQGIi4g7h7vHRWQFKM/dRZaBu
Nsdr6V4ZOuUMrGj7lqQ0jS+Rm95wV7htg2Df1kC7Tqulb7v8Ny3ufEBaM/qCGPOh6lOXYa2g9+l5
qGXlEN7OgxGivLb7cBU1X6ifFEOud+pWh0I4g5w22C7ePkO4dBTNH3IagJ/1EYmM0uNZNClMeLyM
SeOVov6n3auyBw0Dqhmn/3fsd+2KY7RP9YNkablfkmU7s52TuW7DY/0L8vfjdfCVNigNT9vGQ2lB
NIO3HszSxuGPBorF/9O3F5sN8CWuhz0rKJIXB+NNCYbuWaZs0jyuJI/xmARJAHzAyYytSwu8OGte
7u1aR/GgkAO1qaiDFn1R1x9R+rjucomL4PmS2LInxy0yLgv/se4erPDBbhT7eI7WnPSB83Htmh1o
0JiqL9oqBD+dYMSKhFuOfuvecpeYINzsKP21UKo+3JE3dBPb6iZaqNB7uYQ8UHw1B1K4lsgxlPKH
3BDxsx8F8T/Yo2nkaSr3uNSBihcdDOsJtk7PZqOrCdiW+hcw+1bjP8dbg5fR2ezW6QCat1eIexkQ
7BejHFpyflEsCUQQBbUr1apC2Z9G+PKKCixSKHoqX7vaMxz2HHWjQs3JjQNCQUboeiZDYAIGSd3b
j7ua3PnisE1Ohxi2N/6T2F6wruoNIW+GQ+hZIn0mTgbEXM+Dd20mLZuK42I5VHeYWYgQQo/UWBot
jnguGuRSanDIU/kdRJba//JrXYmnVmpF4N5+hIt24tRKjL5Pnj+RdFZNIV2Cp40u8bVfLHGjJAEM
ZhuUpgmipfzA0vtR1DRtEmesdXJkW0UqKRoiy0D7l/yDwLiL2VmwvXL7EuCg4myVr8yB+usSAcwK
3uNTFRdXQAABlPPsAJLzZLH9ReJxWHKz2p2ypcrext2WqT/Uskqv/zQLn03Fe11zDhlqRSxJd3Wb
o5lAylSfcZd5nDDQkht2RIYu+3owxV3tQoBlVHfufw7QOJZiHyK+LWfPi0jATw1TPN8SqForglkf
MaDt7V3DugTuyA+7vMwpzvG2y8xfSJfUK02H5DRB1AozIT11BgBnZcJnwwFqltsgLAsccTk/7und
8QnV0Cyx0JfO26Bb+lxe5FDdQSTjzDLvZLfv6gzzQuoula5sBiS2fNaUTtnfEYehz0OWZFk+AYsH
9TvdaBdPQhfOeHz7o1pD06ZM8Ei+DXuMihlDWm+0s3/zwxBYeuYUy25ES0qmgw+SXnsBlb+zDn0+
g5lrC00Btiwp47a+UoY+WOr6uLUJ5DlKr7kPLlUXEsKMHaPiet43LmxTGad7jkBLqEPcQEFed6in
rDGbQlm57eMamkCps+Py6ysfdXxWLdNXsYTHnkYylGuOUwrTVz2kkv3zWJuHPdx3FPuNieIDGt00
bL0iMF9i1uvUBLOCyRCCXosGqEuHupmDfycfRxYMoWKbNiCzKKQ5CPbC8gm4TxqhCghQ6Z10i429
AIyvM0SHeHNnS0hG4kYEjLy4puu4hmq4/LThP0MECOlaNz8h9Lhe9VVvc+AlcMJw9cFi0yYR9VaM
rP3Bls900AIrq9a0PUXTd4kmSiVwNnOJ/0Mn4NXRKKQhYOaAhI3Ghykjs6G4f9phBO8CsSJJnzeI
L2oKzLZ4Umdwzc3/lpB3QKhbeoY98CvRDcK4u2+PvRrUQZj4VWBBYfCxmPKezg83i4H09B8jpmXC
HLI8dOKR1zsnuNOkPTrVu8oshfgwlH7uiKK12Y9LgvpqWFNmeyH0NsQKIOTbmenX2W9BAFmMU5WW
l790ERhRsSm3aB3PMHib/XDEvolpRJlK+W8FGhJSGPchKa2n8m1DkNQm7dGZjJ8C9GgJTL0HNGcv
rxnUOAnaHmHq6XoAML1lEYbU13geZH+9fc4BjItVRxoOoAPQwHo38Ti5uVshO/iS5on5U0XADWUz
LezmuFrP5ulwiUeoEYaEe0TYQ+v1eN/QggXOamogKBiYL1aDLCKSwzNMPpfYAZniJooKJzRemSeN
FluIlSghAv3vsdQotO78N8xva2IWXk2OxwXfkgWQQM8VxwhW2U8uoBrUb3v6k4tJQdDHxRQFaiMG
9q72IdVhe6BZ9TpilZW4T4bifDoO5mjMOj3RTshsGnJHUAmv81U4JCVhf4og2yFPugsII8EjHNBp
lslk7seIASYhK7s3CnIcgaJJeVKnY0TPnXy+/jqCp5oPPpw9SVZr9bF3ecXxNGi/8uTHYNYJoINO
anMvxAsxnEwhVysWwBeBdUV8KopUXLOYslYYSGlaAvKBYamee/8lzoB3IxsTOLjc5TljC9qQrUDM
WIDfyUi4tTBFphLlPlG0+lbzz8jw0Cttg4YSETTCn7DjIOiMCjjCKoXgGTx8JJdiofmRjpZDE+oe
ZDkVMSlYCry+xTz5Hc8JKvinB96w4M8FeFWZPUIbl1Rppic9RVvBOf/royF+hzIYtE11Rz4sU5MK
CBdegX5AQH/lIVASRV/hzBxYb6zuxhD/f68Uc6R/1cnYY9VF9/Tto1ahz+Xt8VqX3MBKjndymQCe
+jbXl9Nsz4LZGwT2oFgFuWG3hzAYWLGhhpSwNq0BP6cQSvJtVA5UQOxg5Yu7d1c/Is8gRd90TjeB
ygAZhB8wKrf/bPBQ02Bi4h07k5T0XI/IRElKbs+CxceoDnnRifjGXRR2orbhRv45etOoUHvgmXGo
RQEtWwrg+7cLxRF47yk5B6yYWWC2Efv0WmdV0WHMxklbaEFSUAFehAIsvk2ICMBGKel5OsF4Cuon
16dR9t12S181QBJWo/2oCYWifuUViAK69x70nBkD78uO0jjgsWV5FxKdjfLEDGIIosR/7VQI+hLv
gN1ocdWqasYn82rLH4i9VgyYbHKbYUl+vw8tO/6Vl+ojN+vTpZdaIGmv1XscFJQUc/t0Jy+LQPuK
JbdB1naR5wAoeufV9vy4dfMkh3AawoIwZ/GYdTdkXsBn4I39cItuokwN/UHJ9FVOOyjsu2uod6B3
Y2M2Po5pUMnrBwSvS02vf19/eVPAYDCKfWY87eidOmjYLQ2VoE4hAIfgGqWTuwYe/+GskGGk0Vc7
x2SgC0PBzK3PHFaK2A2bBan59gyaV4VENmlQ718QL0D1tFy290uAMUQtnTMSbqeLJQhVp7EgdhJd
gZl0iaKXAZx2hG/eQKyAwZa8Zm5rVSmgYyYjLg+9SE/eV/laFamRDsMgvYb72UW5TX8dgSdkJKua
3QPzIL+adYoCpbdKLVfuWzRCtak8Cd5lIPkb7rut+3MOehP6k62qRFQTGCQ/L2MZcc0y/dYXI63R
FuIHgKRpbQEwMuZSfIdZ7oHRiSuk3F+J3I434YPxM3xYYoTx2ed8A6eG8qC8SAnmgEfZYExslveK
n/RECVlK6ObP8s7DuYKxsk2MeCJGNYRJZN0CJ9h08/E1I11wO88g/riTVOls6mH7ebVe3NeaX9iP
WE4qHEbiHWIfQGjBrrnZzQtWpOhDSpFPqG6vOl1V9x1L1r/lxCICpZ4d1nwehaMW75DJQDAQ7lWN
Tf+qnZXzY4nAp66/sJ9izBeptJDuCAUZrIFPMQwVC3AzUqf+kxgMb7KM4JB0L9g8dxfyUj2cX5rw
aXcryOXB+/HgoU6MrQowxoUp8JER2fRntazkJvfbviygAv77K39ldjSL95MLgdnjgNuaBqx7Ef2s
AvV2YOwAgQBzQ45bIZ2HxqGYb85nNVdnEAbjTYsI1p9U78VSMBwCVrwBMp8cryPTVkL7yjpADGcF
MgQXzpSfZta0D5Z61uufqTtW8clpw3ZLJQrMRcbyTUAKxOr8Fa8mlXeqBjY3K6UwBN/ZYCrufIVO
ecuo2Pz/WA9b8HJnP2ZeWxHfTAKKRVFqR32kwT4o2a7BkDAh7q8q+aQZwaCrLix+oqzLjY/qhrvH
ZeE8CWHnost08USqptFWMWxmsla7utY67koRWlpsWzUsxv7nc7MQ37CaIlRIfW4UpwaI5fMNhbeb
Jt1yO7OmEXrfslNsAu6Un5DYfR5kGt5ajMu8jsC0zXVAadxGRkzQbP9itpeXu92Ny97Pa5Qj2ohD
Djl6Xmj9HmUN+wjmjGooISKLMul2oY5hKtXQ2o2/BMEJGzKemEjtZw7MlI6TJfMp4GaWemkXNDXY
ygpEg3wRw1gmU7T8GX6/SQvbf84DR9qFeB7BPO2+NvXFKRt8Uf/xD6qfPg3VwG/psGhGRe6ejwM2
I8STi+tRzDXbp0jsAQDKbGA4vOzQPQCGizNklNHJLm7Gs5ZAu/r6ogwOmTIx85e/5lByjpgke7bT
nkVBnIz5GkoCImZ2JHBIczH2XLFlZ/gtopB/eMJ7mWap+0nGcrKp3M1zFYXpu6Ls3WFHdJp0vYcL
cBhuGzZXBkO0byrvieB5WM+lJoa0yN20QVLWBINIYyWz6ozdZEoBIWmK8P49TxrmRkPZwt6fo2Ag
gwjAt/SibMaiUHhsa3xzC2AUg0LKkbAppB5Yz4+JR2/kJ4VY02fcV3AZtBqPa3unvQlc14j0pjWW
BWJ4q56j0oIkDHYwBwoybW6V1RChZW1UIWF9YZT/f6EwA39vbKJ8KwonO/dX0tObPohaVcFGFujj
HhmgYbJYUchV6lZyWWKJsGL+TAOs2LvyA99V0XyKM0+hICuB8bHR98DayaJWhVzAjhzFSPA26qPo
qeueoQhTOAbFl7f5NTO3JqDAwEb8drPJFWxgfZyCE/nPCzgcc7o5ZUnN4ClqWLF2z01SiIReRjuT
uK9HaoANb8xo2SG4zjsqxh6azs70broosnyAvkJaebqj+3vgUWEIHxersaoXYMufq2kJZWpMx0Ic
3zrkHUUOY2irZfTxWqhbHheJtFjeNUJLIib4GMxrtZnNzsj5vFTRVJ7Bo4S8b87Fh9XtmrCz9J9F
Na7TJs2+sLfeLcCCfAIWf+qL/ACi6H9Xj3oUPvjnW+ShKXWnczOlHm751g41RKW81FToyF9U2B7Z
03qxMpgbAKvqRriSbNgHLQ3bSJMWBsg/svV9qTLiRLhbGggVHMbAuUE1y4Qk32pb3wA2RFdJ8Rgs
SK2W3V3BDTp0QsRZ4jfvtItZ6XEePvvHQBgXdLO1SpeVyfGZq3YjReg3hPHTW9v6M7MHJ0zRlIv3
mZvTMSc+L5ga34WYyVavYaeA9a7rp0k5+wUXC6l12r9AS6EW6OcVJEs5ewljelXnjs8NMLoc8tFr
9GFMVukXPsNmurbHJYMjqmnEEkSX1cWmETInvLWdnwW8PiQZfHe8HmeBYMhxwooWr+RdpHqNCVOD
6KjViieV0k1yn+7SQvZSt1fNc9rZSxE7BiZrxEd2fbxITjsU5Fw5YEE7ug1hUONEm0yshlbGBvnC
QumyXaR/Dvygun+//enUjNNvFb9gx+SGjELBWsiDP8CYQgwkr01dXAshZ6IkBh058tfIFjQR9yqO
e3gCzj5c2qBRfHRiT9V9HFFOBeHNNcLcoJklmddco3cMDb2jfdmzFUnp6yHbcckorNClNYCty2tf
9YhBAlb/zfUSQnaR1pvwhgFtxDw42182IGuzmz3KjR34XRtSjuu3inf12f7EA3sLfZ3SG4o31XX0
wArurkFou/S+9dKQVn2Wmvx9jT95Kgc1ixHQDwoyfzYAY4Wdk4UJRLjjYT2fRkQxNhw3AcfRoP42
cbHkjYXnl1/ijUSMNy3myG1E7xGirh4uQQ9HsRm7ePY8b+SBYLecQi56Hg7QAOSxVlkst8aFOORz
t9+BpPQjWoHboRp2NlSOrJ6kNPKR36nHKaxl3ATo3Eo11MkFpKLiXnmgDOSA/AeOAdTGjCHM/d57
TNCBqCqq3+AmYnze9ZMBHdnHq5+iG6JTu/EvL5fpOx8C0+Ugz0yVJ2ogs/I5voBp4hQpn09Lz2H2
X/A7Et/XKVMKBF004laOe5qgLvhhC9obbp1PBHAieL3ezGZgMjvfDsQomyQLpQtjGQHVOYYvLIAS
766bTB35e4hRoXu6oNCAAYSsLC0KX5zpXQJSYcx9wYJKtuX7fYUdN3eLM+bIyBtqb7PwKVlhEYNg
EWaaNBrU9yi/MwiLoJEn6PGX4UIVd78fQryVhPN3e7L9yT+x06zuTaeztK2ulHxDeREJpWAnwvt8
ngGvquvEl6q9w1mz/7t6DRhpHxTE7zLMLzrH75+l3F6Lg7pEeK3Rg563H+e3fuYu/Mg0VfCgIko8
ToIaRZCmi79QhuzWe4ijxlTgyX8EbC9kv6sOuGYUurQitC0wkk4h6ukLAvkThG08O5XxV8OwK1Ao
j2kB5ZMpyVy2OtdeYw5a9IQMxvVGaQd+HFBciPtHm5eLcpjfy0ucL3AIPHuarrXgqYvyW2WNeZg1
1hJnyUQWksadHMTr1Z/ORkYKKFYipMJVXiKST1wN3gPHncuD6RoyGsj3ASZK/svoVB2KG8CrDVoy
TKHW1G6ppB/nl+Cbqu1O43a9uf/8XiXJAIEY99PP5ZVYvsruxSAlmWeoXlLwp+17irnChTD4GFFR
cLhJYTFm4sqNvgXKPO4HM7+q8qU6dUBeb7gtChgN6V26nQuzr2DSpmd45kSt9B/ujHvUnIpzT71A
RU7Lj/VPUFf8ilZGUPBZeida32UHkl4qtAy1H76lEtZ1/9WRqQQVOcdeL7sGzPEymuvIzd16ggcd
3H7SNJ0+fkIfBQgYpufNuFD3zfV8ZfcAtRSITqYo5s9M5E+T5H7yys5iHrFWmfY26TDqBT8TcPBc
UWYDzobALuAK7r0BqZwp485yX70RGTiF2bi1o39Rfa4rMIrgc69VmV1myzliY0NLxnx2zRkDCXc/
ob7K7Ee+4UdJ1zE+HJERIaajcW9RF/XofhDCY4gH0sdTcpUHBr/AxcmlQGiucmsCEM8iOYo5rikF
BJY6envcz8CGtCcQ+o+bMj/BBw0ykT/qNwgbCpKl3L7P++AVvstOXN/5GAjqzkzublagXJE5Eeuk
UKjhrpwtqOvnN8jbbcaYta53EQomrnRy8YKz8fQG71j4KSAeQfuwZUMQ37QpQia3S79jT1v3ZOKB
IDhTpOsDLCLwJvmIrix6Zln8+UGLwngqrxlaFDo0/SHFYgCQxcms5G1Fv1vwKgws9LVpPHTA9t9N
YSweffqjdIT8k8hA4HhGL99PSYGANCNLG7MxhGCaAuKZSct2DnK0qztNIaTi5o/ZhfozyWbnAatl
/Jzl9il1H6d4OSHwWR1rEQj/Qnf3LcHaap8hMDJFnyR4cxERWW9dvnFlYYMDYRprY2D2S9atXYlc
LSq8JRSUpe7I8cD0k51NdKlht70Zi3JYGz0x8/6jfUqF+avj0OcnVEfn100s4CTa1/N7yEl+wvYA
7uvz+AMZcmw62/wGkj4wBYslLb/cjKZOTXE3yEtAu8US4kWO7B3yxOOSp7aYl1deFZcE0MYp653p
lAz8WTyviH0F6fMks4h3ge/RtsSE68amsFWCRDyUOgVFY54OtwB2eH3lyz/OGN2lRBNgJK0A96BB
r0aHvRgDjYjgEAF/L3vuiWVejLfztPmf6+Z2fsauSiJq/uF4Gekp01ztswc/MA+p5o+kTxxGdtXR
laVVblkuk8HliUDd5KADs8tXLq/xO95K9IjJCy/narFCl++pCP46FDNTB/PPXlZHxf8JsJ2MoDty
H2Yzv27db9NLunnp4p5oUMWRqhX8MX7dKzkqtK95RXK3Ysb6MLL07YLfDsQPRkei0mOhQI599QgL
6n9VcowHReM2dh/tOrcl6y8GoS4KIwZUS8yYlA4aOmF7cGYSxBa0quFRetBwkHQCKL+m+aba+bgr
Jjb7S0cXvIDQsHBFmXdPzsDM+tVW2X/x7LPtMWWMwq2FPYSrNnN+jSr/NFR6qsrJS91jgkPga/DF
venpZh3bBnB/UrWoWQYIqvi/TzgC/EmYdQj7Co7ql4LMyM/YwZcctJge7RfpoYpW3FJwsrmUzUON
K5Sx3EY1TnnnaTtP6H49VrOn/S5e4RQhZs45/tF96IpofLJHkh8Sp6+FHUfMa/89YHgK2S/91q7Q
mHV0bJ/zh7G/dZ2LhNublULvQSAZLWDS2Z99awf7Me4yjw+RHM8SHmTGGvqxUABU8PdH54eVWvf8
AfRxVCIZC/wiQKecvBCTyt22+RFzsPL6t4g+FNHDRsvpCXcWEPqqDB030ZIv6w4tjwSwP7n9MeP2
TU1888fP6B79LYQ78k14d97FpYRGSq4BTokkKtQf7Bg2vXGzCHVIaLseL4BUZz1YmfbYLAMg2umK
wPhAl79OZUYhsalCG/T9gKjMCj8juaADsPYmhv8vWCS/r4AoM+d0nO3Ax5GkGv3sxwQBSPBgPkuf
sOdM1jIUDNc8A+Ty5V31RK6DdV9Ppn0ojzx5KBGtNSxCk8Qia/5y30c3wMOJLaedgfWeC/nk0D8g
50gecrKRCHKt592keS9ZQ5kbPY8z3aXDwWBahSC+8AF5hhFYHcfeO6LgeFdLy24ZEaai/fdERF5P
V3SlJQnDNP7SZyDFQjj3g3HB6pOhuX8WwevmoSRC0BLnwY5FXCjO0VN28QLbyW2AUDBWGRo0p7MM
1YIEqjvrmZp8UVIyzchV2QL1m9c0ioy1NlJ9Kp+CG40qZ6K4nq9XCaFMYDFoozYua+yIWAGn4dRx
hF1XjXB+wsmOt6XuzVwsOctk/uKIK9t00/naV9WS8zSjav92BGLbxH9VE73fnVD1IKLXFituF/k3
jtZuMdmdWlHPE0D2ajGFcf9o7+SALQm6ErIaaHKbEF/IC7y5we277LJgXeM70wAJ8zZRYHXdaQDY
yUZzLfYUSuKnNeJ4Q5sHTD0hB0nIKIMddJGYjsgb613KkOIwNAHZnNsxi8Q0Adlq5Znb78vHwcEc
IMe6SQU+0QOPTWRz6ozdc1i67b15EluN53zCCeU9uYXjsnU/N15tO2qIVwIY7yl0kTjxUP27q8ya
ns7O5QM6cUtMxkDR2COLYPlH48qXii3nVgyvOWRxW09rI+wkTr9V3NufyNACtT6LtQQ9eZKQxNZO
eskeKxGWI988evNNk3N02Udo2mWDgwPGHHJol2c5FBLkY8CbTsqyXFaz8rIo44/ItGmunuxvUtQm
Q/QZ5IMXJPOwqViNfQoj524hwJ8F4elDDg5SxqjyJ0onJC8kBdaSz0zz0D7ljDsNui0HNOP6rPNN
t48iE/980h602c3rAVkRPvCguyaMT8gkbazt4NUpydumlyGFe5Zc16OOJvlAAQ4odzSEgy9p8ECf
RQOOD1Ttifg1UUAW0MgpUjV02+3nNakDdG1/Y/7J+JTOt31u0mbeawGxC2uGXrHaYuDTux8JEaAn
SqbZLvjKOrgkt1SlAg0wthx+70zdHF84ohwIhSZI0Nya+5nXpMIDvHJcMcvlp3qfLRRPJh4KEfcT
fxmKOIU0GKYJu1UZ6r0ruhePDeyiMgO1dYQw//m1iKJdEU89gT/jTbWCthifotrElexFJixUJ6Xg
VfE6QGPhYuwD73pOBSYRcDCtPBCToq2ce4jDjN/LWJ+zCvsjuoAiQ45K12Vq6qFfFax5grnhCVjz
WFw4pPLSYwdjh95dR3WIvSZ0WV5TfrkzK71WrSoGLMOks0xYrAyRSTdz6cmbIjV5cqOhjLnI3kcJ
2SZmULM48RCr1YLbBzhVt9Ci7bagPIXIzDtubx6KqgYVunBHkg+TkjOt0uEjLM6t1SqIdxj4yGQR
yXXJdfjHg83n5oLmPxemF/KRS4WOAge+Unq8G7vKTiAVesBTycgUQygjHaoUh1RE1QiQNurSajyV
I8tw742DHsUEfFG+Ko9vuEUfA7wO+QG/MyDoT3uZMP2qUYLSXw24BGWq4oalRqs1BvD8+dAqr2R3
Rc0gtoStoYokoEneXL4bVdpMe+7AyFmye/ikjMY9Z0K8tCbKv0gZgkycocJjA+dNl9kC+cCGNHH5
mHMcfdrk4Q8vn1MiM4Ml/upsrRKta4jQNIq2mne2jcAQlMtonGjZYXTDZ94QsQEFnYi1XAVaw8vX
Xxh7eTsJJYMPcsZ5FaKHvGBDSmLkLHL/eKyPNdO8N2FwQ7uOT/WDanFf3KNAGM15NYzeQ82ACgER
oW0SVeDYFen8ImF3Ob8jmqZ4l2UZEwQRFGcr1CbJy2mUKKzBgHHnDFZstg1Kq4+6n+VoyXm+cq8V
ILffF2fV9JuIlL1qPbYoNCRq6fw5BjJIQOkv5wNN/GwMpi1MnCvN+TJRivtwLKlCpuLWqjgjj6FR
H6Bdoj1Zs8omZRGV5c4UfjsgiNpcy+yO8iHj04kk66F2ni2Aek/GyFJ4p0QTaWG6PmCHAlgsq0yU
GjqY1vxTWtz3t8gepA8tefN7BUMTfqcViYXi7lEvz+iyhiMQvHUcL5hkLM6pRdzxdRg9tiOGbwwp
bI9+ETIuKyGLhF9RbT+91LMGU82VwqFtDo0mJNY470Sg7lZzw0uksYtjuoqldmbanTWVJHW0e10u
4DVDFpo6a685x2b8jKdymStx0BaFhtRQARPi49R7jlBVmK5SU6QBz204Owegf1Dd7NXRt1LdvDnL
R3sK3g+jVN7PycSk74Llr6Xvp7Os1PCAhZ8MCi5LDY5qXBSHbXu/19CiSwhYm0DvkLYxtjaDsw5Q
iNFSJgM8a1/6gqtwngXgo6hE2dkdBdrKSCkEv5CEOOIWhBUSo2FTnOfAUW5pDBCcPq2qUsXfkKtU
yqBivfemc+XL9P6KmqsTK2bRiyw2hzgehfqRniLnZaIb/Yd5E/zqPcULX/tUG0ipqHbBu87mhTwX
RRxRSg1AJPvlevgIQu7pEFirzdD7zmWTppKiNJ0lesu//GLOxWzAsZcLKzLu+UNcWcri3k78PUhL
EYhohx0vhO4UQbSiGA3FFX7eILnekYk0WgUbh8M/Gc6w2iWDZsRgNQdd/HS4XeqRd6IyKtGg3DW1
td+03qS3B/zIUrwQ28KcsTzoBhL8trD3kYux7OlcEF8rSZCB+rmLltqcrTIxC/gsJqz8erzFG7Iw
vId9ag9PoOAlRZUgD+2BL3KUPZkud55wgschlcaNFhSlW0CLzRsXDKRlz3Gv2Nr5fL8NbJ08Iv7v
yQOvU3qVNy4GUfu8UEzXQ4ac2c6Wbeahu0OTDz6fx+/dRtZdxOFVJNqoSQp0TYqgtmCAWqUx9tdi
FCYe78x59Ko7h4phrAzVPYe/vFCUBd+9JFFV89wiDGTGGiQXY/Cb7lRlyVwitwojxInKIts6sg5L
Ngr75ZT3/0ETEQV2YNm285pptni3SN3rmnz9LCYO4kdJ+MVOR7MSAavd+w0eendQrr41LAPaTu4m
Et7gsIg1sv1PRDjc2ObfYiSK5QX/oyvbHnJO0klYCUsk7ZIyLE7HjADBhFwcx/x/JwrxkmzE+mqe
XxlkdjbfI+O7C7kerXFEmxLCYvLJY7oQFFZaS9rlnuTU9bg5/SBKQNGstD/P8kEIo9TAEec4XN9B
qUAAhg/49fm+rBgADvTRirEOQsMOf8Sd1hNqjAjl7xMoZTGiXh95d33OcRSLFg7FmURSrstCrwiJ
g84j2REjzukWV1ULsO9b6hOH2NHgW+/YfDQz/zAIYM5/g+k6VzqXs7kQIab27M/VfIL/jg7TLKdk
GGEgXgV4VilQWM0kQJJgaFBuWRMMZekOcoRhQ9KpMa6iq0Xgqj3b+DQGcim7DCy3z7eYcZICY3qB
to6DZ3rzqbQbWirvsJW7qMpCkIrUJqzQXhyjBUjHHQX+LOQVEyZkIpzmmre6hK7DeMmwMICz5qTd
3ybFlbH12wZ5yRYbssBRicrss1eDTTECLzHF4RmTW7Eh1MawguYzr/gkwVE9q6Swpn34ZBYoG1QK
SDzdA4b7v20aIqavRMwwRjQHCfyXYYPUqElkx8evDk3dW22IteUM8SzyGQBEVuVDw6kp9HOZ9BsF
/tf4YyzeHKkGkRB0O0APs4TjxEX6tfwTIu0sUduEm52deB06UCya/h2CBvLnwE24Esa0gaEOKzqB
4NGnyPMFt7DhsLFke5l6ekc6wZqad7J5CEqeCqfnjANpFPMK/HHXK1HwUCLh9xV9TLr9bgVCp1CI
2qz+c511ihRVwCpAogTomCq6M4oS0rsJdp7A53qr3e+YsvKZeyemRG60JFPjsLiUnRI5nstsvVXK
4lXaLumXeZsCTPg/l4g3cM1Jp4HWCCUIBQrWx4e4E8x+dxa04QaXsF2Ys/P7JUtW//QQn++gBHD2
rsHEpvQzRRZo1lgduzZPwcza9scmdpmcNXWXrxJ2QO9xUPhuUf/ZgkXq6YEWm6ZvwzCQnavlmZe8
8LrBXHztL5jP+aVPAKqr9iTOQC0gLvKaYZb5ACz+X1x1sHN4muM7+UcaJj8XD2fjVIL8q/2lHuIK
+uMoqQ/cXzGeaJ76Zoqx9G0nRYPLvW404KdYwKtkgd0gWheFV+g43yWA5naP7CTQDxknFSzdgX4S
lGVdK/KShKaglDXXhYT7lDFYwF2CnIJaCnNJsgO0Hxs5L9CuQhkGoXtGYvzFoQkyoZaVWSCoxI5+
eybxDeKQOd9wNjXF2HmzA2v3BsLt/pvVl3YNf3eemux7KkQcBAd37YZXP3TvVz82wrH2d9eqhNrT
d6MMmVpY0GTmEOrjTO43rdnGv/nzTcq82czKk5Y7kCqH/a8yJI236UOb7xv4FhJtH8Zr1H9oNAi/
WyUnnLXaumhJ+e67FY4+fpz88wE3/ZGwvaFlOTbQfkTDdbz+6fknNpEbkjzKrofw+CScj+XNVwAy
sYT/vUJnL0K1xE/j0wTe0/GeS39u+UMlWip70PNtqUP0OyUzdXicmVBbCPao0jsCOcVLaZhu8bze
eiDR7niO+3WxjmwVrb0/BnNU97Q1TOkfkYFf9ig5RK8/TDS04dG/S4BxCNDV16KgRlWYlxH+Y1jG
d8m5cP6QNxom9M/lgjV4ccQVkTRGcX/XpS218WKHFLgxzB/U+js0Nb5WYjvVQxYv3gjORAQY6LeA
sd4RYx/8X8vUZn24USADVqobvOGPKgwPng7k1cwBGvl0HKdfF/kp7elpGZbv58IYXrn9SkNlOdLS
jNAZcWTOHbEmX9fxMzRsqf0dOCAnNuKYHtbFxqfHCisMLroxlcXrZJsYe0JrHVXSQANFywBPFzP+
Rp2Lv0bOYuephu20MMo3PcEjM6JrMKOB8jzYFAh03LjWN6mTVGvxBVwh1G1PG+OEZeDA/9+BZEPl
hABt/mdEWpqXRFCz2IO1S0fMJKAduhonZWb5b5A4Vz3zwmDKrVEDPwWgcDCRccJ+sdqJP/kC10n0
jOdZxGsdd403SnkSMogOEyskFZrqaFwVC41jBkPjcEn9GaVtStNqmF4E2IEe9EQAD6MVTb1UIM8a
g+eixpmHNi7pzY4sJaeOfaTxyVJvOPO/j+4hyW4Otwj6Nn5S8GoZMzqdoak1utqYIE7RwR6gIqlK
FMNjmjrE4hXN17F6TIWcxU+c0bokLCrYKaivrVI+tJQGl9SkGCcMLNFhT3WGvUoZ8cpmZL2sIEFt
yCu/K0aeuTgi2bdQjzpLvQgvYRf30PGhLLEFK/X+k7n6BQqOJJM3qHyMclhuMN5TJ4ppUANu20DW
RqYt4q4kwyJAj7cMCwFRLB5nbmHB+nuiBl9h7mBdi1phX4HNVPTibsDA1H30zNvZCHnXAeMrvC2B
iNxf5HwbvZmWiHrBSTF1l9Svwhg3FT8TVgzICZwe/452n+ysG/vPYnDiaKgld3JwPWn9/AyKNIVJ
h53/doWJ4f21x6+KXbIyrPwzY+bf7pWZ/puFwvK4dq4OVEfpgcMEOlcpKPiL5kWYSqmqisZ8o8Ea
FjAV0A6pm/To91PdckNRuwi7X2rSSB63rB+lmIYZlenm3zA8dItRpFg6qdkY5R4v/XF/4OnaGVW7
bzGrYxWJTcbw4FkpTJO1cneNMwKeZT9rc6EorD74zbfIC7OZ/BU93eUBAp6wUO14khjOFJKLvvJv
kmUVlU32PBHlXY3kkM1W3Eqr29aGqjYxL0Mx0n9dLV3RKDRlUNmpp2PMYI421thUf7YlO1OkjU3y
fOhMp+qEoJGlQvkF3es+1eKmp5CISUCFBTYQFriTOTz+sed2bfhFJMZErDY1KH4enALitAcVJpaL
Y96f9TcNCSTHj09KT8MMNIw/5lxyML2BiZgwSaJtGCsOvGtjAhPgQB8wbh33Vj9VOrHZJDrz45Uv
L0NpZVdon4+CLhFavDaphmdJ9T8CX6UQg0qQis4xiN6hi8zWp+MdqQP5wxE5Eq7D5A8UHCD5z24M
C1eHorbEXqcFcX0fwftevwnRH2cv6NTWaeNj6ztaW3RXN7GerDddQb2QV0xXVobsaTd1E5rZlKla
FjHYnVKfebB1RPnl28JtaQdED4cjQBgZXW/MvQ1+vVreKk+SOpOvMCmT7D4fEdzwV1KFfupf006t
xHx9BqJE5T71A/V1q5m6oibU/mfslcXnvOQiY+gwV8tGmFf/fzaRbsiBchkeUzkV0Yj3XBTfDnNm
o+o8O9eDNj2I6PZMA8BigTKuq1u1H0l1sk5uFIqzMtsJ2sIiOQluz+uaecb5lYLWFj9GDOF6fUAx
lYqESnxLb3D5MXaOPxURcqA+kzYAoopEOBVf43piDHBcWSjb/hwCfziyIxhyPcJ0jRtDJYszj0sX
Mp2M5AFFw8uia4ZXTbUZ2RFMOmIFZf2weNQpJHvGmBvmIEkeQRd5uYfOwIBzGlK+mufKuCBT2nX9
ZnHjNUA6GxaJVcFwa9u8ylaDLCazbhsjRQoIToDNic6pqXzJL0p7Ync0JYDAZoyQyqYebbzGMVvO
nt941BvREveImeZKVgK6k9DmSBvU3XL3Df1n4GZoYNWWaPKv4vqY+xvXOWHdmdK5dcCpNkoIMm5S
Ba3n4HMd8AOKDkEuPp+xiLjVUi7U11Si9iOW+jteM7JbdKIPL6HDQFOn8/IZ/Tw6r6tPboYSQTaT
uHAMtKllfywknHDJr36JkV+Ufkc+ZW406EQ/EidLAU0dsyd0ambAa8rdmzhxavnXKh/xQNpPtQBD
Wd5xLKrkeRdNT/3YY8czRVSP/hCrEM8VU9fuEnMDZqrZTL1oXA/IknUjxh0fdEhYQAJjgZaZF6b9
dw6RSoeWHaMzNzh6+AKlBjJWvK2R1Gk7mmj5Kni7qWsp4dxTLi0ufTY1GJK86WTLi2syaj6tD6lg
xb66EAbpFsglLeonQJC2PUedqABKTT6n58MU/W3p8aXvgFbGfd3/c2pFS1CefvRGW6CKXmXEScOB
ms3tyVp1lbkG+PYkJmH2Tq59rgNtd/TfszFQa0avVVusGWnVXs4sy/k5F7dZWgrGN8tcY29QaK+8
56KpG0Ry6taI4kdxoLm2e22+wp8EjTYJoLYzGXR5HBKikLJ/gHwAfZsotBXYtCZH8LHojY19Udai
XxgRDe0HzyefY+ck/UZAYAqJ8g/holLY0mHnXYWMbaSMIUKTfYjjn/a/5gMfghGQwNUfVEm+bfQM
a+z8YskdHqrbxfBUrmoF/mYU2UJ8mF+EyOVsAhh0FYsWryCtl76Dl98sLyGZoXng1W1JH7wT+40m
/LmKqIX+SwMJIAIpIf9BSOY5qVp8qG2bZ9EobIDsLudwoJIeMfPy20rhCRvTq1Oj+dpnmM1VVy38
tlNRaAnaT1AyVzEc+NSnFaqXnop+rr6CmcS4FZxTp59mIAC6LL5XsjEd1Q4n2VyBhYBFNwe9avb8
1L0zubUseGydE4j3p3gowTgkfvjriHA1gMcIRPdZIw5JE8eN4nEDiAW2qMBmcuiqxTRF8LMa+8fx
gRyJ8gOqBNkUr6sl8QkZMcWt9dYbb7rdxtz38kYwE60SsKFpOmKt+nB8fPcyr/GJEwY4mYFPoOXD
ob9gK6vLBdqWZ/iIo8Js+lFS18iDG+PFtkrLkeSbKVQRs4oRu3eIim4sjoHmSqyiwch5IY5ntEGr
rMMObPq635qPZYkNj5V6F12VuZcF9xlrm8aJV1tGZq88nwc/963etr8Ff2VKo+f3beHrtF7IQKUJ
u4E4dO3BT2FaZwNxLo/1f9vPHJwK8DHnEB+USpcpv4S73OLDk+k7OTupawIVMrb6p/XA5VQXYT+t
yUMVVLXY7izSkADSH59c/uOMR0sRfqE9u3K1/8HwfF8qkuVinGyC/JnrrRQqLw3tWuOnr5/TWVP5
+1DNySHhT1q5napTyFQEb+zqzS9GiY3aNTmKjy6NCLWQ78c1OS9n5HdZXrBW9OhvmZWJoneyENJ6
H6AVsxduMX6fDdJuiO3BwO38JmfBAOkdv84XDtmmPIQgUhI8UT6TGzKw0g7iFGYeXbI2F5/b2vT4
JKAB/Zok7edfHwArAyGcIQg2SD+J3hS34odFp/C4xksJLW6Axgzd44ASCfP4jgkwt8ZlU/C5YNuz
bZ6+GPdR/4ndyOoAD8jS1DWhrO9aQL58IzeM123eKflfv+wLuVtLefLDwNWQLwWDBDQ8RTJGUlIf
o9ri/mg4/UcBwq3sIdmP7ngLCJmUEOevSKUbjkpi4FW0ZSU1ZNEnIowyAlgXfNtApoe8cwqQp/wd
xMRJhIFvbIowd2oWNUSA3ECTQdr4kOnLJQJpmWNaDzHXiwIhrktAa9twYJublReKwbt8oqPveW4O
XPxjlgFN2mtPgHu2WIPX8E/DP3rSmkLCD+zzrC9UYHKtSZrp/KHf0rhFgV1ohSqGzYIsXyB3sy2i
FgEbGQ3uRr+eJK5erFkc9DhGDbrqrhiiMHnIj+d94fUI/2fmAUsRSo7Pk6ns6jEraLzuuCFjc2pB
H0nPtBzEMtwZy9T/nTHGgkuqNeeC3gBBNXl+eXZlbWtFwpDKTW0CzxZYGjYXXBIXLCS6+DPYQRjJ
P9f/29q/t24Du1Cx/MbsDZbq/kPsU8R9zpNa2/sFRgnB6UNdFyoS0rnbC61AxbmfpjTPSpE18MHy
hSeiJQaF9oS0WkHRSkK5P4XK8gNgaB/V4dzcnwyzAvvI0ggP5DkfYNqmq+K2RUMm62vh8JcUaX4+
/hAlVawgadCx3qqTAQ/J4UJXmA/3o3mMU+wRy0Hz3TrWPO8exBojKffcDAuUTSSKxoLShuv4g/bV
FaoHDQkhFLUqV6CGpqHRvPTu4K5UZLf5nAXzAc30C1lvMlkZ4bzWrjGNyeHaqVDyeAlSeP42mgED
UWNzSwqPCKvCBmT3kRv7tEHmyiPMCDjU3wtMqyERKwh4zLf7H+LaOO4LZz9nbNYtgmec33px8qjO
0IaZL/KLIP+w2RGosIeWj7d+lVXenzo32mummLQiHaCUqRNi8JqWhQy9zTqiX+c8b2dP/X434+S1
P06V/f3YkM1D0J7TPGqlMMK6hW0rOADZB6V0rlkt/BpVqSKFnyUAtnT/5SmPA43TZy73N126wJvq
qQc37zzhA/Lhk+iaD+m/96ecIpiO2a8da8TjwZGyJcdy5wgbmGUIHuPgD9nVKUIDInZaddgckIVI
J8rUz4nWfYNXifxo2rkd8e2Gt8k2WyYjyJQjgYn3gvtsB1tAs8E1/xRzCFbyoeUOGfyqWGQwC3Wf
B4Hcv93PObRdG1VumNdF+G3Y566ZYPmBL2CUfHAvNNcD9rJM3cV8sEKdNyq3strTHEBnb1hVN1+U
HQg5kmhVwQTNaDt5Zszumh6WMxUAaEBhUPa1DVWp67xXfNIxskXXVbjAymHylin0o1h7cS79qRPH
IOrguiErNb45r4Z4QUuKPYHM29hSf+1iv3j0cbi06e91Ifcut7OSMJPamWnlDP2AV5BsT56FSxbS
Oo2Jtkfu1QcbBUiA7vnHcMTSHEL57uh5SFB8n+k6INgbJ1r0Hx+LAUDlgi025kJ6t/9lFYkrz7pV
cVYLiT/hj1dfercDmxvaN9KG9GCt5XtpUImNFxagsy25/jLIb4n4EOiWqDdn2xDzgmHpDlaqTY3Y
uF1YCYGSU3YQyr6sVf3AQw5kTgScgMDnevX91RpDyIrQi1AYYkRRzyDp6f6fzWY7yBWDsfcDdjSY
XHdPD0X6Uk21YnkWu663eGg1zjZlC8pqKacyUKGLkZmIPGwnL3XEi6Boe3dOKpLcHKlQx6bLQHDe
eofpyW2DdGWdPth5/5R6Cdd4NhexbThVoURG3CRHmj/55qG8IMaFSLVQbpr7dgmf2/K/j7c+Cn/i
9z/ROEmShsBlrzGv+kBoQvsI2QyYqzSvegnneqQbSjp+20X1WuxgekQrLOwUZhfT6U+SmZyudxAx
kTI2Uo2z1rpvWAukFq4VH/4H7iQcXfi+F9j2iq98ej+g8KHccBjOIB5gusJKnGZkusAyeSZQPZ+1
aq7oa8x92wSsTs3scRHxUjb9ds/xZwOAitt2vSQj/ajqRRcaCcuxMlNn4qt97nB2gbYWyt20wICF
7SrbrREJbCiSFI/bXdAxUShydJgo/3TwhICotgTWwYNKz5psKa7KOoLCdYhwpfiSg2Ks5ofZuW7M
AvgT80vvtcNmx6tLwxKiB1y1pMHK53psPRcBfpgxhey9tNuQlerIbHoBk5C6ERGZ5GaXSj15qKGG
cb+URp1Yb+tys5r7Q3fY026U+jMF93SuuaYQfzO5aSyYgQ/3/XUB3zAYxVu792nd5hBBgCxCUuyT
MoeDbNxU4iOuhLys+DcY/Gvo8tDnPg3GZqnDfO9pQCgm1aQWUop5Z755qK98qQ39q5RyIMBBhou+
SKkzOUtjL5hAhRBpdr+WJE34lbeXYVA1SU/Yr07g97OBMK2B8WK4v+XXqK9CJab3Go+RQ3UHXkRi
InATVj/rupfOc9JnKMpkjg77qCwXks1kQfBHTfOJYd0Zx1iQX8c27Xp/mVUnXBgkm2rMRE37CvQG
4lmN/vhjnjgfMUdsaN0qRNYjxPtlTEY9Qa6qoTp7g/HaswuOcG1JDV3k8WJy49UO3e0DZJa42+ZA
tSMzkabuP5BfV8RfrOP/LBh0H0EIGHZSTgF9eZcEWfLE5SvD8lKXGoZhDIW6vFl+6KJLPc8GJr8Z
qTBRcuEFw1CgMZ6YlNgapYAbqZ+5CDqYZ1T6FTKDqiOcXKifFw+R8w0RmesOU0kbCg2DLLAIUgtJ
vFcN1+tsssQRG2PFBCFniMgfHP0A8ZCIRQIuc2Fno21fND1wtZ5F3PSi2X+MziRzUOQrNOUH3D+/
r8O6vVB7IeWXWJKAB7S3wiWizLVS0mhUJA8JpnDERS2WX16ibOv3nVMThogdOXmCItQjDrDihnXC
SB+OC6EIgAezG3PIx8yfNFXbyUIg2OLuM0J+dVwmZP5/Y4e18TXEXWRNT+Jj/KcaP/ccLKXmGU0R
NInzIxEhBZBcGlrWcE4xxcBBuLrCjMy6viVk/wTuRSrzitKeE4jrTL3K1bSLef4HyfidTz9fZCQJ
mR8QrAtjlW5Vz5fwj2bMR8JYEPo0dOL+ps/7FaHAUwcSEQK0A+e7w+rl90DPYZalp0dq0WCPPmYr
Ag/TEMeEube2rjNR39fg36Kc1JyHDC/7d1iF09i1elsv2m0wsiB+FgTyfGkdvbm4ZVtg/B3lEzNC
tB/YccqVAG2nNaxz6XSIBtk3oMR86dKmE3G3wHoXHETQI5awVht4UXIf9nF0guFZKcA/48i04t3R
EZj/ANIoYPNyLICjBbJM5sN//hJK3cHYa3JsgO/dM0kLrlTcQFTrq+sZDPBQbfqSaNm72o94u17o
FSxKBB9J7rXIND5pQSfclwlqrsR9wQvUGmKBzfwqXYPxUWf6RhpWdVg17JaroJPPnr/RdvkB0Gx6
2X925968FkRVcVzCCuDBA3mvcmyGCiOuvRAxgXlJr/loExvXrKgb+S7d2Df8sjzwSeBF7HkiabWF
la1Heu1M0E1+POZB4Uv82/6I+cZBUQTBJdYeiqS5ix2KidAKcbMD1vlEmsgUsTqvek4JhYEB6O8F
4U42naauDKpRUpiuJXImJxovfX2t66zIfeDfZCFsJXJT/rfnimiaQC+TawKsV4RsprKELee8/hzI
80T/spTyRH01kEkQOffPYRbgrZkTXB6NzZi7O/UqYr5i0gGME9nWPEyYwPVMGNgfFuN3vk4Vtt24
J5L0ZuxZoUalUoCm1jD2FDerqare2trFplKDX24i8cGSQ7LD4oZ93NZF8keWwIKXADxWp7Nixn1m
VR33f6p9lgVxlduF1NBiSOsJSN1xC3Q1XLQcDu417bPtWJGqvDNlbCKqLPeFJluegbMmdSK5I3ju
LJ9Q5hZ5AI3Q/ZWRGQ0cnrtIJYV5c7SRCw4nhgOCtDLyXmpR9gOR1FPezdcAUtFMhGgqfVfPyMK9
1rzhq/X0NO9E3NwFQmsT6lrCwaS5ZtOUcELxd5rFOxPzLK4U9EdApS0bHJafr2IPisC6cBlSW0qt
BUfH/vio5whN95T9eo7TX0N5z9eykFN9Xm62naYt6URWOz99mFrKGVjeu9ZYS4qo5SSPT3E7cWBy
sebjkmEUScxk+8ZXkFKvH0vzvHb1//mp/AC1sOFqZZjFMtoqFDn5VruMk+jEk2eLOjSPG9fBwKjJ
yvmJmq2j4WACDkev6I3UnKtGKcIfIEA430bWEL6ghuuQy2y/ypddkyWIu6OnLOJqhNvFdI5La97q
IcIZOv6+p4xeAfLjxSImg4mSTwokKTLS0EILqyg7WLCnnvEl6eSdL7NjNfJ2J8UTHny/2wctlwd1
Yp6S1TFa1+cbjD4if23Lv4LBvPaN6c7U1ODYV8wb/VHa5vaQa49ESTO5zv9oZLJF/jvFYs0exvkr
+XlRL5uQCc8n3PhRKtGZyAHWQnLZpXWh/S72bB8k1kuWPAKaIZgFDaWifJHCHek3mWzeqyc15AbT
uYStrUFp0LgE3O01PHsvMr4je1rcU1+Ib8v6dZVoA3GKqD3qOiiRTc7Dgki8u/wp8kLGOQl6RKGx
28gSLef3q2K0hGACD1XQt6+ssxY5SlUm4hhcpYxlHsEzvDs8HR0dbhjXKtrooYAuTqmmbFzoGQ/d
dmqT6ia2jjFTgQt48km6tnYUSEkoQRDQybHZRIi9s1hOC/fJahgMtlgVQxVbhZvYNDKcCa9dDnST
JALAM075lR9YXdM0fhbma7Q6HxN2aQFucJY9o3DOSX8fCfUjZutUUf/SMweHHE2s0Pz675mE9BmG
K5p8Ax39Zns4K/0EQ0drca6WW37xk7unj0+z3ajTDpnD6YGjsCcCuniNuOLbJ9NTFOZgG/Xja5tb
QelQQF29imt6albgS18xMv2vXEsR50h9WxfH4A5lv6WmnFhnhFLtKoQuW+Vk94e5/fYzknIl980t
rV/kloYMEHvZtQJIn2jX6DuYmDsu3cmTeZiq/saIEwLo1lf9S73DOflvu7Ky2pvZVKAmS3LQGgp3
hYX2/wZLG+w847NgbzIQSRzEM+HOeGWwl82ErUuKvd096ZW8Rzo0KaykTwuL3fmm4BGz3WHR6MGE
yezobS2xw5q4ONKfZPX6r/ngBRRZsA48F2DmGw0khJe8FHJbKZLkOL5najK/EIuxt/PyQlHoB//Z
X3LxvwvrOmrpyrVd4CC4rAHjMpclbgJ5Y411l7zqzymLJQc/zqgvw8FQyjEOd7d2LAeSTBArQR/U
8korkYexWbkaPbezKhvsdMNUW8KmTXixKsPTuAvFY1wSjPF0RhdnhAJDwYaId+bEa6gF8WZoW/cM
MJRhc+MTV5pfZy8/npFEBmJ0wG8ZKqc45oHPV5IcjgfvuivJ0issWEhTFSAeqBXdFGGsQR8CT0gB
pUvu2lZFYcSA95BT7FgnUSrTBFqzBUI0IR3lXrWsXhu0J8IYu6wvKQ9LLrxkxJhBlKvGAHl9K4RN
Fo8Xw4jWFt5AU3wHom4x3flwf+yukY3Lqwq4xryIDLstNgnGwFloBzDfuASgo8d8WsxrLhXO+BvS
459p62Tk2isbZcRW63Sppy+MYtdoOlMzNjdqc5Nf9sndue01Z2fPhota4UNNdLth7rx+5rqYi2Ft
3QMEkboQqWf3zw+q1A6FMRGsBxzwkwIc5SiCRgbpZmI+9rfWUBzAkuuhBrAr5Q7icj1b47H6SScn
O619h4AaBOHdg7ERnGC852rLHRIlEkh0HnTgwNgezavhuFAyGIpUn9SyB1gbd8CZNwLInPSlmPoc
OXq2pP6kcsUWQPgz9QbgtSrsp2d+kLFCwjWvsn5jZ+OKrO8j9HXrskzmQFRioCSJ0rl6j5kBBckU
dsPrcfqykOWm3/1mQRY+uaKS2IHkfBth0bi+gYMa5YqcOAwskY5ztdwRUVga3paFRPYUMWcGmTjB
8zCp0ej1ux+kgSZS1TFFXNVnUgJ/upy1f0S34yq3BrFXsfZhJJ8VTeN9IBgGux+ulLSBtSr+8uvp
9FNzuKYZH9/tp4wU3wz+/M6I6yu4idWnQvEvMX7hMJiY1Zc2NtzOLTwftcztOcMAV3q1hDWTPYp+
UJBcpc095LmCH/D0fuGwkWNiY7mzJeBISGaSFQjrdDAfg7LoUl1OAWEMRsoHhkeVnOpoOCOBP5HQ
lpZXCTpf/QZCjHN4dsTthT+aD82JnCYMHVwQ5zJCkY04T/OxDXUgyYaqwNP2kZMnVwx2fn5BzWoo
IcbeJufpsurXsvOxCupuMuwj06KZpyYSW3wUGd16RMJapm1wZxjj4HUMZ1W6OlDbAhBAR+07Julq
1edc0gWfMZSbYvep0zyREXSbP1Za2CukV9fP8fC0x2/Xoaf3oyjykWLH6STGFGk0KBtdLRsyqBl5
Sg8Pd4n67H9H0UJuwLNJ3svA+WdPAI2Lkreea30WpCPJb/VSHnU4FlfeI9WIK9C7FVKDHXBXtaAE
+Y6T1RBeytMamVz9vP/IeDZ7H1fhHBuRDwkKejbjC2kLqfPOg+ioW5uUDaThFUHKWJgtQWnjIvtq
NXOBgUZohqmFaUw/frlSEvYOBAGMxQBXTLuD48ms4+s/pk4jijsjNI8jA5Q1GZYRXSGtBBBhhFjn
xOEMjrrnHeNOJwF2+Sjj9tRVVuKpteexLJMDZKmyTwiii1SfKR75b7EcWZ1+hIKivjBNt6XfBU6b
CgHMkxn55eWHam0cu/j+pjJTyPxKBSft4JmiEZomedsKxYabL8XaqFChtAGy6TEZPlkoxSvZS1No
q39jxYQ/n6efphh1tJkQbKYhtyzBY9KxS81Dl87zu25G2tU5yttO7s07kgkxIgl3PTZQXFxg5Y/7
7QxDMb2bcnuRmd7cKLSbDLt/bL78wLjPjanXhTFGCj0GYgr1q6wWrHzjH5vKLYtdVIG7gvOAPU2n
m2jWivrhNAeMQxpUkQui0dWYaONRMTggMJN4Gkjbf6Qby4L+PFnG8SXNxckkAZRlAG4420IpkyH1
Aw8CySCAyjNIZYj1v0b3mESp+CjFjZv+sXN9QAdYKgzPe2vcm4xFNeRrrWHl/i1HHlnaStF3WSad
C1QpZ8Ae2bGM7deXjK0TDQvkmVrEKyty6MIxomztn3lXhBoSlPdEF/j93ErGQyzHck3uWZH/d6FP
hZuBHzPB7JmvYlu6GxjsGJ4LOwE02KKlX7pXIKt3NgWz3HczpEpnLBGGy9uTC5xVw2f+91KqOfwD
WC9Fy5vupMaAOyl0YJMt88ZhqwGbj+udmfYJvO1V+Gifurn0CgTd5H/LNCKqpGSGvH7FMCVC+tKj
dUMm8amG5Mm+MpdDtMDAjsRADmtREJHTKV6mmuCesVcIphmJkHkbJFQPdYUMwW5RF1kfJMDzinLC
uipFmdqhvq/+pXBAxr+dMwfDrgnJPYqwWSrLLwNyUyp4A3+MbB11Q4CUMeHptwARhFFvZ416NbL/
dZrMkQOKNG3xfSnoX89Od3GsQAd/UnPj9w//sdoTlZPuU2ipOGPnDIcsZUkuEzqPbFvYaQZPb7WD
qbvG5d8WhICfkPcyO+Y/YeqpIewNCMNmeMf9ynFS5JK5HbBd7X64VVR/2AK2F1+jggOrkHfHgIdK
ArP974fKEk+Zm6aRMJ61TCoFOc8HtIgxIZmohoqfBYqnyWdY+qdfjGeUjuzddZW1Lz1CmCEHgO6Q
3/jyklWf4kfRnZx3NMWBxAxAwFhp6VWepv/XysnmftUIx1oVVCRhZkRxhVZDIdwQwueh9wiRqPWR
Oai8ZrwKGA0j2CKcteqKPMQv5C6Tpn/vepf4wQq9+baWpinI0h8S/R9TjuHDruGLH1OLEmynI3Q+
EkJDCyUhluIgeWkNQR+o5r05IaWwzPAwPh1Oav2oUxwympRvAJZynZwjLzhuhFoYVGeFj2auzc0N
KpA9ByNxNGKVvNw/ySlLaLrRZDnG2X4ROb4GRh6NR5LAwUfh2hqCIY/9pLCt6FwIbDKSisE8a/z7
qTCtzCUgXKY0iZa8x3lm4yU3ALcwWqFaLWDjMkLOKNjI0c9Z6tiT8c1zvfgCGXa/hMWE+Do2OEF6
drJUQg0+1JDgFMv8Uu1+hXOHmUVpP60IpkrjSQbcK85Z4YMxvPypSfcpROk6Mo0tWHMAkXnEP2D5
ZXqk9CG/nZ237tloJ+zOQf065+O3Dsq7dCRG/2hUIF/+O5YI7urWuSopO/ZB5ZTo3OUUFbjVxo6M
d+yGwEiIdwzY4jtj9S2ExB+bl9dL0xHB+AFuTL0LuqwqqORECPKCSyyDONk5uNWRp4AX75L+UcO0
sPPFjqv2aXOrnEI6cKJSFLyT2sv+vGnLZxaCgZ4TQgn17tmWB//KuW2gClJbk2C55TrKZFYmEVVX
O81MuZJ4P+9k9QBEAokGIZOx0Fplgz1srYMeCAIf10nOOKpSsLOzV0U2Ahr7kVMAfxjFVaqde4TX
E4xhmOHmuEEtpwy2pXTSbGhIbrzrmCdZH1Nyk8j3b58yTUZ5AFKMBGjuq4i+eLSsEr+VLVY0qtrH
2T4UAa+BQZjUeFBkbQ9/Ib7hJ6BN6CyxssQVi1Q+79xgjQAH8dKpLK7lJlhrT+bKG7VUZAhJ3X4g
jFGmNO1RcTOFqBGh9tvSLGSp/yTpvK1zLwWvBGS1hst3r0z1KpA3WPIzMUrCHV8JXPTT9ZgenjRQ
x1Y/sCXNa7CicOLuAgCGf70UeSCiUh8RPPzpg99xLLMIm7ebUjYRW63t7s7SO4XN0F333n+TL7nd
KRbZ6Q0BWBr4uM3qNAUmAOXZSUoqlBI90SPqqBK49Wj81UUQs07+6rUkb5Ff0hJnbMET4KiS+NZa
pJk5cxsnQ5uQqjDuua5x4dbbzDUO+c+bdQI5ZvES3ZFkYK/cIOQP1NGiTY8ZNpdoJ/6TDNexmSp/
iBiM5fLb/8RBdJL/gyzmIb9ODGmt664yklUmiZe4ylyLnVZ4LtWoVuYyT4uN7cxv5FG+/p10fjFA
I/V2071GYIl+tGv84aT1/Z/cNcq+Z2IctOmDvLkig9lVwM9l6ttPG4KkMPg5vDX7Huhs2ei2wO5Y
ITr5uPZB+Ac2enyGEdqsQzcn+457mYRltST7tb3tX1FWtS9EVgURAxb5/0YLiER66ab78RBAq/4O
SkWqf2Il3y+G58/dnt+V2uhrQg31kcCELTWQM5PzrVbLpeUqKHNQM+U7m8XZ+6pNIR8OERrV6k/o
92JOWbzI5z7AIZpEaVsF+22kGvafklGMBLHteQNlkqRbOyd+2S85LrokZUr7m8ZfS5JTMrj1WoIm
UGxmIYZES2YMUebtQYuLuTqZgB3lJc2894oBFCp3BhOXq6jVWSPZbVz9iRtH9YwhEgKYDilRI1wu
i1c6mfjILEpCTnTfN/1lOooQ6Zg8kKydjBJnfsKojbXnmUyU2Z6OyCzKU4t1HuS7fZjkQHppmu/O
Jse81CYzLCkjiMhA/aXhRZuSxJsIM+IVrwfFC+kT0Swbo0ADzpcvj8ahZjCsMhumW3HwM8x8bc6N
lFE2UJ2WUPevQN9MN72SndWiYLgJ2iSypbmDEbqVK7IFh1ycC84neVclU822myheqweROhpYLetM
9Tw2RWBgiEuH05AJ8bVHD4AKtzzE3IWL9D5h9yDwWSblziRiP63wOzN0DgFJQOp/I6eWFTf4vNFH
N+8WzAY3TXn1SyATh7ekCn8DOtjwMCItn5fcgFenYOptTlA8g2osvZ/Iy//y8t7Ut0Am63pqerKr
cvTnsyMqBpNKFM7ZHcbjNDNHdwxEe/c3pyW5GV6+WhVYXdbOQZYFbkcnhbfE6sfBab8xV7yy7dhA
KpnWescKPJWivLEtkpP74ZmOvXBVo92zKqB2hk5d7Qb6U8vZtn3uXBSwAYUuhdjHNOTmFSJHd/c7
9ClYB1rmsk6nvh8QKmLXQDlQKBcnv84y8P0TDMq52k6MYWEoyxFAgWo8hxrpu4wbp/fXl4b9S9lg
3wfUz3mmXRfK7R+6PfPJeRrsqUifVpu6IowfinKG79Ht2O2TlNfICKqivD2Mdpm9lO4gO1/7/dL0
kwaiZ4h2MBBXx10wAUy2ts2k8yLxJ+UgSkGY8UvAXeeic9PLOFTfZBu+PIvSwRv/gS0xf9kZjRan
Ug/BVeZd6LqdKSTqY8HazWp79fUzxsupZT8VWWc6kGc/Y3hMh81ZUnbr7cw8ejHdzW7Tef4VVW0i
W89VPU6RsX/JC+CztiYKIpNEgtOnO2IOHRFU4yiDnZ8WZLiCI6SLU/eKsK/dBHYOcZzA+B8+cWXO
mOWACvtJX5rfW3KMV/iAHwpfN2CrcQ7LsX1NbgSrW2jFNbSq+JYF7RfjUcnnmkrm1Uty2hVPJ5kA
FCPW/B2o5T83nzeuVIVsd5QRBeTGjduv4Py5Rubr/Xu3MOkLcUpF7zg/HJjDp7wMfhQNY/UwegsP
T7zprzk/LX2tHWLne/57oqW9L0wa3KP+O2HMl04AeaqSIe538kDLhYWvC6V9TAeV4zLQg9VBAEuo
iZbZO82geZYNwsEPpXQ5ituSnBTrAEXRgrgxKNDBqx5Pmf8M1NxwuPRbDqFaz5mt6k1p/jyvR/lZ
6EH8zZIgTabZtk5xb8V2/uD3X/oE1iXSyoTrWZ3z8xztjhfscarWI+DAnrXIQLc4MGrqBGO/OtSC
/b0Q5iakOEqU7AHwv9eZArTlzy5984geSFnZPzjcDY4NyzqBz+BD6muhvHVSccdBXT8v99l0uOoR
Kb0IxX9yIx4uu53VK+fcRiJBlJSN8tGXOR6COCrqtyqCsaElD3j7MeNrUdbl9dMbCiF8QG0wq3NV
D5xSspseOiRgo4fXvttlE5SHfWJpYLpFidXk1Ct0/YrGxuKC3MlLPVToVEh3arnGldZNTyhIaPUL
nb+u5cCv5D/ZZUgLzEBqQdNZkrVFBL+GrbDnqYCTJkE5chzf7zP05vSZLetWsYmAtuYhFvIFOnqV
5Yzt/N12v+ZlVIewBoW9b0GT9tyZAC6xdEB1I1N7yMQP30h+VMzrJWjpkeiJ0bzxZlpdOzVE7jH9
MWxk4/P118XUk+6/2HHg7J5Vk9MPGAQbi71YqKNufu1CcS77D+ZmuP1tSSCust2ZtC3bkJJaLw6U
iHD7LJR5sH6TL9ME7XRGkeRP60G0qJGI+KNNYNqfMnksC2Hd7yFEUTL9iJsHpEDfC3EpapRvWmYI
tO3hcN2pPXAJLWsEJ7hBjeq0vPzo9wOm+8F1NizO5Ybr+oyAUuvWdn6D2rrqdil1GYGSOTfRiOyE
Scuned1XgT98ns9TXm6lTuwhYruH+4z6DXmplvnTUQAyRS+NzYkyhbzZcHuAfnLCvfaHNWBS+M2I
iY3nenYn6U+Jkl1PqomlQfxyYT/t6/JOxGPJrD/sq+M3SxOWhp76gh1jgcGnTsAPgn4GA3pMZIAl
39WDQlX813tf8RUd8vjbB95DVMbrwXTQpGSrZ/mnQpQ6sZfw8E0eEI+G4A2ARYkp3LRV/p/TSeKp
FW2D+yNFfZ6ATd7MFqE44wmiWKdZSRt8V59aPftn+p8z0Au0fc4SYXps5fmFsw20IhtJArwI2U3Z
b6jTdXtbcyH4vm40ZWzI6+wDA1fzV4zl+hYi5VeRhSPRFh8U6iWKkmxoUXVyWQi2mhOr0XWXf1Gi
7Nyk4NG5ZwXP4mNWLfg5VC2zOtEaxL/2Eo63Pq6A8N99U146MzbANBfv9I7sP8fr79mt0QJVvB6d
cyZH7QX7y1mzBmJZS09krt94s8wmgl5W90u+ExfqQ8r9Lwg24Bnmx2DLrjJfUyG9PJnSc07z72Wr
KMDezu5ohtSwcyhzoDa3s0yoHsrZpnVsGDVqMzOvu89vl/iyZgxLLziwiiYAMY9gG4AzS9uFzMsY
JzVltSeCvg7w0ajFr9pyrNm8zspvBOk8g0HnAc2AC9reJM5nvpuwYudqKAgsg7k6ECg5ev/tuTm/
9xrgKXdamFPsk60rxJ6Del529zisVUTHASvpPXuBbfkhAgKEUb5yh0flevMH4zeYPom5LlGXMtAY
w2iyb8xF6bkbsQja/DT9SxTBg0bpjq4FXynqapKK/dlS4M2iHTqCMaZJeCdp+RcFE6UijkNAx62Q
Jb/F2H+dmIv/El2vXDbJpND1RwcoLq2hkQ8PC4G/NB8otqyzTYitKnUt+vyl3NS2vCn5LLO6Xiha
yLDScxO5VmBZq9uIOg07HYmIBpWbYB7RieUbh6XaycIzI9M9i4pHo9m74sHrA4cE/YEIlGOtAYog
aGv+ZuxP/zXZNdavMAiWBl3vHYRaAB8Gta9WY1bBYePewIyAX86H1OuxNQQqbq1+wRQAqfg8ltXP
XbzChqziwuK4vb9pXWmHsEUwF1Fdr+CBWrNtb85dFLbIZGL74Hy3KzD+i6RcrT3hvFLAxwbZedQZ
9PucrApM2yHuRUurmPH0YzoDATN5qtULrcAm03Xzf0TrwhwLOm34oGKpxpskdr100VEEco0TREZ7
vfQLKbiFFfx4zc4BnZ3MrXekqtBwZ2Em4N3n8BK1BqxT9g/O6pvXRtg/lTVg3QpPXJUVSwtxzIcj
S81qH9BDq/6E2FHVTDWCyzcsGuwz0HOOtW13Jy0fZ6yCcDG0Pxl9ioyhXi7+zx39d46BMS6RYDgt
NhSj5Raw7iOXy3q7ezldvconIRhlWRQHlg+TxX7k2G1zAhbw3gFOF65rZhn9a7wP6gmqmG6f9DEd
wRhlqkU7tERl0/0Otkjq0ZTDgzAYp14Ig/i8U9PAbYIPf6Yo5UqQx/pnNYZOWXFm7Swevnaj3Xyj
E9Ia0Y1UyA1hez50iA+6u5r5pu9deQWimUzl59u03MSNuEoabe6Jg8Y9bRZQ3qOU7z5pcGLOsw6m
XpweU9z9Wr2HbR/QqB3BdazKn4tH+uh50Zz9ndyYXHESDRSGaGM13+Lnte8kamqrpcZIOXaPy8A5
N9RbRAmP0DBsYy3fSBXfvmH/7IiOM/N+cA25idgu7bpqv1DiEZksxCkwLqXQrjDw+4tGys+W+jkr
U+ZhTOsry5fZH9cQgRTzHLKs5S9opQYpjRCI2xrKGR/yybfCzCSLhJJ3aBYzZucIPbIGekONXqU/
togRfobeePYPsDl8sCHTXpxJg99ztu5ND+ZXNn+NQIxDGoZsHFIJxOm56dbm+pOsPifTx4Ws1EsR
JeQqcwbgp9oBjjfG2WsmmjdywB/xmfSxng4yMas4ls3LAZT+WbKOCurRdlVJ2nyTq64r6kggGusx
D0ab9JFhxs28vCQMgMdWhH4NHP8Ho8K5V41VVUFg47nhO4lgtV/2wzDBeA/U+WMWDzzuiJaGnq51
6Wl9AGmJt07PIqSfXPXCMbrih5kwY3ntPMfLOeAhQ6PCv7qorMF+LMobVNEIOfIAbzISdv5oI88T
ZP+eorbDO4ufOJWfVWbinYPqECM+KiPY7ZwU+bsOH/4oUVvbMjRyZs/ypfxH8Cc8m4GryIy6deVG
SJBhlm07+WojJ9XCSt7fMmbzec2NJ+LLgyaeU/F5zkSLlzTLTzVbtpS3VeDq+G88w/0gCwum/N6n
II+W3gbMlCPIUwqH+na5xbbje4oxyNjei56bnG2sEhZe9KTt3WSAN4B+/oIjVrYcrbxZwfOVwIP0
P7mZjzsDUcQ/tycCWVmJCsakNyKE69BjgkB8173seXwPDCpngwA1je2cyw/LC2CW4hrV4AqDVvHK
QPkPpXH4VSar9yEZ4fexZ51GbcOBz8bGw5+uOifmDSm0rpkTE331EwzBIaW6NKqq+riaUbeAHKzp
XHyDsHsF24PyyiuQc8e77MkEJqucXhF3LIlFgevebXqZ75rQTz0qtUeInBydBIzPMp0wE+Vm8Asp
sUqydRa2AD/LixfxTLnahd/0qDyQYlUsUq8hLOcQbubP7AMNeX0ffmpBni9Q2B/zdSnYksFEUl+a
Epyu82/XKdxWj039ia6v2Ra0B1HTrXO5FbZyvRNSnnXpRz/RibczJ5DescMEb2Kkf+dlRgnT8hhD
Ux3xZdfvrJppdXIyDG09+gI4UeX/09B2VutCElkxs305xzMxsmYIaeqaAj0ZHJObDNSF5uhOJLaa
XSH5hNPBTHLAQ8ibXUYDG4CtiIHQDrV7fiPYbvEQb8mqqZ/kfOoD8mbpoAwh+MVRI5Q5VSTzHgf5
dUaaIgkbTTZX+Lxc3Dy/ggsam/QD5qC/hsv+pOnzVwXzE/Mm+cYfIxjWkFxkfDthj7WQ/b/T2Fk8
IM5iuzN4aEUodXK5ullsPICeEXNV/ier+/Hrktn60UpKMDiflKi2khweuGFScgbNpncOx3sHul0I
O6sP6D3szipRWuDN4djmuMkPEASEA9R8i3g1RWTFxpXAAhdxRKl4NeScw3n4Hu2XnEoJylhUzIOv
sxvTVBptzwftxrR1v5eUOLUbJM5ISEv/vOGj4pnPa/X7NLHwFwOtrOQqNUYfwfBigt3uQcTJfutz
CKRSlojYB3C+PRP23rtAVoC/22yZPFk7ctnHKYk9/lCcp5vKyY3vT9vyyflBX8O3+XtUlkohKaYu
jc9Rv+WUtEGHiBGVmd2IiAS7U40A0yray8htyyN2QNNpAUooeUa203NnWLmWWV32/2DABJ4sVMes
E6S1nW0Diymo7wz11qUQ5c+9ZMw14Tsfr8/znYIhtaWLnL/ux6nSdQsV1Jih7hGDlSU4/E5rMnSB
05/4Is/B0ilC2mfxO0RcDeYIFBfseg5125JLa5DgKBbWGlo5WXaoETc1ZB7MNYl48vtqushVBg/6
xUJ6Y6GqsG2vLvuIWQsEqULVjwMt3H0W0fWPUo7e+MfXnuKHMlPZYzdBPt7wGjM5O3aAReou3wIn
rbQn3hIh22XewO8lNGu3jM7gRc8avw/LKRC/CH/FnBfZKmxO+Ocj8imSwNrDKI0C3IVg6eBpFawQ
nWDb0r9i3Xsn1z7gUaYsTnHE/EuXXSTaPj3Boca5c5YcPvyhy9Uo55xG9GKM4Mnc5oy9C7MKQplY
99Z6egoa/pXPcylMmlFGt2/DPpxZ/pScnaWWq7iNmzOOC232cojk0z7EYuza1udnpA8tyT7HAsOT
KdkMkt+hG9IrMo7q3xWtFHmvXPc/7yJZn0p11uK4p205TTAkBLK4xgog4TOgKJn/qs9219bMSBL7
RPgRoxDavj5HAO9knkH4DP4j1OR8hZo6973qNDWIuMZ4QsfFYyQxzUx8K5GNFQ3Znjy7+Gh31S8b
q7qbZm2DeTOcQcQJ/1eXqENXez2kwsXcqMawjPsaUC/IdOOsOXp9Qm/RwQiAjps4f/2f+uvceabj
os7QoJqop1Ptn/mh2mFEpJRJwZIYZUdL37kgZQto6Fsqc6eCHs589vXAr2dIyLLoOVf8t9i5i81S
kdyJtMnJhSh0E3uhpRtNiCTwv7UHnBs8iFpPxXaLi2sge9G5E2PX3s48g6LFWLgnPv8+ZczHxUVg
3fGhPCEpH0Rg0jovTKOv1bwUtdUUORKQhno0BJiNvvibYRVT6XjKDNW1pzQb1ih1QzGOEnc4fku+
2z8T93w/XVSZmsCDeqiqVbaIsHASEiD/XrEFgtF26mhADi19439XSiM3moVXzvB6LY+8NsZS/iiA
Y2jebFT7/wsVUYnstEaCiCZpZ5KmJOoAhyrNiiltj3XdOmmVecnHgzQm83/TMPChs86XswLKg2ij
nXqzeRzwo1k+VvQBjjKY3pqZf7GRQfikIo+5ChXjWzuDuWYv/lwXoUPPjScOWs3Jwaa5vkD4Uzho
GkT4922gM8Q+mmifKDHI+0i65jsnkPpVEXX0Gldh03W7Z7Ma4HB0KkPEMQfkZHKJP7MmHuQ15XQ3
Q9BVjJ286JxTS4kQq0Wq0DlTQ7me3Rbzn68tHgBl6eTVNEB3z54fjgCwTC//jq6ZrPDsAttvc6CM
VacTG8W4JeAkk3ytQPRgQ+LSk9gSKnd22EO3eCwQtAKqKtq88H2BABIhiQ9uVqGtzgH5qp7DJdXe
RQ8SRMQ6owJi3J8Fn5uOk6+PheBjcAMmRVt0Cqosjq53S7nP3Kjvnm3jNaKVV0IbgPtzqtKApcGi
E1wKn0qjvcq25W/EtUL7/MisqjSdHHjnqz7+MDp3nagyLe9psFLP3FWL3P356CcHCgjzbYXS+Nie
4liX5L2QK3Avq+4PxIPUfmBc/VhQzRgXDLJ7sb+C5R/w8kFybP4kKr6UaUqtnQsi5taVw8aXlUHK
vBU2SddG2b+69PsOdr7b6RqiL9gpYCOImb8xgiRR/82fAAhQmCi+ZUnE5rmTAMup2oBLlAgkVp8V
PHknGbN4q791paDgtulwtsR8MGj0iU4EkOM8cAyw90JbtTm//7CpO0ZaUv8u7n9ZAiLHUQO2ubwh
1TC3I7lDYZtBwMV8vmscmDPJch0/eg039X5H/TCAcwqUsOJRaFyhum+ZL/5CQek8aoosnBAMgdjL
ivP72AxnW7VEwAQw9CNL14c7Gwtbrqix6dlwcvaK00CUH/lV58k05tJ1K4bnD4tq67XxTiRE24TS
q7OpZz2z4biA6rI3BrOhTci12agdwbTGMigbb8NyTPDDEsyo2F0RejQt0Xv79WAI61De2Yx5MB6t
sYgNE5L8kgVCTb1j1pBTQngDF5OyzpHj0bXOyVPeqvreA4g0a50YxvWk+LTACafwkM3uKgJGLfLF
XM/4otJNxY730wV6OXFfrBzmglnCjM1azN54I+Ox2RkCsqmva01fy1vgww8IHjIB+j/wWkgmiJZP
65LzsixvKnSMDzmoDSw8UAhCHH+Pmru0aj7K16RAFSv97s4ZOaWMtioCJWL7f3ttVDegsOUdkXLP
t4/sVky7Ja0vguc03xc059p+xePBc4DK+5PHCyGmYTc9V8a81yoF0/3b1653Q2Y3Zg/W3VtoX5Jb
w7TZtOE7WzOAmceMBlvMNVr4pQjzmnMIyqqKp/q/KzRBV9Zt56x2s204BgH45SPH7yIJGuAgzrqI
ULT7Rb5FHRTM+AKvnF1pZamAG/ID7NOBdyZdCqD9h1Y7FJVU7FTOUb4lIDpMdQeMQGmDLLamorG+
sxPdFth8zZxTVQV7W8CnW2D/qg8eq/9SIP41Znflf3AWn7P/tVhvyBp+kDe4JCg0DVktNt413Un6
rr6uyybx7yNU0B7QH/3hJRvt1lqkYqYMFFh7htIVmpGjMum/IJ34HcOa5taZzm0ubDrqYOcksYUX
MHkeTCQo+e/7lS4dVtCUPBhFoicnybJ/GQDc3QTAV9/2z12odef0RTgzcoUDJ10PyosALldRiT+I
SpATsxwRh0muXultc3F7lyoD+xS2ZeadsVbVrLcpT9PwC/iVVymaWnKXk0wplLDfbt3lk07xbGMi
nrB69rlISDWaHfJ5tLVKYsxeICoD+BmKNK9DervvOGPg3S/YnmBVyVB97JFm1W0oVuQWP6ztQHjP
3zJ60JfTwIga4IKvS3n5TvtEAgZrDVFbxg3PBUFSMo6Zw06KFZn90N8Mp4N4vidm4pC3hVmTaYSx
x7GbaJB60FtZ+030cjN3mEJNWv68yAPpO2Xjsw9qVd4agA9KGSoh64v5vy4egUP21rnKXcfA0c8d
SHa2tNSAG9k1s/dXt2MrxrR0TWxyG7SLl6vZXD9wJSz2Lwb8UufHB+4BEqv7BXimY/wyqtdNIEog
T5l20os8dq5yFc75f3U+CoBdhHE3QaIJ+/CQsQGsVv07Fe0hPoWWLpyV2beEIDQ308jKUP8t/GON
8kMzJPtCArhcDueCUr5S/lmP8RMsE6U9++81cRhDU/JMKb7N60rOaJ7/fZnNjIKd4IJeaxu7//+I
9SDck/3cKPq1mQyUL6Aa3YwSblWM3Qb9lf+KYk8sXK+n2Q/nRboAE7mQGSmxgM0VFaT6y2dF9bZk
7u3cnMLiIZXu34vDtyEL6yxBeuFnW+edSxY26HAHwC2HB6qNzfycYIhFA2vxAWGBFMEPP73LJL3D
MVBmzplV53dwaLw5GmeTYWdWSZgbUFeNtc5ZiJK+G4xWXfMIpeEuzZcLZPQOYfHqPW7zU/zEcQ4z
mMFT2O3tojAYN2PcwqYMupP+IwwmGw1679oEegzHFG2HBmjxP6+OOXxa0qXCyCm7t+5GSItuhfCq
DHoM0yCLEbA5wmBUn5C0Dp1wZV0erurLJU88DksZ9+MTdjUv0uc8DLD1pTI5TbTLOXyzvfQP6Hu2
7q4ZAwy0cOTJQ3E1NUxTbd/dLzOi8nip4PMpuRxa06G20Grp/QKmDP1v6O7fCH3RVIZbMJU3/SO5
yRA2tTteGDjxmANMvEdhoXPY7YtZ5ZlIqKENkiy5EaV9Eb6yFnpNIiT74Khhu94ofwo0DXMSdpxu
8+X4jHSViLrgGhhoojcZ84DJgi/Ny+LPteyRLMWl1SYu6H3ABDzB2mCE+Z4DYPubjsC3g44DWrDM
WjXVdoXxWer3DaErzNJ+hAtQf+pxOj0UX6sTStL7d96k6JMCRpQy5Tpo/dkzaqGbLg7PbD4vl7Zl
uqthCn7fiV0CnBSl16bitJAXCSbWOoCqeAaI1KtYhQXdhtNOWoqXL+PjSB/OdNwfvmXdThP1dohg
M4bXBA7eQ7qfc/D+A9/2nKmj4I6MnTAA5iDSFEiWti/UAyaaybXQeOmCq2ghRxMWKsPH59i5QtBD
5NCck8+7CpYp/G66FqIVHNxNde/ZHzSgOY8z4JUXdK9Fj7FLk3I4vNHV87wougmANHkIrH78FeY6
fv55Yc7fgGDxE148ixYCs2+r+YQ6AP3MUn1lvktkSpxP9Wlfmrbi3RladSXWyzRCRwOHma3Ed+Om
bNI8fkHbzNFahfBItm9Apjd2IQNrOhU5sRSkGtY/lvf7piv/J7t9hwje4UQaYNdNiXTbHV5FkAQ8
ag1zXcZ/clUK+hHZjbyJemsXcZqltjyhTP47acP30Jmy+4hA6dlbn+o6nV3/A/Hx/hp8TPAOicKT
y308DXB7qwKjY7IsK/LieSjFZHwTO5xZNfcc0dNm/nloqYhPiJKdsG2z4v1cu7GK/6Hpk3Zbf6Me
ZbcTjOQBnOty/Fqw4XLKzELJ/GVq7Bq5DTWpEv3nKEFUE7UorzwpytM5C10Eph1be9z0J/0oh7h4
zjRgI/qKoPNKuiPUl9rG37rC+q+I7BMXNk3xLYmU6TjSLvq/F4d8wcXJT+ziGj/tdwXucJOUx8ti
x2a/aB1oHoCYamapl4bzMacSJlWzISlj7nEf7jIgpJ8ozQPDRSI4JBbI3GWHKHgPpGBsX9zitf6+
x0scSigwoUSlaIh4qRUwhucu+kNadoEUzs9LA1biBVpNeEUUFUmXIkpio60My7a5kGxUTmNKmuyH
wpe9WwjLN+tyg/WaB7Ecxo/lvC7RyQ9t2CmBoBunxmgCEFxwZaWy9BtcAWwPfhgdwYSPpnfHsT3Z
wTiLXyXmrG8ITGmtQUgyxu2AbzxfftmXnkDbJyfRMDtkZDtkri5aOry26O1nA3Ov3KEQUKYQI++t
ZVkBVfIIHXCCwaeEBCAZ4poPjTS0lIBE5dorZ3E3tSDNrTZs0RidVn9sS1uh88ndS9hXXWFdYC2E
hhRUTl3rRwnFGveVjDXlcNcE0KPebIIi5ptEzhChwnXvNNpeDhwdMgGaIKnEDh++U89XMYgPtFL+
KcMRQcGfOjqs4yYQGMVRk3hyuDMnuXYlNvIo/hkjZ80qflqyZRIq3kkybYj/vqKDBBD+ysQmMvRC
kcUvdbgjIFsfWBJI1ZWEZv2O2dJLcWXIhUaDRTCKt6siVDxU+h0jb9sqkPL16PFpuTTj7qmGorje
S0xoKoiZlEyvH+m4yqjlyuq/rSx2zNG9YkI8zsbLX81MHtX+N13fdoZ3ijRgNmJ/16bvqXBE5tW/
bnX+/vshFW7icU1YuKT5FM7fs1Dffl1bYw/YGPRJNJHI/lOS2YDPfnCBKuMsgZxhNXd0XySTv998
ToWFCrjkXxMQUjdjzlbdFMSzd5p9Z6u3hodUdxhRzuD6osKxF0PtQOgKGIqAaYHOuA3+9TXvbUqZ
D2021hzqdjjks3rRvR/vVtjgSjGxirwMk4QOTS2WVEMaArjCACrhiCiO5c1OzEX6A1Ugsn3iBe13
hfo0eflRtjbRrauH7w/Xz3g5SFbUupwhn+Kb4zFr/hxJ7IjFanjfGY0Kf6qogaBrf3rVZPH4uR62
vSDFkuFY6bfSgKpnlM3HTgDS3HFHhsnNqdRXH1qzMAvCsKeKPgbQ5q+nl1UcEFQvV4bwuFK3Lw65
DGiHyXW6eDiiQFuIkXX8RzuuWPhWLn4KNtkhNq03RFRMbC3gAxjdxWDrSJLtqmRl/3kBNt2bD9Jf
hY9++DmhpPkLFHIVEzZD3szWwDPdTeMcp5o0EU8RjRKeXYmujAUAyWcaGpwADbKxDDLlV51iWNBv
EEuBF5m15YUBtXIGfL529HldFUeeV49lERNv5Y75K3U+1vyhgBDXgfSqMKJDrLwCbHEnfPXjPevG
Z81yjcQT+13mnGlkCuS/jXm5Ex41hi8FxlmR2rK+42RTR6wWJbiCrfXhznzrnDuSEGk7NngbCknD
eCMMmFPlFtP0760NrXNYhhoT/jULt2owY+FOkRmcRPJg5MpxyN6zcDyiLfsKq9BtQw8pO4cqqxI6
STgqIHHY1I6KTaelopfOx52RNIJpg2aihv+eZ9DiiaUjO3+efnouXFyfLkp93GRhkgX1x+EtlSpl
ww4IxUFwGReKPPHDOqGKRlygNMpffX18rnkmXE0XeR7us3HU+E/IpOziO/8wv+xlXpn0g73QeCv/
3ytfj8Lv8o9p7cooy/AKk5GNIySnHodU49zpJV6pG/UgDVngFmkU/4unAN4wBQft9Csbl+LFk3q1
Tfb0eiAURJOcs6ACBSskmRh4hjEkRYcpOSREvbr5EfZfrlWiLkfn+KMPx5j6KEDeQHCay13ikL5k
AaQUmjU8MsrHenWPh8orpGKuIsuK6DgOMua7HielyDs7VLYFsZ1NzPd5Q1VrR5qv4KPYgSCIp2t7
ZEN7BqQAj4PzOUbcI5+XgOvNrvhnD9aOdHWKXIEYa66tRC3XDer4VvC+HbX/fKVRelw8tVpv4LuI
WQe9pFIn8DtIvUYbzmEODkoWCTb7xj6++xsfI5DhAj2/rPKadKBFloQVTRNdoQmSSEjvkNRpUJwp
S67v8eOwBjS3k7+q5PHI/xL2CHDED4Ta6b+HWoDGnJgFqZFWdAZbVyahsJhXf5FyVvqm47Fo2nv3
dyNgkY6ZsBPOYZYv68tvrO6TxQvuV2b8dsinwAn82JvamZqSwnyk1kAydD5RxD1Sl0J1ea9VbJiJ
aBUHNEqSoOMEMJ5dglaV0N5FY3Lx9ZhtPXAZ5NiB0HzeTdLhRgYtdHYc8FiJwhmEabLdKxmIdEj1
CnfVWhykC8mg6h8Oq1K/EGU/OyzxnbuTDbZ+YR15Tzo/n7BWq2ICLHN31AObAwAfHg21Y59x7gYK
sXBwxfHRgOc0pxGBBMjEdouWRoWA4xUHU4Gda36XJGtIgyExAB/ekMs6JDlszpswQaoq5HemWddO
pk8zoHtsCd5OBupNUEzMeOTrNGiFVCLYkCQn/Nx2/Og/eYzVtBKiYMZ+mvxQ1yP46m7/8fnkKozw
x4XE5Mrj0Ef7nq+7QEAXWASmJfEkakt/0B1smhuTQM2MJS7xM2VyP/ZgpdD0IkvZr3VhNRJLYOZE
xsba7i+Y2GFBRh2DTarOOOQak8Wz0CS6F2UpFC9aZ/+qwZBx3BTiU7VZBFzaj92ua5pYy9td0AYf
SkfivarIqlr+FRHzWJtN6QxMQTCP/yXu/KdjndUa0INIEg4RGaa0uz/zRz3PW79ueh0Fkw22WGOT
ybTiIpp+jxaXoXTC3Jonnd/YNqK8htYRvDaJ1vNyeSQzc400UTlH0Om7iZRAbeIZs0pEO5kiHdID
7Ymwpr5zMo58azfUxlrsKHeQFQAzmDCKeuFGTZ1ceUfXPpF0c0Fij67VBvKbfZl2qZGxkLTsiBhS
1wY8gL20+dWaSn2GiBnIZ14vtwVfgkdPHpPZvwpKd5F3DmOQdwnG/ZTauFqETsQX+jtEzm5E3X/o
q23uye49/8KTIcmCL4P4zaDIVprXeYL6pgY9DCnN+9Ljut3Wa2P+9fmGGAPop8vcWn3p1GrzziyN
c//2hdepgOEnftAqtF5GDAydXgZE813bmuhcSzKw6uD3vxoo2gqdMPYENtc0Lqu99Il4jxlqg58x
6DR7Gk1MIfaUy641Ud/L1KtmxQ37w60o2g7g6IGQhsOwsNZLPYKjtp7ghMLenHNFjQDfYssM+Ucf
rPLwd/qdBaxQgoXV0mTGT2QYj8wF76z1fCFXn32lxXxKn/sIjAtG/FPBVnhIn/mnmOx2on/CCHEF
hvUfX9zg8J5Sr0H8J83qrxb+dm0AzK9vpiIxT2TG1T68LJJ++BooVfypQISkoh21ZyROeASH92Kz
DiMXwMnGzH4tMoGGivhBnkA4PY3H3L26q4uEte7uKLuK7NRz65leZBpkM+wh+G+W1iXwu27jYkr2
j7hlNWV3/8jKaPU3+u8XrzwrRhZ+bfSSrfsqssSEOwPbGz6WzMEivWCEDvi4un12Ay9kQ0J/IoEM
CGe7BBpeSLMpxIiyaOgySkB+l25fos9n4PF2o3dj97YOqExPmAWP/2Ey8oXIzOqqS2JlPf9BRBi6
Upyods9rYuVbaPlETbKjKZwqH1qyQZpg27X9kR28Pipqzpij4/TPq+amGISkLiYdnYSHXMO8nhb4
SLd0GNzzvn8giaF87IcaBsnzm814fA7zHVBgI9GJInYqGhMHn6ohHvCKz4qlLXCr1U8mSCY9fdrW
2r6ucx4OZgHio0eTCqLx8+0qAuRna+CCpGkBNLP0DNMiU40cMPZYb3I3PD/ZYnROOVq3MOthHVxc
iaKomcCNeH8TSazZUPiQ3hFOGjJqTiXiVAYtuojUl9qHnCuffmpj5TBBaTzlShMFTNp0tgLa18vF
7Dd3AhGv5hqM9uHHZPeSgj2uXfPEJo/ELLBrucFp+WUMvkkbNs8e9VITC+qsmB7TJgTWvFvz3tZa
aA23nWj3sKnQb9DFx8UsD+pMTzzEeTFoXkvqO3J+E0rwZoSsGUAFP2+iv/vuOiiZrxmbOlmS+06l
ozFDyZlLecktohXh+59zxA/fEXXHzDGB5kd1Bd9/UTe8W1jRYoQ6dhFOmpbRMBAj52JW9k973Fmk
pOJWzMW9S8m0YJImYxIoHTuBvIOFksskUQX1q036CpZLqImej9F07N+RJpIfrYf9YV7NRoDI2aKb
tsTIIyGMecT3ywWhcRynwDmkNajGkr5XMruLyIzoum6MIsMFPbWz0H6//rwoHjlgOvo4Srm823zN
Q48y/BWNCOIjwnYjkwyANpxRlBPKKYxWWXgdoM6Efn4YDImPukLbWbYBP2sUHerJfNOUHqkJ+EPj
eT4yq/jG9xLfRyrxgpUKBsS0/3yPyM7EQklVQYQZgi7wDkD0R8oclxUT9nyuREO/2iUmhpiez/4q
H46QeYMKhgGGoCosperiPD2qjwKPQg1heUnX0ANt5S2VZlWvhV4f7KlGzog1vhOXie5TpKIU9NUn
wSkTl/a7cC9VhNb9LB67mTp/KkrjFfu9FCE1XLRCq/+6CFF2Xs/U3tAe3zPgvskE/PzmEiJV87Ao
TGEOnaMFlMhbL0SSHsJGctmV30zReU5C5ImmKHt/0zdk/K69K2kk8OCW5dVZu4Kl02FyezJzrkVO
iQDQmn70l7oY0PYa0hi/R/sivxGiH9KwQp1U+JbB6IBKrOVAYYu5CsXfshzckZpBukeNs9ZqkoYi
FrHzORvASe574MwD883UGYmx7kDoCOqpkhhXVeHfRtsxJbo4kjtZ5GUIQotFPk0gJbXI0szwJaJk
LNeHYITkVt/h9sMOgcOFLZ66kfBa5udlfvPrkPLUGeu6qiw44T/cLO3ehTynnrl0e0obPi3oyRrQ
ycyE5jK/pcQ+pkMHFEeTJLrO7jv95bePJjfrH68Rg4TWzu0lbsCJ5zI7iTMmH/1eXycIlgjTwhWH
E7Ckv6soloZI9LibV3pt80CJrojywE+Qqwvs6gEsZvbX7bHJeVymDDc7nSxHHNoLYKF5wn3tb1xR
abvWwDyYK2XlJRNjSpDs1O2n879mvzolVU6fd2ilSksd7PD1jqA/yJBX1su9MPMWR9y10WGsOgPZ
w6PKntDfdsUnt1J8RU2zTICka6kBKDi7MkcSEZbam4El2mf0P228UAug4bB1EiBF5zAgxGAJDaqZ
5JZwSouIoOJLPEiLlyNl5oDMMwSQ00v0AUogylSlvaLqy3VkWInNXZXCVdpNQqdajqJZc4sjeGhp
FqZmVW0aoESymezdD/o85/6G7jzuLmcyMvBrwIa/0NY0/czx0sbO3aiRCYTo3AgzZbE6mr4/+H2/
bfZwXVdKFsVQTk+vYaB5RICo/VsUJaVniCTtuCBe6PTHFB3UXZxs1Fh9hba7gpi8EcCaI1Eqljv1
U5Kh3oHczTBXchnRYboSCe9MpU5EIlmBnq/Ot9TG/CL6x6xZdP0JuLAV3FaPzN5eEdyHLb7bogGv
xfCfMutTiUiybECadJBRTzFcipsk1dxF2mAsfnwaU5RTI2MH9K8fLCA5nbW1IunUj1cCDRlz5Ah6
Ol7KAlTB+d1c9LIfvLe6ZHF11KID+kdYJ5BadCHoddMWlM2i+LCAOy+Up2A7Z10tv6eSa+XBTnvD
YEc4Dx7zdv36X+69u1lyQd/Anux9CZI0NO6Y6ViS48Zh1RGzBRqgZaWVAg4UUOJ7BuJcq28jdU9k
cO2ALCRRn45kDvD9RZnE275wRyJxghBlRemOYitbAdnwLi8ZTEtoIJ5XpDheEam6v+EOhpWEGxEJ
p914II8NNtGJgiQJzY/9Mt0evCiNg16vluiMPA+L7v/pssank0+9cm83wQwSVsFOgLWwa27EP8Zh
j5kjFMybaK1DPomVkkKWVnvlZUOSdQwSe9GNwIECxT7ErEyyzarDSmIHtAHlyFWGDj4sdIUr5VoI
CNfrS8WafBIvKLUPIdlXosY01NEoPLS6oDafIXdrHjfpdoM/oo+jVG2KG+nEYato6lZbzCNu+Yjp
EQulHBm75DyMJW6k8zgIGmbaxv5tlGmAegJEHAqjkbCh7JHeNvvF4lGn6WWhvVkPl7R8tK/H6LA7
OSkq7ltbLTqKPPVFUDUThAQPaJLJGMoCFWKjQvr0koYOVu6ywJ/QAcKl4kaStaXQ3YYmNBDwlaeh
eeTdZE0aHssgm0wTlfoxg2Ocjo8gwO2KOTgWUMmnhbKtwsrdb3MfxZqi7xuQb2OiAAWc384eMLiX
W1b+YQF6MbOU5VM5CkujHK1NsW6hjtunoFVjHMUrrt+ZFkaaoIY1GhVwllL3Ke4rRJJjnK0Z9+bB
zGNeNHLOaP3pKggSQdhwFljkU1yMXJ9Z5cqfeLbkHd6llut6fy3pnUr+t4V+taTzBWHncWDztJPq
Ur+584ANHr2IEp4lok5GWm2xbiw1o95Y6RlHhhREnmfZza14hlp8uy9MNaumLQ0nACJFZb7uHDzY
ENXWKImkbf8uhNNRM71UGHo1VUoOaMP2RdY1V7QgE2xKX0hWdrNoa4mBDnprR3fjrJG4iN9ljV34
FXTy/TwffrEDA2OanHqqRIahi5CY/3bDIewvxvjKWE8J5fEabYVohoRryvt3IlsvnR6s3213F1Tw
1ocihUlHiDIFFUrB4xF6Bh3y/TBOpIfyWJZ6MJbh4i0OHFZV2WB+fh/NiXbMkPb2ZqVAoHUjIIpv
Rkpd/M3YNKpfL9UAmMiz/SctbqtkNrRmmm0RGORjIgbexOAPBGid1+iEfgdc702bQX/IILQnOxKE
iBQGoFQzKmoMN/tTt2+UeYDeTzf0vNL9DYmNAeQFeGazol20dO87MQiADDtpGvBq09t4tgNvSQ0w
2//tPQ1YoG2F2MxjuhDPgFdFcTfXr1d1KbTEV26LsyojVUbYsWsNqv7N/IJhpLsz71VLunKT6RGC
jlThjpUPi/Yx39DJ6CqO/BRcBV55507NQSeeg+A82HVnpytMfA/6wegrK/g8bLtWKboN8UMdtrtE
wz+/FrP3w3qGSASPaWNxVQ2Ynxb0uL98Cb5QqTlmGRkDXBRufM+L+lEwqARo77CrxobGrIN4PDYB
CZhxrAui0LZgqNvcOM4s9oZrTOIhOLWkgKPH/CoQJhHdA6ZowZQcvyc5K37308Tys8DsnbPshq/3
q/RF0Cmv4Vt2vXRX8LrUPCKNg2ZjLfcDqVcO9cstD8YQjYTJbB6VfI1gFc5TOdtBfh7bjGbiu47l
CYqpjmH1iPp8evMDyPCCkuEZ35A4L1rhNQ94Xmcr7Wlb+k7glwmInDvz4CIJWoqTkapYmu0xvB3x
Wz67ic90iu54CgA0tAVToWq50ePpUi4zNhq8VWAmcuNy0ZQ9eDrrS06ztKhztAhMOQAedP93bbBS
2/l0fypYqvFIbX27S6kvHx6u8mxmiUAXe8jhjQCvFaEtkLohTsHE6RHGr0Bv8XyUpL+76QKXIBct
3rjHwjhuxqSBbbQXdLHNktELmF5qxXUdoM6Yd20k6TR9ER/az8wtmwtbpYL+Aa1gWiyqhnOpjSOF
3Ymk95C19SOfvrMN7F2yqToN3l401FT9nBDmefuJFZXR+8ctFH4K4aHvj8nmNCrmJnjSdk5JiTr3
E3xET4UaSSvGOHB5Ii1NdtxNyKx1ssu/GHH4g2UFld1zlsKifcyexTkiMenum0/ekQTvHM6eYQ5X
YgWixSVtjtOaQmexbKWI7IMCCMDuoLDSmQWtKvNGjcT7KSqjSZpp08G6QXcF18q9IUbAwOeKkREn
U10p9nMNE/EpiRJsse3cENqV72MNvx56OGQm6fmdX6KQqn0ouuJx9pvBlBqr2yQ2leY0x0+/30k4
/gYzwdvONRT1Di7Q6KGsajK+g93BRSr+zf3jotQFC1DPu/lmNV2RmgSW1IppzEs+EVypEOAhoQsq
w0W/DR9ICMjXC3fJV/35Ph5hrNGnW2K4fPazX7iv/+4WtJkaW8R2pg3+hDK662I5tSjnQnEwRfhV
y7kRORAr0oQSjuk6+pp5uo2/wQd+9Ziv4mVEKfVlXgKS3gLoRjX4WBdXfOVFFoHemNr5k2jXDj+x
BhPG0LRJ/4aTr39iOPxBKYc3xFqXtJprR0RtTY0J4sm1lecUBpXszyVYOEnxLEfbqgBZUP+u8Zk0
IeD/IkQu6ok7znz+EDgn8Zi09Uk8D/ht+8fohPGiMVkePGNXYKCJHIz6hdzYbyJr99F8xgsFfg55
djsW/FkPAvkqONNp7E8Wl63WC8kZi4pLOTvebE81q4whhX632CZQIEDjXkNTjCFdeQ9E0tilSkka
iYWMXj0HWa7pQS3IfUj9RLTPIxyXpQLuUvscsrzM6bIidOopo60furGdyp4xPrclEQ4SQOXsvPo6
NVEomY1Igoo7ClRFpLZ5LEf9Q6QeJ4hCWdfx7Y7A9hxtBCLZeMCa4+JlGn0lgi2047icv8DW0lHL
rC8xmKdZUhPiQuNvEnAPa0vnb7AaBDcu6jrhBKxfdWRjKfWY8KgV/Ppkt4G0Upz4us6TdVu74jk+
uPjA+ItnlccdMJE+GFcjcRQWHkLMwJUCiSHo/A99NmFb81RcAglcQKrhdMpFZcekutwhfaQNbJs2
wQXlr4iKL2kfjkC0W3RajPOnkOMY5/iBVAAzq4v6jdsKxhEZ+G70OR9cdcXWC2GtpumJvbUSKxKd
ta0AJvzxI+f3HmvPgtWwmyF2VToWgUJPqf5arDz+muxx5P3C1eGlEmfS91jKfQPdyH6r+sZ0VI17
P5FQw0GyWewpXZGWsMrlNIFX08EQhw4kb39trADbbdaePV/z080jnBul6q+oHoVwfL/P0uAqkN0M
xCqK8VgpqF4lN8dRzlf1Xdo6nbqrQCE+tyy40TEOgojRT59dXXjxftnGAxGAmHXj3TycB6m6ErsW
KvNoGkfKigAqxejhgRaWwX9o7kq5NX9AWN95X0T3YHi4i6NfeUM3YSWXp1WHciKCqqR0rXfiDyqR
tVyMu8OplpHNbdBHOmqBgkMp3SqQjdBIpGhN52bj+OhvUOvhaX00A78l6geS008tDoPbiIlQ1i5j
bQrTst43KBZvYqMvzECqqd7YY8Fnl/bSiHvzu3d+78kj7HQove9DbtEmH9n7r+FD26mgp/rnG8RX
dGyU0zqF+aqtpH6srkkcF+xVlaVADyE2pKF/ncH5oI4TJi0CboeWyqRvcNo+xQDeu+XtdQq2piN6
H1+Qxl0zl4K2/vJC7lYxoXBUdzAMM7qhjTzAAqBotNoiLzIgPZkAUwV/jUXwkOrU2QNbKrWIslex
du1hVp4uMwxzFZiq4gqfrk2wOqzEFKdsAC3TWZ6Z5/dchvA5y2Q4VkxoUqDuaAFFo4cRdNMvr8mo
YDg6nbDGz4C9YHesUuSwoz4bbq0iaiTSNrRkZ1066Rd5suSqMxjTeVvsEbDm5N9f3BtK2x408LU5
yZ5afI0rVhQuDrNM2g6psmDDC0NokywrFAd5NNp3EVceZFCyfl1Vwue3DMpd6hFcjaxQ2eAh7k/2
+YoWEKNacyMat7GeuOejGaWZIvECfrYprRcLvwwwyCdgyHhVCky3IFgJ3o/MO/QwJmf1RVvNS8Sg
MJv58ABK5FELwivZteFA1i6BHyBDfDQZuMsGZhXnH7itq4seoXYdKQfb15/QFTBSotUfwAK4GrjA
ZNKmU2SJquZ7WhnSqNPAItJ+KHxInVVQErY6T3wDUUfneL4ynkHQjLxgP6/A0+pTHLLL2AiXkZly
Y80+adqK76DB9rS9/o8i2uNl+sjhIal+JOlvhmtiQoHkLul2FrC/GuyH4Na6ISDqksqznRqOflzG
BC/eLbRwDme7UJZ/7tOxakj/+p6YoZTawZreWmbNDNI/NolHs0Wj+o2C71CNNQuRNS8gN/LbxTws
/R3m57i/T0qMOU/G3agJJ2Q5jWeyj7iScKmfsOul8d1hNIn7u/WfBvr3MVtAB3ErqfdIS8omWAL0
x6swIJ6N58s2Dcxn1nOKHABH8HwgcuKMscXbT4mmjx+U3yUhUkw2yRpN8c7C5W7Q5NQPZApTfhR0
Fy5ZLQe8+y2BNyui5l1iUcellgyTJ44ClEXxg/aSJ9Xcuw/9rFgqT0j3MwuXxaw2BJ1M02qA6VLh
w4/C03uVNm3Mm9Cqu960l4g6BHlfpumsFDdMnyjC5nhgGrRofqJXCR7sGlsd3NuXX70IH6wTqVR8
X+/k7JJtyPGCsjOYceRvx2JHUpa6ILVLoSnU0ld5rGxI/u6DqnHXIE14oyLESLqpM+e2qKRa75W1
VNWepN9aq6T61EhSs9SFkjj6BhDSWSnP3bBb2Q1GFzLjIpORT1YvhfxOZ5TqFogndrWB/f5yCIgj
rURNwxTbaf3Wjy4BnfpPKNd3w4oTPzQLNwBxQRR1vH6N54AlES0+EykPnstCMSSUm66RU9Swuj1D
1GAYHUpOUzsBK7S1dtH4AOcgDcOxzUGb77mxYbzD89OOes5PjZvbpt1jnsWTquESnjpvsihvRiOU
Cn7cHMgsazs0znYHepUIJ1e/wIVsIxPru8HX+CrJOZXJHtuC2yxexCkDkumc0mfMCvQRAMuXaiLv
BqVosV5XAlBWxyes4DKwOtmJvIpPpOvPS/zZoGcnr9OphLLnMalzFkesY1Y2MS3sv7jp77xX2NhV
eU9ss69xbxcpW9ZL+8JGB5NqxACpUfBk6mf8a92djJqrzN+3uvgX+BOD9mYCGQ/VyxDaJ9trmB43
2rg9affiZyPxnsYgbWqG82JLixZQo/jBBvJd3PBTsBqThNhIy87gnvMYwKN9prpF5qMNtf39/nRY
PJnzvlj/X5SW23kSpg9GG8PEzLzd8X8FTXbZJ1jXIuu1x4pSD3C4HmAOyhyT054QZE6xXx5rYgCL
pfM0xCs147wnJaU7WUMnaMuBEZo/2fAKfRsVl7AtRWz0uHfFYcr2pfxAj6vJ2SKtS7uxQD/oVJOe
0n99BU5PlemoZyxdEyx6ZWVBV5Bkzpdyz7XmZDYDkVFi6HLfZTlYykEoHpeAyfRCldkKr7lEJBo5
sdACGtAK5s4/qWoLlhmsDPNCDBQBV653W6CErCvN8tjRmlzYJkTbCj0d9FjevP/crjaxlzMqzU0q
osmLm9iVjzjeDEPRiqufCzdbTLfGYUuNdf8u98uwfimMACZuM7o51UW71sFoTjBB6ENS3HFeIKgY
6wee/fKbdNqxznt65kuDby3NZr21+Vwk7b6nrXdned0i/jgmx03rCA3ZwbCW8AUpZiPM4m1zBJ/E
xf0pcSnySvAM32TLk0wn/Qd19IExD3y1fmNyc3FukXz2bJgLf7jh6FXMu04frYzB8+rc0r/ICqqI
xOZp575xQLfTGqRdynGilUqtkzahnTNv1WhMKMX/px1AOnD7yZHpuLPFiWDhBHGg3WCe4lPuUXoQ
j3Ak/hUBZwU/G+pxtRz7mD+uwzj70fjBnKwQonjQNxVe41TZXiMsobe2s824hZcNLFxwKq0qflNe
Co6xMNt2GcyeNhAumd4Wtv+pByeUbDYgU7U3otBdMab70B3KIeWJING/JcgxvauxtziCUbBvs0wm
6nl8Sns+xvzGlJj/punuOhM1h1eXyTFFMnvEIPrwrcPYPPstfGXosUHSXgTKPY2UVfFo6uAMclOj
5IXg3LgXtwwO7tfIZ/VjE06rdq6bTqiQXc1Lkwh8YE0/y3EK82eeVKe81v5uGC3KWEA5A4Tobyp3
K6SVHHWQqcs+9A8bZOgE8+hD32CIl6AjnfitqPgt7vLcnxgyGbdy7Z1v8QeomkZsuNoFWKKA2GIA
pW2Ch4fOma5pUZ9/+YSfQhJRQTQi2YEl/ZmrjEBo7444Q14BID1UXIpYFaf7muPZkmBM1lMqkuVC
VhpRTXziw5jCrsoIPVSh73JPwRnNruluQ69il0uFys9iDixYbGey8EPd2XKfqfZG/KoDX7ELqoqE
DAN87qVqc7p0rIibBwNMC1wAdYzg65nJSGgn89ZaNrr4EmsbMEKU/utzxBk8tMklLItmVir4Zfsj
uomZVHbZOBsovqgnQPiSmIzLtrPklH5J1MUD5t6IgUz8jm0BCFjHHoBUj9pj91yiX1eOhQwzSxCD
Q2MrgruvVZOpii6O+2PEohJjzT8ZOT3ouqZtgdlbLFfWvSkM1mEAaBi/Bx86Ds0XPVWNDgwr7igV
+6CEXlX8qnhgZiJEoK1rBHkKkTIM5jFH9Kb6WqJG3nuGbNZoKlxHFN00mIQ4xAzcxax6TEYmTtwd
4mtGV2ak8fDA2ncg7mWJLKGkMdnnGcOsyBWLVS+j/z8wGoRwBybsCdQlsGJ4K5QY9vnP3XILW0dg
gCQ7pTDzLXmrl367AM+wEouvUPLsZlnhtGO2VCBRltc+KrRTFlVUB32bH699EPw5hi+eZvFoRoPw
GdSjmAtqDC75cLErn9SqDIG6AEGSZhEaEvDF7ITvuroONdL9HbV64V3weJRqf6K1jDSWy1B3SlR9
iqz4LPphvKGHWo+WNfAigoSaaznNsR0N0tW0oOjHDBGvzKjSWh20BuNFNz6rNiT1TRrSdAExWKmH
qwsXV+2CFz07l4Jgr7QwFG0qczskqh1d8Hpgg2iNNs+nt6CAuHTd4UyQBTxuWpxsjgzl/cN0zSk9
ZPalADVRJstMdJTftbsmcnc4nZIeUzmip1MSItqn/L54sGJq/lwGxTU7+daDcSDzdf1exmZSHx1m
6q5rMno8jEsWfav8qhSDR/tOjUQBW34pI6jcXVY4152bScTFUNUErb6Lnnv4uJdfUebAZ8y/amB/
zMacN85Yyc0tU2CWhOnUKJOe0rL+nLuo6tALobgjd2vqp4q592uga9VWmANFukdW9o3WrHlzxoRx
gE88z9otOS+WGtWyWZQtO/akYRkoQkRwZgiuXqPvOejpP8y3UfgyZBFES4zq2pp+N1xegVPs3uzS
ndqUaMEZEkVoiSUWlI18MbIB6yUAjyu8dR6CXXllo28A3iHZE1u6/CTkb2yC4KcOh1Ng/noQcpMS
oYUhgcD2K448GS+7LfRMtdwVSElT7YsUhtMz0a1FoJk7GNma5OaQ3UgawtdKmHseA272RMFEXoVG
dklKOTJ3cPcyMHZ+IxG/F7TuNjIh5hQ/2QY/gmYEIbDWsUgyyOk3McfaqsTZfhZpnXrH+YzF7OwI
U9o6iNwfnmKPreXv+ATLXbPGi3NSiwNeG9qiAg5hhC2SF7D5WxGjkG0veXp6fDOTke8o/HajA/jW
jDPpaf81cNTdUz+Fi8Y3d7G/lWyP6Shr2kl38fd8rWl0pKNgUTrbgYc9J6+oDpzzPAGRkC/cXwlL
4rF4vJ0+K16wkL41YwSIVjmvdrv5JX09wE9V6zVEQUMCi5RPl4RGGjURMfmrrYTHbCntcnTKB2gy
Kfb/15MpGVKBskx2bLC2zVq/70F1LSjKsb+wFpSPV/8AXwGQ9B6W5gzL6YqqSmM59hWmmfXaoQto
900X7s96FjQx89zkihegAS8pDjVVr3TLpf4GZ5uqMvpfn73SHVmRl38S7vqgDRbun47HBSTTURLB
cHXlwZ5z4zAzJwV/uPIWqEmSx0p97NIMJVeE2wMgDNDzp8KfE8flaAaDda9RdXCcNRoAZ8lH5rTh
4eA0ksi+MRZv8oLr6Q7xgUn71RZ/62h+FDUV2XJysdfNPR9249nTTt8nkLEV3MJSzDc3YDU7omQA
CqXn7yjsxsFxgf4wxvGxoAJjk3z4GmauV0MPMCcnQHzmdbif2GnKr8QsvtKmHiSHTdjl6YFTLuOR
Ud3E/VaJoBuPLYqwfWZcPp4ZAk9fnV3ij5hN2iExWd68eh6onQod+1nDpBO+VWDO8fNVivO4h6h2
lb38X857sH1+fobZoEIWlVFHU+YdJbNczLYzVw/mVq+qj3aQIDTmjiB0XkEeN7Of7w7+byedNCoL
UQXfnFU4QNynYoquuMeq+Fu7X2EBWEnstMdZVm2azdh1UWY0WqysIwoOeL3395EHQlHH/j22fraI
DCUO4A7ieCVzNCbCi1qkixj40nRlBaOBPG+6nDJ0rpaPFDJwqF59WWS0M/k6QfvNVmnutdjgwa5M
GaG2jAjecf47myqJXPN5avsiga1hxuehxsMdtm4PXiMEIcQ9d8edPPwuz3SmKqGY8pdlUXY+GCd4
Lr3ZnJIqU4lclxpkflpp4I/gJI2Hpkoe110IklJ0bvdZVzOO3fQMLTfiiRVHBJ/4ZlRcuvJlztO5
jgvHXp46cBpGw3Dwz9D/BbwhoAZR9LLzhw954tIjfZ3bRObGTRIRd4Vk4hWtbFE9QoGF7fy8ND+i
1/7s45AdyoY5Kq6sfI4Lj4zcaido3vliQfwJmmwK0RwLbzAOul1Cpmyt2tHXoHnQrN5+QdNZ0yo+
FVMaoeY8v99vgeWDCIDRDIujBnmw/u3Qugk9U6kqD3SIP7mRdFs43e6Y2y2c3eokILKLoK3fQG1z
XE89DAlSnMx9sJqrw9N46/wOaV3QpK2aPIkaAw9lp5XjL/9PF9VYM7kq2rODl1N9zwjdC3m9aLAh
tDjyBnF0YvryeTxQ9eEbB7rc5KzMzPw8mgZITWbKS76U2wr27SsVJ1hh2qN4rV2CIWcr3N8b+iMA
uH7ZC7tZl5Yuv/xYXkS8i7h1SMLm7zxuH3+H8s//bOtlCUAf4oAfjxCfwRkGOc03JmOaNoNcIAg+
f31xNRIvWL55lx8/SQwNEmUle/GoDIbhLZqpx6XSh2tbWWNDCJLzITGiRb2UuZMqT0CbPo6r3J+e
YjhpjZR1fe+IbSJBTA41c9kYCgcqt2oukdXdJwCy3MBJHvRwoBkCOcAIsMBdtcpzAChLeKRDUnqm
BLC3dC+pUq4WI6ULvbjzNdWV+vLFWe52UqFI8qeVUu5aGlqReZxyYLzWf9Ig/y3tkyi+8NeZeBCl
r/oCj2p+LtQejpzWqapwL9+j5qH7TLjirUF86PI+BXXFKk6OQNHQTLOrd9TcUf/VOLFlL0TXvrYg
mONnIieDKL7kCsKd4awkWhE4sRGVGDEWC8PTlCRcQm7Auv3Kj24SqPpKbXRWB9w4lmYgYM6F7r9O
dd6wEkT1XXPesXuJVcpMwBKJfCZumsK0hVEFY3VBe09i2VgWWooIMNux0Wy1cIRZ0n97HsQlIs+/
E9u45HbxLtOOg4gwzZ64JHvmV3bvrkLoOV+8wRI3i/vc2Z5VPmVvOmyFRiYmN5Y2+NnABWVKpi0b
FIhlSx1Qewz3yZxDz1Zrlozcrb++LCQrzY4rXAQ6xh+BW0ST78u9fnaXIwCACBpXoA9Z4tedfKXX
pJpxU1wralDlPGtBCfHW9dNERezSsUnR8cVY2s+Q8gGHR17f2xrxtCo9aE1gHGIVUqSJnEiPebNa
6vMDnhyrBxik8ezSM/oBEeXiHMubBAJacDSACEj3vYOIrSNBZSq0cTZzjkdKP9WJPN245WwTYeNd
ee9ZGur6TdNkb5gkFmmQ9S5E0sXl7sPPRd4Q+AVjRIcPVegMsQ0EhjEPo74GMm/ovUE7Fooz5wf7
zYfQx442/AgIfAcnNMoEGMoJewCW62VG6n1s261cU+jYAxAsWJdKB1l6yE3T00PYns2wFiaMi4c8
l/7Ml8gZSr9t9sUpwHWIQFX2A0QjARPtYoayBBF0I0K3peO+2V8ULYjKoGtVfkdbvJQLaAiYJ3Lf
YwWG1L8xUXyh3tbQrd11HVjm0P2l3zPSk4zoe6VXCrjFgE8qotWbVOQtKtuJg/QD1hqLJ1+1g7vk
Y1cSXj2f7TmSWOdS4mGXGjHHfxVvDbk5DY4Hml55XeCkYwnrltf4eKR6j/YEjHcNvdQMSp1EnCDB
sCvrALrVo7rtlDbQKZErW/u7s639ycyd9Zl6G72VlFeX5PXHYdy+BdbC+k9qJ7GYiIwIqWCcdAjz
1c/2GJHO8SYOVpHFL+ccTFH3O6+byj6ddxK4BNM2N82bJXM83tdJ60o999BBHvu2BaGZxBx8l58w
/pKqNCvI9Nu5nDHg3gqHrVatvjJ9KT6LNoP252PGV/VjEQe/oKg7jubxjxxA2c3W6+ATXwAeamJj
E+UUQpORuSvNKiVK6IjduwVXB+8Vj5G8HCqH33K/q8EFvDDQb66lzoM4Zuu1liVoLK0RfGJ7m7lJ
qd6OK4xh1LYv7N/K9CH5GiDw4qrUwFie/0amJ2l3kWFS/P7vWu77MVph4VA9aqoA1Z78ke3r0btj
4DXIONlnz1FtiZ+EA0uyM90KWHCnLz5DEugdcXzevnQX0AwUlxg91NSI6Xawo3vkn5ByyKySUL+K
QfJ4McPci43d90YJqqSvH1CfR7PathrYPm/HSa5lwAqpLp43YQNIL85/TSOALeaPOVoyd24nEqo+
tKjmzVpyaqmqsn6sqIfT2jPJ2j1ZImjCgDTEv7/RlzmAOyd5c/8aKq7vLbCWbA/cmH9zStQ/CXiL
AdtWGSaIvDAst+sYCaseiWrOdHppNqdqH8dWqOsaA1nZZlp8VoSSpDs5qVSk5DMh0fznynjCI7DA
ip+YpDjR2BbZXuX61ft1QNfyWrXehNyLNAYpMbG07KbOf8MXCKr230hjiZSdVeIOm/pYUPUWzh1z
ZIEGdL0IYHyYEY2eozkb0ht+EfPmzxfuZXRSxkc1RogtJJ18gATyUpvrEg5BBtC+6obxEszh+T68
Cl5/BVVrbl38Y+LUVA4k1tjZof7f90XjSUiWJli1XHJ3/Aqdm0dVFe8pMfdeJMmx7B7JZo5EwPvo
KhtWZwwFjdzQj4V1ysH/eR6XMOTfsXby9OVzS6RMTIUnfB41sUNklywITlrws1dngpb3SXzD/TzT
McWNHEkpaFSh6+P7Iw771drWr1o1dMnQLFcKYgfFi2ZNhmRPJ67PJTU7epbWKmsdXvn1nf4pLJ2A
aKdSfCUw1MoA8jeGrkYqE1apCBEiDfX+y5N1oaEzA+HTNLHCy6QQVsQY2gnaOSCCz72IfERreTE+
TQtViKgSj+jq2xMK5PEW3oP03fx+G4Usdn0VDk34IeD+5UA1wKLWoin8NjXGQLwyccmuDgIdSs4I
IDqECHJUoizcFLLCEYM3MIPFTIWVRKhqRCO2DU21Otn0KQ32TtYujt5LOQfCV3z9Y7Xc9JKB9bSE
PXqYRWN0tlm1OB/jLWdNPsNBm5tnIsif4e0gvQ3L9u2Qd/MVPOPh6fgaNKqhG5wNqXSL7NITFweZ
dMIkKrJtyDzFxXQ01NL28VuZwkS+vwbO+G40HqNfvZ9kikn3xMgEapTxLQWMpCe5FB9WNMRCxiwn
V5xV4pSebt261Ad/ZOFFGBWjOcx8aWiQQH/PK3MuanqVUPtZOz6NVpf+8K86hjDpD0cVhQ+geJpy
LxCZPMP//0r7dp7Gmg0wqHPxaxhipkOCI70Ls7l5ieI5dbIrdtnoLXJM+AIIsggazwx3iV3lE7KZ
2pTAcScf0rCejeFndFJAThB75zpbySI81I1ArmpryNPIcdPu2J4wYP2RDLxAHepqCK5hgjiMi//e
4zimJPbxmVHPLyZLXaOOL2sZnSRT9Wi62tDnVDq9QfkTtkLd3Uikmen2wNC+Wyicyv9qAU8+ttmU
WVgTuWTvoiZxo9Oxv5AVhtFfGu48FLBiYn+dH5ixUK/568uFsIoufKMBmvHYRW0ZNn5xBHpeOKO8
917JQjiHFz32P8laC7BiaNCBpWWC0e+vFEiaNuGN/JdVVqVTdnwnscsJJIrTK8mhg/X02EDrdna5
xhOAJkWspDXjA76PgiBT2BR+YTuZ6hqKogpI3AyxTxkUh8llOG3CkEeEP24ZPOJpu5K0PeSpAj40
4k0vwYLQRVElEMUVNpBTWdVn5WV8Aj+BdDvrBOvEB9JgDBTHQeqGGiAUEbh7CK57QOgQWpC27YgS
z3AwTTsH0cduwzO1leavbN15Ll2lgZYqzaeBRyoT2DP0obTHLj2gOGbTlMHxUcGXgYpWSQEwsPYS
oX5mOTeiqU00+iZ2QsknHv/zORmTnpT8NFQChW4TTHA+UUDu7U1VwJeyjbpSxVAnPCmrFzJ1WpwI
vNt2+fffS5mDtrFBiHrFg6M1hRegvzQ0xCaSaQbWeeWLLvQVhIW8M7yCwbVzjwnsX3ZOAl4E77zd
uq16A6piTmNvF9M9RLqwEWgQctIC+b6EuGaYN5NZM7FnJhGIrAqTNdAP6KcLouLZ0idq95hx+zIr
iRY71xkYjjIfkTBYc5DV4Hqde8642ZVbndeS8YpFAaTO13z6Do6Z4QsjcT0uE4D+j159V9vozaNx
Ygz8zY3zaFhZzNBVrZqacLMlZK7+Aoe8o9oTh2XsdUGuZ1ZaBbGmPBykt/XX2UGh5zhEqiOPmPsd
IgGkAJVn9SYNozuH/kD9yO6EnplTYhSxbU4q+pyH51T8ejCOtUqMpvxZrMbjEymsUv94nieOVtCx
7zYBCPnXwSjHM4YOR649fO6vx+UN/Ev1Iadkokfx09Raj1qeqhSFkiOsOto/rnFnmHuh7rx8xTla
cgT7snW0ZfU6lMlI1C5I7kKc23uGOVwvM3VRN/O5rXtWT62F/9JHiao9sIT+TEhXkP8tcT6CJgIF
lnWWnkB9Im5PUF1M3PUWuKbpewznxJ0tXwSigo30AVq+YmKoQb1rCGmAz6/p8a8I9ThQnu9QiIZi
TABUKm/jpQYL/mGv4DxXa60MijEROEOrYg/eb3Xum2RBpnL8dzeLCg+ndLJ5sCOV3AuB38rKvOGm
lHCTv10SKsHFNJZ0VekhLSEgbWgABPPHag4rssGkN16mL4tRKa1c6qRaB5H3tXYBLuxUfC4dYEdx
rwJUK8T9+ydJzw0aezYKshU1S2SH6SgYbZdnqc/PVZ3rxPOE7JIOO21jJau+G+MdIX0ODeFVyswz
G0bKp3/rq6VUA6VNl+qKgGRzXZx/YQRPq22BDcrrO9h4JWE+3VVfKjlbWp0UAKChG5tK3qMGxXxy
8TfuJPWywSfoJx9D2yCxTIaDpCafPGQdHRJ7eqZGWij/7CkectFkNFm9wDAYWTsOsdodM8TxTprL
yDLxunIzi0iYbqyZdA8fAXLaKBx25TjTgOkiK5UbdR2kD7mRzGCjOZNn6iH/PrnB7VReQ4nK/1QZ
RGAQJlZLuXhDtRzyjko9cbmuiy5UWpJLTXgNmSr936F0v4XjjXXYKRLRbENBlg4ThxCQEv/5YZ8T
KJsTWy7Os9T/zi2yqX/QH+A7r8BaOvb1CeghtI7djboE037htZ9beXHvfubSKj87DdVwx+leADSh
ezDtjNP+ZL1eaBiCbfApv2mskQx1Gu1nZzA3y3uhNQi64SgnwGc/nDMPrM6QuLycdwudNTye8CoX
gjtHEZD5JBSyPpugur0pCAsQHZmQbtsJkQRjqHmXlyYYJAnZFN9YtK6YSMap1nkbfSQI7Fd+H0J+
qzgSR6VpTeNN1dFvChmxYncKXtZJYU8XgyMhwqBlTe+zxFJUr2wG9Exxkbc6NkE1PYqHQRH1Xvy+
ppmp9Btu4CZvyL2z8vAUwBDSSD+JSR742l+QgafQXXolTMgPR+7CaFSI6ndoXU/RhJpUK7VgrZca
lJyjrVGr9OmoWq5lSSmP5N9F4OsVhAN6r/QI2PEGZesNI2maIK74OG4dPYObeqdNTsuro+GlJo1Y
ovts/5EhrYZ6RWQ2JiC0O1KaCKxuisehFMjTHKHCcBX1iHPWvsao8NJ+mS/6tdlmfuyQC/jgOpf3
KJjug3/bSPWrFdmkXClnxSS4ZQAkRdkjptoDlcuJA1mPJWGgPXapt+LIiImouE+U5t7jUWfYXRg8
EsGxNtJJLMP8o7xArRkHIo6VUGLru+pFsRKhHA/1G8vIQzgpHe7zyAhkpsGf0EPPO/Pw1uq5yLHm
2gfPvQLTyGN74vWeFKks7JEYwpRIFjbjYkX+HG7pcyXFuHwvCddONDo3vAcEfbI8M0cy0rxkzyRZ
oILW4x3oGn/fk4gJqmSko40buvnAylpamQBHmmzIuPE6TOIOI5UlKvY9h6nO67wMRyFgP3CT5nRn
cfNvJHoIi2CCM9oOgafEiIeIQdhijDKU43WvLiDFmbxXwnuM3rebIiYpT5EBsHTR+o8uiMgjZxY2
nwFAPfRgPMCRcdf0k5iR/n0P6voJOmazj2zWbrzEgEPusliNWDMcBI5dzxXmhrb1cqcRbdTm87uO
1XJ0pX7uHR0u8AsNZT93GU6CDES2wmzjshUjKjsLSQSEFxJ0FWwRYgPHMbxrhk1i1f4kUtmn2gtn
Qos1MBqQwnYHemXsmn0fVNCyDVhe88iygc8nUEVQ7P2eawDxaAzncR1fd21URb7wwRbwQFTt8qUy
RlhrmNnbnoOMnPoWXkxIK9LmP61PYiK+q4LoC3OO3L6/rwF9vg76i0wOBT7Odz9oLuDZvOuTK1Fy
d9Hyq6+5ryE5ZIWTRl2XVTzcpJbrfZze2/3WySSFM1eHppS+mHngmtDJ91uUTgeqE+i4V1q8hPKD
I9iA/QM+M/4/R6RvyAc473TffipeOuhO94Sb0utXviGF4y3AHpQ2JBuNXyGlOED/Jg7SVUNPgePp
DgqqCrKEjWoVybAYylhIvH2eY9rNYFLTI7+mLXUqh2jcLqXPmN7fYZRRReBPjGt5nfEq8BJcrR74
GKqfg98pEDn8Zy+TZjO7WgVrCxpzUdTulfoZn2HdsW2YR7viCYf+tjMHV0fV7jEUATJqApexgALN
wFKZEae1HlsjJJ3Ng6deXtZJJIJWFGafIsTMVgxmFn3bHfha8JIzoEhqFnu5hxaAx/E/z2agQFW+
zhtxqRZYHsFNW3x6jAmXfWjYeUpEGeaZxAsWivsBcl6EGIz529NhTuDrm1+wRtATE6aDaWMpeua5
nfs7+z1tWPL0oSVDVBIY4oP/OmD569iMKwnEb+8O64F32asP1l3p9qUHzSyMeiWuNqBrpWAj3IEA
0I1NAdP0nXeI1Gu/+LQWcGJh6bBoIpt+i2MwgV2qrtIfjE1wKY3+a5KvjpUW3k9UTwL/a06+/pFu
cFe2z1jRh77DZyKIlMLPREyPlhjZU4am1U2AkHp/4AyLWbsvTizoTSydoRNbqu0VAZk9cwP8uMTU
Ryz5Fyh8+WqJSC5MwBgHsj7A1oCcjHEt21IXqOPdiw4Dhxlb9yscGbaKs5n11JZvG+s4BxcbEp39
AEfUA8khkjRf5iZlG7D+3jR71pJvYB1QtwKrTHZagQAr6PydKZGbib2B8TE6Jnoi8Ox+hyA3UUiQ
lmHFNDm+F8XC8NM38+3a/pFtXDTGQxjCyTXfMRz5pyRmIwREUjMWCwjK/PPk0U/ViwtogvLjWNMt
bm2aBHf6WujUDo9OAepmgkCiY7UJbLMaI1QauT2kY7mxFDgMk5OOqVQexHmMeLxXIRiAq/xJnRCk
NSxJ5+CgHoNATgT1IewF0BISJHK6Sj9IUD3pQwcCY7YvUUy8HpqA/9yh6EdMgL6vgyhbPRbU+cTW
l3W27OnRQN1944WimpiAwumhYQWREfjfFirwzGJUewBaZqQ4qnc+usCwAHaG5Urm4jIQ2yKAo/Oz
EdsjL98UxDV25C4tuV1YsV9jNM+4tMJCLRFQsza/p+40ob+hQfO4p5aoKJeyss/Xzv+A13DY43LG
crI6+e2gPBZ7ZISVU0BD8wuy6gNijE5m1hzzkk1Pu4J5EvMJ19TjRdi7Yd8fpF9U29/N5WZbDwHU
VFZIat/cAiDIPQj4AgMNjoEQQoX5/oXev9npso22c7sREi/xjTl0isEuELHtzB7aDA+Cg9hscdEk
jCj1nTA84Oj9P0wAwulwJxRfewXrSraENtf0vJ33/HXoMl5/sQgJ43x3F5UL/OJOzmWzicaxvg1g
8w7k+kmKTPlt908XC8lqILs52oO3okv5mJ0YkrmqI9Cx0NLhdaz41FVML4ajlvfUDZbGVnZKUpv6
4MRbHoaTWhVlu4SU+N7s02A5eIULQ/pJ5PJz3tZmPbhGmW3NXo5xVapbpqwjE/1njf4aY/WAFC7/
7LpZ8X9UW1HvoKMObe07p8HKQwS/co+VULCiCflBhnhsaJh5nVgQVfC5XzxlWoHdmABwehRQN7+4
g6NiUGwXwHunzob9+SqJleXAMe80y5q5mo3nVc7yOO80/OrWHaZHfZqhXVRBfOgamqJXjyEvRIdc
othNKkgRIWjvIw2ivmmido69xDdvPmT/Kv503WLP2uDpiApENwyIzGrYf0tWkoqFsVN7ELMoh+s+
SqoII5XvQRxFUqpIcSAEEp2/ossvALQmT+VUAzex44eSLXcUVjUOTyzFT3umrLIIeDiyVh2q5A7B
hVm+onb+uQ4DGZfUTv46+n0/BSp6lKBz6fALkV22ZQ7zXIg/vTQcvvj66EUNBGX6Vz6dSfFgPprr
H8VPmfpVKPMqpnUAD7IDQtLeFKWK9NGLO+PG3SBNKcc8znMohXPe/N9a8HUMPcQxB5vgFSXf0422
tEOIhx6wjtflzk02SVSiER6/70S4cuHXCiaU++qDBa8BL0wxGHyrS7nfssCXFPnnh3TE3l3X61hP
WH7HOOWBsWcu8KcuoqBTaTQp5cdGl/Eq7/v4S66oripxYL/lcaSrd43DPgyB6t/hQS4WcWaxlobf
cqRCtBdsbkajCNYKFO/p208r1j/T+TsEBNFpfSlY+QPht3qTezL0J/qVC6LJF/Vk9941Kf71iWBa
YHzmn/DB/qN1KXCzeC6ilk8PjKHRKSH+Lhe+plmfJXruaF4qD6JG1Tcqno8kNIp8ujanAFcAbOac
qffiOmsvIGHyc7nh6ENXMvXzUpa5Ihy2YV4Eayd6j3j9UQS1fjZFfddaX8VYQjvTKdO4/AbVDpyR
oq3vLMQWjKCaq4p0NUXJ4geDA4jpOSjWzJiLdzU7daWzOvtsyZWJ5uiO+nia9/lL2LEQgUDc+npU
VHkwesXA3reZve5qW0kw83qDtEWQ5hOoVq3BFsp/73HxK2ngzqhiQZuyHZoXrdzR9lU7BIJS+M5l
HA0/kvbusU4LqiKAs10mk5Wr8n3mKj8RWv254VWKsoyHkTjLjdRskYz9N4Dk1pBaFe6DBYjkEn4T
18aUbC408GWEbjz7SdwTvjUK9BulFcsygKeUvYmJOdRE766xwuz0lzUbicYIqAOQSxdUjL3JilOa
zQjAEWPKkFvBmDauZhSUoxYJmU2o4+ntNSQ4Iy979hQupK/MQux6xzNNPaOcPJyh/G8YEEeLcUyh
3fBYQAycT/ma4uQS4lyXAzzx0BmtQ85WDKXRo2ini6nrjWbaaeKHMen259gqgYFUO+deL4eREkli
i4Z7WwMCBB+wYUxPA08U6OzpmMG7dOEsXehYvcbp1WAcfs1X63xvLUzWbEseTPK8oitfrLddc32Q
RAJV4IL/GMDUR0xUvHZxhoxvgsPhhBwc1kfhgu0ApuUs/ZOmWahqFh1vYN2luxkgQThfjLvw/vrA
/4Od114NnWFfkMfIJFFCowTB9UeAJd8vQSv124XpmDGDuH3MMTqBBJHTH53tdhQqhqfDKFHrNOUe
B/97174SYBtDjbM5s8p6WXMRD0B74ul45NxvMHMt2Rg7vu1l+TmsSbFo+srLXpSPfBNViEVGerpk
4qjCV2T2wUinK7U43fut+Du78bCdtXS+LsPeB0r1Eny1DzF5R1UL7PDECMOlFPU5llZz5zAS9Zk9
QmxVIq8q0UrnGtdSbBJGA+XsdHz9zcIBnQ8cSZIImXnDYpy/Xztp15nNT9ACDli12mkY2aLT+3j1
+uBKBCQeYcwbCGTRRpUPkWj04sP8BmvyLR5dNaVwC8L5okyzH0mNaUUZofdH9quEifoXTDsw9/ub
UEwJVvgL7Zbv2SmgPiGBvncbyZacByCdt/VuQRv9F+8XZq5Gm4PhyuXJZbg+x+aHW4/Ixrl7GcQF
c7OGqS6QYpDZQa+HPFXpCEDxz8OCc09jpcR0YTajx/7xo71m7oGnZP+ywwNZ9ncrMmbcgDLrVzYt
UHhBQnSTI2Z31Bug0I1iGmQ4O+/hlBm+RexYNKC12qqOCulnyydSxuBHQw+UAoT91nCpm5qLKt1P
GF/qzhgxT40Xemfy8+rpoRQa4v6D3H0iKyiVHH0IyMbOIzD8e93FE8bSPXt1PYsqXkIVkLMMqKP4
YdT7IclsPC7nzZvP1FK8TStg9x59vDRvgqZqZnbfSbzeGrRb7uNM6pYDjrvqtSOb6OgeHAyZ9O4r
97oRTIIw9fUgLPhLE61BfT90dR2qwGDMvhu/QSIytOSV53gR26O6kZAbnV2q56HtQgM4V1x3OvcK
L86muB4U1BFQDvuPwPnF7qY7V0QJD/nRwlZD3jlYcMBEMJiZAVNYRblLgYLRf1Oxbdt2rBeelIr3
C6BOU5loLJSbzZ5L5d7k/pJY+2gBIP+3kNZvQ8DDVOn/69Lyf53g4n7G3fSMAIyeslRoIwFzys8j
3hjxeKS3/yHkZaY7Fm2bYuiPH4DfZy7Hf53YkY6bMsKY497Cjplk4ecbciRgIKmrG8EvSHFpNJJE
gUEzE96zUVl5BwYLtd3JnBYRGsL7B7H6AcIcYptOn39gg4n4yqoZP3aVszEgWGmU6bMPMPA4CTfO
m7IioaLprc0C7D7P2YwnJtB524BXaGmGm49km+/3eWZLr2tBRtph+iuc6CyjNeLrnkwwxe9Z7/4F
yyqW52astVzZF3eztTYWQTtMMPseY3Bl8W1v4P9s6c2I5cHzEPd6FxnyKZTvMZjWdg1aRynj3xU2
XWl+VOEZ/hwGE+C7Ce4eAs3q5ZREu/TIQeGrWYS42W01yeS8fD75fxk9qexCCDNymbNT/tUFOAVU
nOXYw2xiEGmplK3mfz0TtXzdBLVG6DvFHt32ug+Ri0DM4YS1o2sGlGujiUyWRXKaWn3cD+N/wiVm
62BYeU3RBsqFFvfP9K/gwXgX3E4+ixsqRxOz+tTUH6yMBFucBt6sBlZKJ/e0ZEkubGrAPGT37J5U
AEI35onxYfXOs0I/QZfa33x5wkAXtfdm/F0ti8jG5gUDgPK98RqamDg4wupbg8HW3Ue16Ers6XWt
sOtOqAIA8Hk/gtKKAt0QnBBL/7iqe47cfw73iIi7qPtJ5GGoLyfQoHXz0Mjevg/Ypxj+QUFW1ytN
uD9d6QjamYgtJXVTuY3TiTvK6HRPlApZ+TPMuYPRoJZ3tZpQfzK2nsOKY5D6XGDv7EWMtPX1PGT+
MrZZ9YPXiApjkR++xKDlRPwyLe1mZioP7w0f0YLVFPX4uDhPvNCsM8oT63/0GjOlCClKu/Zh5Z9/
WTx3fsaHyufQS3OAZtCyZOsg9u5In1mVukrImL/iEFK0NrsUiXabgTnicDThfFl0LwTyrv/bCkne
T2o/y9ATmJupYqPzyUCXctnhVtBYSDQkyBErsOYImVGjkLDOjajjfOtPX1fPHSkj5AUAQhXy92KI
Gg13x3QdDjIlL/JCcevxqg76eS9qcP2JUqVWeNxSCvFJUlNEQ0PeoB1neiaVmxBhq7TWmHJ7FDUf
+RaOAyYx465cqwcM7ufKtgCeF+YrVXml1RxkbZ9h7e+74JpjKnvZf1dWkwiQZmKPVeG7fNRuCQts
wACVQOqNj8Rmb9TtpzBBAoW0DY0GNV3mValJPcWDKM1y+qNoNCa1FAeLgH/rzmVGsooCQgwQG0Zb
LM3AllHaiU3x53gM862iA8QrUeBII11vt0nESGM8k/MJWieiLUXWCyWqjjR7uO4auIDktueu5/Cl
2Jzul6mhI8wbfhL5ApidX/zWOhB+ktjhdFeHFMU7zZNQHntUsqAEaUPXHrGSliCTlzTSV5s+nbcx
cLy0VjsFIDhegK1P+u7TEAU3saKD6bfS43NuMFPxAFL3L/gWC6hIBNPooPGGmaWNQgoMjF2WDSYT
MIe9Ejda6s+gK4GWif/aUR+OR1y7G9ocW1Czz4kDv+wrW+8rd2POZW6L6c09X7CPbCxYIrJM9NGy
KSuUh8+Z+OQgR9ajTc7Gn41SS1qyecn9ddnJ170ffrqK01DUDdRu8GBZMYPe/ogdLYIRmziodCnP
IbRNnh1BC0JaiszowaVUSou1cdBwzc5oQ9LNuouvM4P9/mxLGcTR5ZfU70XGKzw9R99p25eZGl9N
SUr7vEHLNHsBsW1HVpw6k5I6Hireq6KEB80DXADFx/KpNIEQsmGx4Rk+Ds/8QGf7dhDBNuCA7N8F
IYOIPrCxi+6hsGAQHewaN/r9oMkqtrTP3XayMVbSns5Pqlvzv2uz9KpUeYs8yy07wxUuADZFu52Y
8Ho4BF14tAjLGzEO8pLdfxVBJQ3w23k9MeNCoBMzJnnx7eb/5hhm8EeH+oLiFWduK//+Ut9Y4DRl
3SV1x6VWzVTG8cnvqqWEg4C7VvQqQYuD6wuDeFGWoP3yNzBqpXHI7Gc4iS3kPiv8H2HqN2stixUu
zJqXFk0m0+xAo2L6T5X/67326V61B3suYlc/FdV8OExfV6IlvzQZoeIRxVsf2jCpkhNf1xSJ2Uiz
bh9/c1EJARKzjHpUObPxgDJm6bpzvUmg36h//78DWIYnqsHsmeeeP/Lzoe7prw7JLGDPDDJB88bL
x52ZmlIgzujtnS1OfI1DYjWEuxTVy/Y/GgrKXGDt0vmdaVe0+fmw3cJzcjYGPvuFwdhAwIBz0/ic
R3s40j1/9pCZ5t0wIjldlBHaVo7rAwfyZqv2ZMLgy7eQwTp0wX5R6YxL9JzK2WMYvwPacYVoJIv9
BptbFD5u+rx5hO3VF7nJYJAK/gbUnrR+ulPpsWzt7RVo/9CCZqQeF7VUftqJZRt+cOLZDieN9Uvp
KCHgKSHrOiABD+bO3guunZt8ScH4G8tAtjyjKPXdUydrlt5JmoqVRewwhvju+PbodzqNrhjDgJi4
gBOIBYxt1L+Aqbu3wjQ59M74yQ8ZnLsCWzK/5F461mOAHUeJIH7WbWFJW0+D6a26FmRE2qjiDVAZ
BZmOnIs+L/UFQt7sxvvAIiKvn3ucMbYN0nnU9oQKPwZ7qKbuwuvs9bFezEA6xE4ALuLgN1LX8+at
oej4cxqBwvadLOqlvfFGI00COvqytN89an3vtKR+1yvwmZ8Hm+4ZfE9ncXKA/VATm9fNKZm9K82i
x9eaqldmV9YYPhhtvyO3g+hiy6/v+0hl4gooHAwMY8sWBury2TsXJj2NzIHx8TLXxgdU/sYm3VSX
TpgPD/d/heCyTG2A5AdHcd3k77PjiOfc85nQQkyGRvadxCkzre4zy2a1MuRqy1ZVLe1ejZm822Ht
+W0T+XcgObbovrDCzvsJ54z40qMEGYjvKhoxt1OVMV2BLY5mGG3KAUY1MQTdrXGuN46HKcoYLKt9
LK1CfOFHQSr8kFLBqxG54Wmmh5GwNwavOHCW/XbuBWe8x5RuPM5uCbCuia44C7O+80fSAxls7X+X
B48Qie3vwbgXuwGglUhQgV87ACPHHuCej3L1vZ5F2nU4VLXzJ59265yhOkOI7nXyraSYYsEdh/A+
Vx8UBOHRVTZEnGMN2qwBM5NUQvIWyUmzzCUMFRNwWZQFo4b0FCh90CQRPMM5S+LQ3zoX6SmOHecZ
l8lImUV13A+dnVA6r2dV9cFrjGbH+piaUZq87jqJiZEiYA0FgabxSNgbH/n5yHWpIhlVvUj/9jZ3
xkVt9XdKBxm0Diay12p8bWRq3II2OPwF8IAPFvTSEaJLoKMpOB/e9Lru8Shyy2j60G8Aonema92e
omlkmv9f9Swm0wAB+Ik7ylJcpGNVPRZE5uMV4sr2Q5NG18b4UrRbM8o43ddTvCymIGVKQZyF+woO
85AHpxHHrOvBpz0ZFuJK1ys47VLxZJgHpaUvsbcxLv863pqXznjQmUBCbvzoojKrrxHtji3v0RgZ
iED+MvFPesWSga2ElMgTfM7flHZz3Sbdg8yJYQ9lxqxQedZyrtkRPi5DfiXTyyQw1qJL3zKFBDLM
0ufNS5SFNkiLWgyoQdALpk9yWEDyQU6BtX/2jPG43U2BHCov38615Ldbwz24YuOoqX5QPXicAnbG
ICeRjAP6Ull5od4V//ZX5qVizQHYzXtETW8r3TtWH44JF06gKcZ8faRoEb+vVNpN1MSLlGWwmiuH
U2QZQsUmJeP6QO9RpdIGelbPKC6w0oieMLbtxFUQ9votjQKtoOS0pFJlvi8KkUs7ID2aKdFmbdDO
Lvdvyif22I47wj9F5wHwDgzXUWQLl5uCZ6HvdPRAXIuGBP7xr6dNOrRDWND4MNLmPWeNKFvrDVCH
WYEc2Yxe39iXfO4ahjMfOvU+hCI2v2u4W1yVTnhs35DGrTfXUiceDL+DEmGOL+tsWRf/2G9D8Nde
RcKZsK0Vuc94WFQDJlzrcLTt5wlNhr1JZiS71LegC336ARJ+/NC+Vy9R5pR5tcSI+pcGPMmzvFL/
vLjvmV6ZeEO5m4YDOjqqLVT4v/dGVOGBSRvJkv+r0z0JjMz3dYkn/RewvoAcTdiwJc7gy7+VQ3FM
sfbozQKB+H0L48FZrEOID0Zqr5+WJSSgYPLOoBpqM150zFwBYlSLZfdmsK5KboDQyz73pqfoKKu9
ncZti75EyYLdBASxDNR6Aj3ARm+83O4+A8Zou207ULHoU+bjsND/jVG8y+kXwdyKXFZ+JVoCH7bz
aEWGukBT9XMvBdySaFqQJvdINjP67HDeaknKPgC3LuH9YpWUT9xEtgzOW4Mci6qkzJKo5hMPHSu/
SOw6IqavR7f//xtd44ACsykF2x8cLTsBlK4SwjMDQwtd1B0kiZjtsXC2bdwhqTaxv10O4GkurCkQ
e+CY9m3oI9Lgj1/UVml3+aQ88Cx2V7z70Qzi4sLGs+aFTsRmPwF84EMznkSBXG86nVlgDBS2pD7u
50DmyncuCa4GsGtNcPHsi694QJlBMp+wChju1cO6KLZp0gWhWrEKG/mB/X806RQh1OCx/IyOLpYW
zW1RHhkfjGpmPwV44X0M10DsyhZA0L67xhDKpO/fPYpNBdcPRwQ2iFFGkQkfLUIGkHveQNqzhQcU
cUg5qPOy3ybduMo/+nfXh/kdnATlMyWPAkF+vtc1KePFBflLfUZD/wb4D2txg0m1XsFfOBpHM5dk
CRXTLW72cudxPOeAoWHVzNPk8gtXNWa4zzg31vSfwN5QpdokrmoQJHbeQJohkCZ6FWVq2EgxyjEi
lVd81WTLO7rdENMJ6gGeUjCut2iuuyoMrwTEvTxewl846HUYIBrZ9IOGI8nDB4jNcHbBsAMKePGo
aWf4elj4y3yYfgo4TdN753BA6ndgkU3vLZ3fRXavGh8wXUtxxR1kBH4xC34IOyofyd5OGYM19ng/
Kliq7W0uizQTHq1zmN2SUeKrFq+cJ2d+9RXoQnvlC+BvdF59xnfWE9Aw1DN3H9S5YZgDoDOdsTtK
mlZgUAKqNZNQcAsPLPmXxjz2KwOxpI9cJ0Zkqxkmiih4Vo52nOOGQ/SpRMWPubd1gZTCECTx5FJi
mt/C8Ss/+vVzvlcSIOD4FpyaeXZhh4KpnR6yq00RjXG9vb9psz3WCGHqaZfWiRseUfUnT4jbCKNB
dMtXWxsDZxYAj7El4bnM9fVIUfbTxwDoyAOYFnDAd5iGLPxpRjxob5BVkpLmtC3wrchdX55wUE7O
4xhxZp5shXzo6eUA1DOH2wy1wmc2vxou2MiH7kCGHijyg3H9cWs3vdV8irwZg6RF1BgpO04wzrqN
AvxQ3u2mghMc5WOp5GGsBLF0EyE1sMATU0dYvccthRLHtrIAcU/Irs4foRiYv2D+cc6pa0ByFm2J
n/jjuRtJhanEBblrgbHPaCTDIRbLmv/7pOdITQX8XPNbjb3raNIZVA+1/y6LTiK7nvKaiYmOgvxH
7ENuvawSlMkG2Z+ClGceEUP9hSiO25dINtz6BtqOt86MIkjHdhoPiNqB0EScnTQ4Lily6KOs/8Q7
c469l60Tl4IPcBO4v2mX6BlTUVyXRj6Dy2BSc5y5Lxl/uUqg9Rt1DFvgVf+sBnY8CGViJNCj/FQq
88XHsZH5En+zA4A8HIuAbhho4MTFvFU5uiGB1YSB0ZW1uNqELVkPHLXf2zS3H4He+KiuN8CyU0gz
e8Vl8H1AYVXY+PtM3Bmfzv0kv2uj1ZSUaxYJDdCLtxiVB0ZjHgixEK98zMPs3sXeMgL3LHJtXT1C
sAJh+S+pgDzv77uwhNlke0NsWH51ZJyZJbU8MLq1zay6gxkrZL+FMfEBOgTOG9fNywdME7oXWDlj
P4C7Sh/tuWjedO1HY43D/GloOXfjnN7iCOLuE5hj0h4nqFPlaxxp4EyeYTW+g/YKQps69dCu2v8A
/YJfXSkVVSlgXUGOPpLb1r58Jb5p9ZA1l4kfWtSstRBu3ylyfTqajs76g9gFIlfrNdXwmLwflRWX
eXDyjO7Wn/QWOfz06tOtDCbRcJHMDLWQgJUxnoKP/D/GXs4HnbkvOjoD8yznPniLZPIvis2DZhKy
GSkPsF2b0/isBYyEOAOgkIoLd5asGzHmwKnfghByASFIClaBr2nsLlF1MSyey7XN++FzM0LRmdyv
D8KaKOykjkyRDK4Xf0enOpBlZUUocU+cwIKD/Q2bmNyEXQg20Gp1Gf8M9X87rgnkUbdbcjQMlUez
ThCCVXkZz65ebzG/Q/TKLskMKfMJZfbr5I80IMUqmn3XB2L2Dwlsvn6LejvxfbIX03yITohLblLo
0Kg9ya6HDiyvezoI5z2qIHMJFWRlXGN4CRfs587FjyLt2P/W0yzEkw9dVAMquIeQYAOHfUXOISi9
3+maHm9e//eRWSvvkY1ONWWPyaqpzvzEoZjEdD+a4L8z1kLK6V4NxpHB4KXRPtgsDTm51iCundLt
ATSGc0WU09/50ngcXBmzCERvkoM5SdEXT3hTnPwPkdOoQXBssIgjIGItXphIcBD7EaAMjuTfNqIC
iacSTkQ658Qmq78l+mHR52LJR51YmySVPeAOqFfCkrXdFWKaDR3VN2bsNNAjNocQ7HS5AFbvXiks
ccUeCfjL9JNYr+9cn0HH+a8xqjawQJ5l7Yq1xqiNsGMNnG222DWELsOtoAKvwve0hyFSq6NjfnMJ
oWTArYQShlXPtNIg9hB/FEqsI0QZOWixHU9mB7BqC+sKYbBmJyGvJEcJYdSvPw9POz0husg4bwaq
asNVieYlulvEy92NcTbfzPEaifvq8xoBKtrSQJE8jYCLgL75Q3kHjR4C6O5VTtcH2wkV0ujxgpvX
qBiT4tSicKVcu23zxmKTuQIVdTrs4GJzfwkkxmq33vUxBcg11A+byCkiFBld2s2khQ+txs253KF3
KgXlAqHLy56iBS4eS9T/on3ZIUk7iqijy8acI+QtChkbYrgJas/03YzhZT8+zthJhH8e36xxCebI
T+qgZayKBi9C19AMPmoaXogQ/ma75zYgajeIfbE873/NbZWVDct5uULD/mMr6/VqAMKuxUc2FksR
baU7c3pOwSuPRmiRzInzwD7q2255Bn6ch4AOjCQweWszlC+b9eZadmwTRxn5KbaCEpTVpX86Ys4M
TT69q0oM2h/W7smdvO0B7xCvujrcoPJqFaJGX6aBeQMT0ilkzLCP1TCYJGZfQVCVVnu6fI/aY281
RpC+Z0p1hajpJlRADLIb3DMZq5aGb4mfnyU0PqhlPEFuxlqfspXjcoIk839Bsfm6hGaxLQSt4qbU
qH4kvm6Ko99rhyW0QjOMjwZI7v+WDfDMu1gUPr6CRIB4/YjyC7WUsj8QW8AmxMO++uye+sBptDup
Evc5LVmlmnSMS98UEE5OoBYjItJSCvdg0fdThfl3e+lDc+/5TuF0i5nnj7n4jHSO0NVxJHF6Zu6f
OGx3V1Q4BDgMe55TbcekmuypB/pG2fnkWpcV6U7z7Pjm7SSimg8ORXJeZpiWCFm//QaHnFx1zaq2
go2gMRMkACKu2Q5i2bRl4hDuFIHMitsNvBGDxm9TFNMAGSvmY8F1Xh+TmPoTUuRlH2Zw7i2zMoRK
bx0JMu3mysst3vAoTZ4phDF+QKfru6Pavft2G9/gZcBPw618BcOGU4AZDK7LtEBou+SsuqfU163r
tUCSaAwQ5aiukau70gOiZ1p/oArG95L0/dYYOX9IXbpHIHxwJKTtrd5kumRSRwNNUtUC2d+JXDn0
1OI/Ygc2KEC+HNk+93HZRt1iOJsrOdDc68L/ZZxGKhDIbk/413cKZKBiaMjJasmMXUBzhGEn6+PF
zHMDzZOofq9V/6dBXlfDWGDj0ZhKOxD381C5InzKc0hJ1NmWLcSq/b8lZv9otHfrLVykT6zlvnkB
2uV5bIDJkvH2Xf5vP69cIT7kaXJM6uwMuM2eF9oeKpp7cQEKkMG4PsAZ+L7XM+p8EJqzzg8NTa8A
L22nnD5RPPZ5K03DKsO+tA/3h1Hno3LhyiZQ86uvzFumVq/d0g60d4mPrwWwK4n3DPrGmlhaQOsc
85Pu1wCdFDExH34Zn0qEvWxncu/vkgolfUsrISdNEq1XSmp6x5gSFoSawutvXSgMOqR3bluxfq07
3/4o2eYHYos983F+6zgSjLsB/KLV761f/FNAI5y11wGzoTk4lVIjRty0ki2NMytv53MTabBk9bJe
ATNftkJm5zFcVcKkMcT8sZpAvpQQ6AhKP2i19DsyZXIP+4d0DzdJgOVqxX/rOofESCB/LLE+xdxu
nn9WQBQVkMgHsJgSAU145/7byYC5Zqi73wQb+bEx5oOvCL1ddVk2Qqg5qoDlaf2Dsfd11wllwKch
FsTUHrp6mxnRo+TeFypmEXFXlC45RJz9IzOItit7PMq4x0nfbDZ7Ec72RNXDiQmWXRsWBjva3wZg
ATj8KAbnOP+VzloEogQQ7X33+dKRfR29cPdaYdf2+jCdcb5xVZ56//pu99Jq43NaiELogsdEJ0St
G7DouX7EIZkA078bRd1hCFbMcvHz2l0SK+sNU/P0yo+NGFSZc3xo8sJZ/OvASaFnFQBZMSA29Bzc
/RY047+QONHvu+LJY6cp4kriHY2OGFZMd9oeqqpObRHQsoS19WHfbLZURkwng1VjonyMoAUmGVDa
3dssIBWEd3Qe0JGzPq9P8PzJ2GGfU5Wa6zOUi76dZU2jo8z6wzB14makfa8CMdbh1jKRa3FVXPCG
b6QdZWEz/mTMqUCxCnUlQh6ugaIhST6BtOMNmz4edJODCnPwyR/GA8xcPkABha6BfpbpC2QfEXec
M0/AVh4wHcXJ5DfBAwhNr1RoRwUcxxMMmqOBgADkiPMtsKM3xjnFq7KIq4l2LJASPAaeKOVA+njx
5dLqFdJIU8O8E0IPO7NfKb6fLwspW9gY3fPuznKmZJRuV1UGtp/YJsCXp5E5rx10ZQzduN35u8Ya
qvrfbRYP8syD9GGcnSGKmra5FjVHH9bVt1Sf9eTXBz9lVXP264ss4dhkMH92SxZajkzOC9+gmgc0
U46+WsfOoy5LngzhDs6n0NCTlbYQBNfkrBQ3ECjFvLzxc7aZiWGnkLC234GZFt1msaMA6A+tEAMJ
dABQgtwljvjULzyw11mzOg2wnhmgZ+g2TiEYa5XhaWD/eL+IkedgsMILYBqVyj0ORgR7sQ6M/OUp
u5zMEKgC1sYXgtusKq1DSVtb900hQj8K3PX33gqYDAC81RzkUO9ktfuJqveBJstxKJ+WgMKwg9QF
sbWh0LxpmI9Fcf4Ep+jryvlq9mjc8+S0rFTGfnwKXohY/9PtVzUIwVUa7czY9k6r/bwO0dMXub7h
IrxSU3XwxGIUths3Y/npjIkjYq+gYmTXy2nPg4FFuTb8WuvsFQG80S1glyTJ7MuLABV1Jn0BtxcY
69c0D4KNA7tiH4PEX+nVR2VkhHLO/ikiGGbLsZ30bdNF3P7Aip/4TFyLEsKBYU7nTNh9MbInAjpW
LCwfqLDkRhGv7v4roDw4Qr4+xvsUWHNQdjARAjwSv5vZaCr1nvFv1cOy2rQjDIP78Nq1gPL9f5Wn
CWVsRbVASPw1WZ6ogFEng/V4t4tpJJHA6NA0LjW3jOVS82pApQrIwfD/ZryBqPq6k0CCyTwRc/QY
YGKlYPHGqcEv95jtZvMGJcXpuJ4P6xFb7q+vIjvXvK2suQr0s4FhJzrCgAGoS2mCPw19lukxFCJy
hAh/jjba/IlV1zkpncTo29eAcsik+FvI3rGS+6qUWj2d/wIU8mngBcRq4GMDbstjkcapTsC2IEhl
Y9XvQcPPNJhTV30Oa4gFcndJcG+OnkHUxOZjI3Yzv+yv34dhUXm5CY4LrP2kbnWPU42jA4mz7Tw0
2l5osjEIqAd4UJj4Vz6GPONNiVxPVUwyR+txFNenvMKMxY+GEqdN0cfGZs+XatlTjJLpJt6TnCha
TA7iUhNyaQgxeLj7zkM+Jdf8qGaBroPK3dPl0o3jeETgXoofVtZNE0IEWJya+ik5VxV291mqVVyj
IrfbzLtbxPR0UB11Qb3ZOwqrzF/AMc8ZObKlVX/WT5c/C+qx2PqYwC1uvcPwsOlJjFeb8yIwKknH
37Byk9sxZ5ImIaWeC4oTzCjL08kc0d+y3lCOyPdc36lXRYT2b/u4i7ZztJ1eFkQQyL0gjXJpJsfc
gsm2j0KR0FBPMCmdEPl2YMK5NQZ7Na3NCMsurCB8i8/hgfIxs0YCFRmU2+24xZfO0Bt7yJzWSp6S
Fz762Ovu1rk1IXiXhOaoGJBRy08HOZtmwn/z/B+HE16AoEgBC5vi9AESOiHCu28KxDCH7Rg3rJRA
LMy0NNN9MOcdQZ21/Zugd4s328aYJI6GQMPJkt6VGqSlLXH6NwlCJoifrjPVovdctWih5GLJSX+/
TWpVUZqlmDbdqf/iglv/t0X7kA1Sys0y3XC5TpOYRTM/TSxjyTaw3Tx71q+3+UDtJFL00Nqw+2sC
drJX3lS6AZnER0HBlP9ZL4TLZYxSmS2JKXKTWVr4PLMdx71onduQagHTLXL4TgDSfcJfGnsSPM8o
QLRlmTcfHUGlFDF0mcInUMAJjnzbWv5wS3Sgih5PlBkJtfMcNt6tGHRPTsTCBZHu+8eStuULsCMr
rSBfTIoFEEqPSGWhDoOHe3bdHYTWLy0L4kdTfgg4cVN9vM+y/FRaR1ldVHX+eBSPROwsmadVnhcf
xRtIMCrMLeaPqJ1vXiFLT0D/eNYy60e2cdcQgsumsUnYqLSTgQQudoOCYOjNsuqCGpIa1kt3Kj6z
Q52yqGPX2H9xmz6etnBNoQnRHizH6ZwuLo9yxep+1ETiT/Bdan/DFotsekwNiu6kZdcR5xup5h/v
pgYCdFCxUQtAWr4IaRDuh9QkcNPiZyQyrO9I7CE3csyXmaJv4pP7yfYj4wbnsn7Ib1VkQdfLAPph
VgML90DKpLMP8hlMhU83q4RWG2nu5MbSLk7Dg6ZZGBZuVCML4ggmY2lNR0B1u68xrHHi5USIY5mG
yA2+OejRGzx95whfvApfp+Jyx4KaANVAtt5oAYj7QenO8wFZAN70rx8UX88dR7NTxopbXWY5HXcX
s40Ms+vVQiG2ndjbqF4ofnDl51193RWDkbGY4sfyNa4Uciz/1nSWWJoZgC+RyXzQ1zB/AB9GOwT1
UzC9NM8XBWQRq5ZlaY1eG+BhMM1/R8dxHx4m04SLm8AnE2KDRkUodd3xxpfDGiG6mcEHLFRC0Mdc
+VHbwNKLsufTZv9hrrrXdSyjfJZiM+zf/3EGLEIjnrP2sMrFTS15ASt8nClKgD7pLNUCB/lzG3NR
ytSPmUX2CWmU/PuPnPdUcfL0vgUcpDAd+pumbbKn1FPno6m9o4++NizSrdSPWMYMhpZKMGgR2lMH
u53f9i5oRwS+vUPUUMK3QrN2nuHfHq9UETUXAst3M9iU7LPfFkyM487DBcsPSq0gHZ9FYCZLoI/v
N2LI1Jb95nSR5CXZUDPgAEeRLry4TOAT0DsDM+uUwr7Bk+3A6G9GVlvTZiY35xneWIw0kfJ4VFhu
2LpV3ljIPK24R+Y9m9FzSGdcinIhEW8MP28Jv3LKRVvs5iGXOkM7qt964z7YuqZY9oZRlIpbf2/o
/xaMQ5zK81BPdvcZDBtYiWiat6CkbzVWnh/PDrU33clEW4+o22lfDbxqGgc3nkWpgytQ5UdwfAst
X6gY6Oq+B1xZ4AUMhp/ZjG30qKWFaYWaNnxFTMOeWCV4UaRMjzJGPUtl+wcYdKXzIMPqT/L+AGfL
3ENqIKTMPpy1oFBOXqlTRHk5NoZ+hVWKHpvsqJPzM5kkZnkiRrkZL4WVYrlVXNqmzHP6jJilvYzh
/cZ8yx2XlmINsw1uH3ZTvwBwUhRbDG11qDTxWQNCs0AM94QlxiDqqq80f6kU/+mKEr/2IgGxFGkh
qK16AMNj08rPkjXJPrbp9s8lRCPQn1ZXse0FmKug48c5Gmc0HXUIBE2lg6Ua/Zr1rGqk7rjgUrXH
tswd3bKj9dHsaP9XT3esotyOGUWkt8JqFKr2gZaI/+nA+Uwm+I56JsGAfedh//VRCQ0Zo0pbpd2W
4V33MLvT/NQAd5Dd/8d2dzbdPKCJ2oD+aIY6Fjh6YhJjUut6GiX1disNlFoYlesxKxBpPDBkO18L
7/yr8VDrFFQLfKYXxphtQ9kpm7n2GOX9SifZjdKiVOGcHQ2vLpO+KPTlA15Mu5pbDIeYosyn20/j
2uY9hLjpXZfKrO2aNKko6JuFTwcyJVkRLwQAEH16nQNOpJx0xIYpFdktyeIgSkaeXaj+BOPbki0L
HLzCfsnrnP0QK5xCRGj6ckMgrQY+LsIw4biuKaHf2DtSmIfcFk17lS3MuAOmU+43J399TXPbdYx3
K8/pGQBnP3Jd7y8OcVNfTQ8NXwnpnjTqMkJjkocEBuKxwWTM7vyfg6+M8VqxFgIh+xLIXoZl8/GN
dtrUUsBV7KsvyUKiAOrAMPpU84kqRPqujyS1jeXh/AXcZNtKGsOJz9NSLrGOUxSvP4Ilq4KPnnvV
oWdpP3zI50yp/oEsoJMDZT0vU25J5+kM1CiiqSGPHrscSt6OALp/5mw310183YPFVzR0cE6g+vi0
gxxldmWxXr2eCeq9952GkXrwrtCaReyzlzr4nVYUl6tjQmVgHh4EFVuyFtVWZ8Bm0mly63O1cfUA
LIZbKMuvacu6rj6xpm/LO6is4R90kmgrtgSxtLwA7yZqNbkSH1xcgxH779p5m6wiUYq3In64akjr
gEuzsTB7SJJnMlCKU/81RYEbNuY9a4wcowOsE3STqCPv9xUy2OpFBxC9RfCGTa4nIeMPnBA0UG7S
BPm8sxPqwK5lhoEHPAhHR5GebyofB0sIwcKm9tTitOD15ktP6pL5NsllzEVi+CKsKe1wZ30LrTSC
oUlzWyrXySkI9GhusJN4jwFnD45qL6gNOblWFpOFsovjMZB6BJf7udmuar5ZPSNvBibaKukJd9oj
cAf8QOUVlJsg/OAAMtJljSWOD+rf3LI4Ad6eSc/aaJ/iFZGM1LsvhihVo4wWwOxHGnUr7KQXrRt9
YZZH050pY7vTjWQFzg27wSoM3Nq7VwlOFBHVeqNZFsq5JODv6VtYL78mGaodUhtJ20xfZ0z2moV7
DtidsF8YlZfax8wwNd7+SVPxWM227RTvvYd6OXG3l0ZouTFLRIFs1MMiAUo4UKpmi/S48DuynXtA
FLgju23Ed2EXA3JZn7uLx3dNB8yI5vnpU8XrGliA5YlS+bfMQoeKPunGfmHiOStdJPBQtDC3kJvr
Lf5huN2hxp7xabaCa5yWqf3TOb9yoYdRXU4MrxYivxTDkOZ7vM8+ApoeoSdy8yzJFfDWYA/qShuD
0fECtiTQO/8lnG7MlTKlqaihswXsZdR4Kf6rCKGOJC5nKHW089Zq/dKjzQR4UnriJSNuAGgQA71c
KcFbXSoa23eQpPK6sc0l8X73cHinhiOV/kb6AK3rQS7jYfOVbdazljumR/RFhHkFAGrL+wSh/uhG
zMm1w0r95fZ4dquyTx+9RRkE9r6GcsKIUKbFx3DWd2ftAWqLZN4IlZN8TG3a4fDdyWkCxIvp94hM
1VZ5A89OTHkJa7+Jb0NT7LSpu552AP6x96kluxNNz67u9lVv3LrgoRfMuy9BOZK/lkn3Mex7DWFl
qxrE+QA6GSwTQcjTJfhMmCRCw5WMOv8sq/q1f9WodAvzEq9KWuft3wnccsGj0sQavbLCQPuQjhyz
TqFm9M9x6FIIHLNTIUWQfmKevI/dfrwxVsiGbheSCEmpUsfLHOG+svWDj71hWAPbFuE7mMV3C9BR
WhXCoUUa0GkrDfpEqkTapIBbWjmlf5YW3hn37XClZhOoUoVW8JzMHd1ncqlOBJkpJx72kJp1T3X8
jYarPH7WecJQWej84G3z8J+VDUbi7BxT1hjxvyvtWDwfVhDUWwjlPrK48EGmaKHVhe1XPAyt7lq7
EfrQ3o+fdU3DgPV+j6vCEB1KP6nDlFTXIHfxXbfqKPy79cAfub66pbSgwaVqn56T89kKdfgcKJQe
PgeJf66woeo9dVMduy/LiWqEiSb6y+0bKCsU8Fx65oVax+832786e353ZxmVtEwmLyF4in/Cp3RZ
iO+jnLqvX076FqdGmVWo4pBAyvwkYaROYzvQurkoIxPK2tesxoge8J2gaCt/eTQBGuzHfQ6jjRhi
E4x9DA9A/AUs4oXl0i4VW0APJL4sEDNyidHc/8pbGSkUHq+ZU0pDsm++vkhDKfHIbWVQpr4sgKgQ
J9hR0umnWaUOrKEUeAZQmHXTUU6yD6N3XmrRvo6hDlS7aKQatG4jYfnrVwBa75kwWhyfiQScWrkX
Ee7qISy5Gn8Ri0fhGS+XIcVcodX5vEgn2mxENkzwvr3ipuQoqofqTrPOo60BUhpXKrr8RLPK3FqH
SshFcQ6CFtzroGoHAKgPrknYWM7Piusa0l8jMAn/YUPpyyOHJKRQwK1ZvxzbzcHCMXztC+qoAN11
3ccaN6n5thcS+P4eGeyRyrT+p2DvGCUDFugrbko7oNwer61Kb3ipagBSMN4znn7/IUf0XoWhapNR
nQYV5IY4UuebvICalgi2T3lZOHtYOwZlqyHEKEP0fGqNFcJ6qGlpqKRmOUsFZXZi1Ud4l9uA4f5e
OhUETeEJcR6nL5WKZTLokuJGBwFQkQkaxNDR6OsJ0PqzIbzznFQ9RVVypHwkGzY8UCYAOkiz3iYa
XCtMrlWTulSUubnnZV9hYe6kTLsxDNkkCV2rIfrI/mEMI0hYk2p7qFTh3PCyHznxJejg3A1ar7//
ZvEnuHsDcfvHFmtsaGZ+39uZFncoyZTT4mFLlHSnyMRSpDpHGbaSmrT0MtiMp4KE4hJ4MRq1zUWX
TKKGuDSktjhrClbMVEaY3nNIld0jLB1lLqZtaNXOZRRxMctecEfBDI90DPCXjbC7qUfOgkYQWMEo
juQvGJTbK2Celno4hfvPSM6yD8bNJzqHZp1q5adJNMDoyN/Hfq1Iy+iJ0WVynm/wJUzzPIbzz8TD
WPCCMVkejcSCWDgOzNK8SU4c2C53oGgp/Q2TPPJGNkE+AiLBXIdYmpdll1Wf4zjyzEl0r3fAxlJz
nI7qlTsljjYt9RjfPQJFmre6z3ANEkEPMkpf6HCEbOhn9nRNzdRBVgpubbwbHrPeuM8W03v2Bc84
0d/Lxik6yj21bXZNeCjN9fWg9lyUMgaU2c2UK05KjPXK/EuJBYfRkYBhH2Wtgp2zXdsWFEQNtHeH
Fyhqo3EM299YmyAdibcryK51rKoCCiYCaNyYT0y7jtLFG9XRpPpSmEpRi1zZmGfplNstjmqU1Psu
STJep+01mse8Njm2MNlwv371Z7n5NoUUNd3hLtmWptG9up0uPLCnEHkHO4wKZIJEQlSP1SQO6bGV
5LR7l0vC1alEsL2dgzano9Sr3LgBw9A5Yw7USqWrAnW3H/NmygUxmjLEvLUIEO8Ixw31UMcvZcQi
d122mHkkylp8U+TkY5kvbzNAofktbca5zimvYo6KhurePJtqSgsKRJxRYd8Jr5Iy6H94QPH9QNcP
sCFG6spfVPrjNo7CPnc/xbMfMJRJjeUcHjeKBboYsdo/eFIGjBvDLwaxXKWWKXnRvrq/kKrsuSJK
TWbDy+1CkIbwP7h9byF87QHL8x45z2kAboIqHVxJ1b9S0dlRrUOsNzAkAslK98bAIjb8LfdtFvh0
iwjjtRg9DGcTAlmt4Z9I0+jM67YbCN/qFi9dcs8KESFSLL3F+zXdlRvshpWeVP53lyThiYR3cNnV
+oH8wPP6Ec251NTf9RZEJy7aSHxElrdPnX6KzduZaIaTRnUVWFxv5WegvSlbgEiH2AwMNkBGzaju
Csa4PFlmz6Igljtn9nFOCWhRyc3ztk7MPiDRSmuvHLEkSPbSCo/1l2sK8Eq0aijz019DzFtrp8H2
uuTNcOjDluDv/BSKzvHtelgg9UoP6oKYHBo14e7yRauylbLm/4xYwrSBYID7RboWWfGXidM79KdC
v8PGv5U8JsbCzr66vz9c6/soBkEi4gTAmY613GeC59VHg90gKdts0BtF+Z/ks2ylGYnj4ivkHDOk
MvWNuyohnZ2v9uwyULrr5oZ4LBsCOLYbbDGPmwZu9Y6JAufkeoO4wrFz6xCFjv2Lv+oXVs4roRPY
4muhT8i7rDBFUo0f8NIo6PhBpJjDeOpbOygv5XlwvGD0A+z9oSuobzunDBrVRAvQHhfHw2Tx+Nab
/4CQRyIwtJQ5WT3uHPLRhsg1+9lhDUS8RWOIBl/aSaltVPK50LOU9wivuPV2HTYoKEaNboAsBHir
k/Ymqi87JhoHCmPX6WvTVwzC/zrqt93BozIZHUBVY3vGPmIwe5PZMdCjfFEusU2DIZhyzbIcmHnd
t72F8OLH3gmjR4xFyWmcsGBGKN0P+h8BA/pbvDE6eRHJtUWsQne8pCtT16/G7mwPzSrc44j5dR13
kOzICMWKfnz9FbDnVtU1gqUyFVY0rTzI17FlbN3xqkMlBLxMpqW9wFWmXmjEudmMvj6Gjfci8s/Y
QDy/V53ORPepjaOnYFaOqRGt9smnJvj55dZaq5Nbuc9z7kd2sqi9P1aj7vF9s6Fc06jM5eEPjHIF
aggL+8o77g4fxcLFc0BX3fMbJBDs4RsDzBMtOp+R72enL+11yEr4jWo7zGSNyAwAUouHR3UB1R2R
IXUu3TXwHgF1EXf3FdEnu5Kc8J+rIiX720U2gPDADlB0N6p8+Lwjn+fd9lAOn4MNVPz6CzfUXod+
ASqlHl1UBwf4QrYGUkVDj0OjAGa+kfxcqpwQLZRYBhwjHYyORIVSpmlmf3bQt1uBOA9n/jJgpOD7
0BvAuXDFgTeD+ZSdUVTOdLrsR7YgfJI7vKXH9wWtX8QjTU7/gN8Tw9zH8dqN3/QStAXPoKj+CX+2
mVQR9d4QE6VwNmyiF6pLCEVDhtCmb43nBNr4RlY9U3CFjrjTQMu4RpsFirJt1bArZbLy15u8xHko
rKbCEdaK5nGsjaL0WvWpqh13b6JSqFFTzauqCFAwR52YQZUX4ovQuVtZpZlQOb8YOslnl+DY1RmR
02Zvg3hS/cVWJel8Cjv4V+L7lriIK15jeeGsY2qzrVef+stsUNUsFB7tZ4zPvtkKcYL0fXyRHoyG
Sa4syk9BVYUpVty7caSbIAU7SwDU9ndAARpEwCCvXZzUJvr8t17VAfSDHnJbxjMHK8643ycxffyr
cNTyzWtuDotibDUWXpGXLBGGApP1gdBY7VjHAt9jSIAt2DMdIq5EI3FVyoyKlNWJnSkFd5q8zyME
fV4yl8bSHBxiUdEwoTY9CB08fpPWsCxEkItEYRH7uIwknJOZticMcNQm1u9N3qiy93FzbOlJwSy6
zs4UeUZrehPHL26Mhg5PQIO1thFgGla7ch5Q25YIJFxKdrnx8ePaUTqJVlO/P4OPuulKVKcTkMju
HJiM7Yl57W4RKcsdQdA+5d8JsU+7/vBQ9Vu1I9KpdXitoK1OyZUOlihvyC9zNE5wvTFmqRgpyep1
NZw/seEqujgSRjnh8dR18zFhxDC5TbM92WNmrvmPObOvBXwSpV9IL2QwygQBArAHft+eUXU9cBao
gnEcuzRsO0/0PtQxmwroELTEJdghu8YimFh6XQ/02r7rEUOUe7TMwAQ0NGWyb0I5w7ZUedxDYHKv
blmFD3b5s8nYUq87jzd8nTvzqNaYI6v7b+Eo5oFkHeGVkh6DZ8I5hFuQL0FqZ739yS9d9/z7+5N5
wD8s7PqJahZ1WTutRuKILA7nGf2jWE1b8OIIrB46dKGFIYxOG1RGa3HWJs/RRpYVpDhxfWQBIkhp
dvbcmn9cZKkAl+RFazdTl2+ouUpYq4LcqdtaGJYuBWEqRq/KrZ8HGk8Pnwtia9W9gH1cxhJUHgeX
eNyidtV9yUP1h7xIH47SvuRs5j4xEJQzfGKlHfUqvFSu8ln5WaxskoIFfOYT9aJlTm6fuV0RRz3g
4hibqo3khxAyPmIWiM+Df91/c8NsPXqtcCzcEwp8MS31eLo+boY6NZ+1WTGKbeA9fws+t/nLAi46
EEOZGnDJudgVExPvPwKtLeHJ2loHbYH+lx6OSMO/ts0ixZsF9RzE/8Yydhu7LMidOGIEHn7s1+nb
VHQqyAQU2GmLo82bBXrRPRKHlX0K40WL9EjeInMC9cwkGq93IZArDlLJmztGeu8HSxAAjn7mrUb4
pQB1nEQQRZ0t1wWO91NecZjcsK+l8N5CCZU7Y5XFde3ofTXUb0hv7VRCMxuFMtAHYgew1CJx+hdO
kONFJfXq1EZW6tLncKJBMZHCnBv8PzKvHDySn3ZpJM9w+dHS8eHZYnpKTLhZ48SqTnPY13TPmifN
ahFLU18uHlnrTrwCs60fNuO6Qxt1SNCSKpQJLWKGdC3NXc0yZ9ua7Eu1A1kDqaq7YBM8DLEA2BMK
0u+1fN+iy7Jvdj5uFe21uMUQ6VmKv8GajbX4/oMOqMrr67EPOfau6M4lWUJFxURvTF/y5XHl8/jg
f4wV8dDvsROg1AJ30HdAkv3cuIHaDuB8JbQUjNFNBFytHq2oBEY3p8fzT4NDLPiNd4VeYSeZONez
chtC+hLIGscKvZG8E7MECFdoeFUw0kEuzKSFkF6b9KEPdoqc3cbZyE5hXV8PfKQ/wa3EjbCRr9d2
ZuwP15cWMk/3mOQu8jUDcoD1RcKYd9Wb99VFiUpI5okqAWrfRGgfaikE6dF8BXrtHG+MLkoau83Y
iy6hBl8sBhtQo1gsIhGfRS2I8jIQ8n3Fr7sbly9zZz2umFxjCY+syVNekqGVBXaOFV/vIdNdwZln
mCP4kYO7JPZmetOLiNBe9t8UOEzMz8yT3/tqX63zQ0ySLhcPQ+JtER1pkCWcBlgaKOP1VNScan3j
eQ+I2Axk+LUbzAfuSP9Xb3fSAwLzz7eaQFfPK1porh1BueHxSBG5ZhByCYHX+AB231Zs7W7K7i36
Nj0kcqkcaskruG+IWyBkE8afDINfa4liXB3TIERouoIsblmziuGnfx/j9kZNIySkq6V5vu6O18wX
1jHPtQXaV8/GfsD9HVxKHW5obWl3L68w6/xAQIPkN3Ry6l2aYbggdSs+CZjgOJyaxUWLctKXPPlU
fiefGT7ZoVQZLRu0XwakKz0I+fw52f3P5Rdw0LICMKiR1T5qLqfsqxWrhCnyTQN10YIC25LaYqOD
Feros2vG6iX/V5LpBfu2Pgb0MERrzilEnaSpm+tBNYRke1mNhJ9t0BBPhFfmNNHzPBQb0ndalBNP
r6GoFhap6zmc1+rPdvnIdBXssTh+M3PAhTPyCCW6dQhE/ZQGR+JLkpQtOI+WymE5Ff+Wd5GhuLpt
/AF4dYZ+NUSgbyPcW1MOqS+2PoE/807Oq0lPRQHDPrCrYxbFaCq2Xrgypns3wrpCyP9s+Ld7hLud
LaZ4iym4Rz+LbyZ2TkDKiYgcSZIolaUjLg84KvacNV/U8PvmWs+YdE8pJNlOZ5Cyd4Ob9Rt+3Zl2
SExBlodOSGbMnpV0lKuGrhgEKsvARzFFpzppPd72ExaGSdDn3FdccwA4l2FTsUu5CXYAXC90T7d6
MY1HeZcWUQNmY+4vK82W//r5FWhAvHdtA9S55zAlxxUwbSFyBC0okoIxBsSQ1CeTM/tc/p2DH/Fz
CRFEwpq63oDlA50Oro6Ri56+LR3fcjf/f+dTEoNUvIgIVwo6irYC2riiIILVbmeXpXPW2uY6D9wq
Hua3IeBrze5dB8V3+4Fol4LG0VZIW+5BI3sDv9VDtgz+A0flu0rLiUo/1q7CpNR6f8AKEdXLGbUC
KYpvt+ShjTbYB5QL/FzfQHANqtVrDnbUWQ1hFJMWzKty/g/yz3NQji0mF5ZEN+2sEh3p6K47MM6b
iV+yJdhYPWV+CImmGwHRXdCe7azJMbv4CEzzLgqileLo+MaIE895dnNZJ4znH0tGNzRoGVM27yT7
bQ8SQmF44CCZCIFgL9IkMkaM5LxWV8+oK4/drz/cRXpUZ/vmkIEwG6PQ1bTKoEwSbvgLKMF5MPZ1
uISSvROaruSaMUQACkh+yRUPvekMviQSRkF4waPqryBR9IyuyVqnwnBueM+r2zuxU4PX/yPG1inl
5eWKSz6X/8k/oM3kpBZFNMFByQVl/lolGEo2xLxXrKdxjZAHxDxFHyZeO/596Rnd5GvWTwMZWGLK
+C+zL5mOPz/CRFHmuQRk5pSQz/kciuhE9gR+n1c39bj1olnZMk6ZYyFvsSd6jE8gUvUVSQcc/GyC
gmFL5AJmkNveEZ1301Q64TNQhK6OOiW5U6F8sfqSAO+AfqOL+Cc3W2IzMm5af+ESDCarlNwXEq/A
LqIEUeJKXTZlCJMgUrygf5sdv/SZAUROKO2o9//KeXTmNp58IcLERtR9g5cof4QUeNKeGyLgli2f
e9MK0iMkDZhdBmj/6pFnUoLe3cvQZO7EyaG9TxATSG+6iKi2oQ2kdr6Q46fdfk5lsryXqOtOk4v1
WPkD2gMQBTZsRMMrKzT375zfVUwGGwLc1uQPR+2BMv8j9Bq+Qu9iMnwltG2kberKOSTi4/XujCcF
B+ZW/hmG9KFy9jyKJx3qdU7ZrG+8/m4ToLMJYoH4j8ZxCNGFw0n09k5WMlb2MeXYy2Jpd1zRk3xf
fZn+orvq3KEZ1IUm88g6ecqE9DL2GgV0fReqCPCbh9CdbRqv/0S7zqmrdIiSpToDD5665ygVL6aS
Ft4d2eS55dLbDaL4VBkbeORHhr3TPPxiicu9h0W0njgcDEHCa0DeufaiD1DrPZU/bOAr+sSHzcfX
U9JSJoMJn2/ttk2zobAT3dHvSelA9EHOJJp3es7Lq9D/FlEJc9jej6p+ZeY8cp2pWAT+a5ks7pmW
YgzCD1PojHPDWT1P7HyTIpJs7z6hfAJvuvY1kIcD9gyQIGCIvtzBzUdwfQIs5PzF+oWSFtMiCGZE
eY77GnQP+x2+10HiuxoVeYEYpehBnu3vzAWBLbnYe+RpuD69mI0ILq8n0T2PSqTTg7F9MorBxLJu
+wz1+zRrzv7DqL4wVRCmzcM95XBP/E0AeBgu4QuY0gXoQFBDvwBnTVBDGfqJ09I1TIu+nTRTOIb9
avaZqFETr9RvVSxJsB8714WgmM+CwF5temcH0jaLXjySFrgpi4Ua6p2BTP4ONO1TYW2NbZgOc1Ji
/YHssuMBtFMwsae1kzaQ8YubD6gB7mhn/BEnQb5zvguj7Z7AZWwXyjHUMoBDMOPLhyyhmFyTo74/
lMBhPlgViVdoURTFFODwtYYZTvlhl3HdPM5CW8JAb9lbnfG7yaTjR2d7N9SQpba1rWkvAhz+l5pr
YkgcKgRrmbXKolatCuHQiGETeDqqXQn6fT0Vl6G6s+7Esskr0Ci571aKDT0vhpI7vc8Caly6Yi3b
SIYQv6MFynmr1qvTtTQs/hrkOSwWBJS59o16cEdVXh+j6xBZh9qgTzynrkbeZXylIJqVEVPzvZpY
+u94EEW89dclRNb3QXmKJzCVYDAdE2gXNphov0LeJxqgLcSCNty5Sohb7EkQpYT2TrySfmNOY2sY
HAeOeHyOpgi2eFdTVYtF25LQb0bgJaYE4roS25bUIidTq+DO5dSumWpcPfEJkfMhMGfRRPcQWLJI
EK+1pRxWzyr1Fz2JGC++5QX2GEf0zdD4UKAGcT17X9LV7Vro/jwKXz8UKZf2IFQFJDeA8//J+Pdg
7Zz0htCkUwmLSnH0M78H04DCg0r2JcmEfv0luuRgA8zvbaF4L9qdXTs5qcyvd34nsaLPxm9VSaYt
4CEE0ky4L4MptLJHJLm1GVwidi+reiLAiyrgo+dFbnYtN2wJz4Zl/RmEswgM0q+B+dz/198FKC1B
2XHiNi5ly0E3MsG8k6KX6TrXonzYyx9v9f33vpfSoS2l4VL010dYbO6vI+pRqeE4nQu6U09lvaTt
B5DiJ8cz0InQ55YiTYf+AmBIGt1ckxSUpWLeiW+IgDeMIDlVuIgV5s3lI8sFXlEJ4oaV8EIVaK87
43gcNDxgP0Vvy1HvjuBIIor8C0vt7yaEnR2iZhCzG+p06E92GWQTp3F9u2+Kfq2GmgS+u4IF4DFZ
AaNWRQu0nyt4UnwgT9FzPGk20fH2onRmCYr/B7hDPpXR5YNykyboYuJv5bFbE6QTPDn/Cj1S0z3R
E8XsKRj1C4D/8Y0QmAyU5jEzhgZhd/ncZvjz3Ejco7MaVC8q1Yjm2022w5r6yUOAGsofBWOqWhAK
elYkBYgCcToSUxzmIzmLdferU5HwQmuiValon8Uh3BK5Zh6MdC08MwsMeRZFsYDrix48uNcsKkmS
ICgSHSG0iFTgSE2eW21LznWpCZJKfM5NXLFEPKvubgeG/48Ck7HCACur0YnTMTwHbc9Xor5iHVsM
lbAYULazBA879YNiKgUJBHRrY3vx/l0VSnbiRa1MdhEyS3NaA0VWm39VtmdjWHE/yx7rqY/qG+T7
euNvR6Za7f48hvjRCg1ToQ6lYf72jZmq0o6NENgPLTlNJIt4YdHRmrQHLFa0BykU2AWdBfbX0c43
30ycJT/SQWWUE9FSgFmI5dq5c1Wa88RoGr+RAvnPsqfhcbYJAA+lYy3+K5nbLSBY8IhGHwmIxmPv
zO8nlcN5WFgngSHY+oTtGjHwkBcVgqZn+SnF+F6mskIWf01AybRkrahMVZdrLD2E92qmjwzAnlo1
AhMUGTIs3UUoJ8vPa4DUAF0qs5xgo+ALj4ek17r/uYzSZBCDUGygnmzdmhzwaO9xYgjKc0vn+OQi
5KA/5s2vXiRdALwGJdRmeCYIOrSWMK2Vxzh/WAT3q35j9Yg0G3E04o4DKSoKh7ncybQ+wpjdq6e8
7KOG94bXBh9wUF7iaetkb3fqlt75xWA1GXxG1zkQzmks9/IAauHwkSPzrqnUxGWDZ7W41LxiY5Tz
gm96L9lJbRc9loDdYyOwnvxrK0Bt2S9yxYuMuAQZzvrUs69zDSR/EYAbUTFtyElCxoEtnfYqzmXN
dv/co3nDYN8olvOLWdAnctMXlFO6J5ioseRvTVSu3+zCcJbxl4XnKw/sl6m6547JL7yFWqxwoesI
0+nUNKZ0U/JMw1ILFTymGAWI8atzN/VSAYoMywD0vdfwrVAoe1PN/ZS17h3+NcqxRUV8pqN0hhbE
i7/U+LtLbU7VbOcoC7qUUWve3MP7LIPES0Pq7zHFrH9QiZUBeg9ejIeOCL76/v+oasnJRTbWnNMW
DzhmW6P63gBrrJYT6EIAIc21uhsDqMp0f9BrgPc5r3xjFLy5HCqpqJ/QNKgD8QELJgLkFkXUcmd+
e7XDRMHSGnFkt4EiCMY2si9GOoNwFPWSi5YLjEhiuHxHPNNFLOqPxxzvBLlZChx2rIhcUWZFOS5e
3ZT/whYGlffKl7uA+gZfE/UWChyMMt2J+qQlyrzgMitrkNuDqQlB1bvDFgV7s0pnwOoZDaKllJJq
cSW7snQXStgZc23FWru9ytG6uEm9ITCrAQF+CwD3lwHLJbpYnb+Lj39LJrlsAgiy/8Gyl5MDbB6b
98GeBwkeqOatkyrxQCMREkDTGJhoa3dClgaAYqSt3sSPgxtkhzWSlGt2jW+hUIjqMx4FS2sNczqp
bcbirK721g1OavcuXHiFKMsSgWqNpn7gaZ41s1uqfVy0Y7M5V/UIv3h1trzj31LD7qXiz/lHQNON
fyOSjTYrUyg+UpX1OP4j9oCzr9LoeqdquKDpEiqQjT/ZD0T7zPhIvMfAJNrCnB1xKim6hrnnu/C0
gZdXbBmHaGmlJKDcb/0DhRoAJA83moixr8TD2uLdf9QpluOl61s2GxZTTbG2CDVJxJ4E4pLrS5vC
TPMsF7Zmt+O8umUuwAppyQvaPZOmDS5BBqR7WJBAW3/pQG9wIiHD6sCJcjIwZn0LLx+474Fylqax
TXpOEtb6m4o96K+4yjhLKKgWd1jNN2mWzmiYgRdp7yqNG+CG+zrBFgiKcV9cPa6B90pZXDwVebZf
2kt4rqtMWG4bZ0OulWHrrMyVfy5DZqS5zJnfMknOg2Td3rL+uUoc62jXDOnrM3YloUS/mudw4MNJ
ns/riEq3tWWY54uwmPJMHgfdyo+rYZflbQe/RTfJvgnMwyuCkBaD+MTZcM1qI4V9Jiur7RMhVxxc
i7MY3G6xW/TX6ehmLtU4zhDv6MHj+6BdPIw0F90Ufi2mKHpYWfKrtnd/Gw3onEMQI+AnACFkFmUo
DY09wiBR7sO10PZBbeMujlcVnMOGIgJ4Riz9pbs9GhQjjw9GSCLRSj2rTrVPSZC14dgLJNLscZEv
TpewltaQpsCLd2VNVuVN0V9H7tAfuAD5Gc/QcdmXt0c2J8AlE96oAIfikLOW/x66Smqy/GOZ4Bx7
Ip42YNk2tHdtaJn4BMw6wbzGxNB0Cj6zPakE2f/DQR+g5VXaMDQ/dpWp7RkiQrWt+ISPAVWqS73t
2V+eityBwGqd4AAvfx2t+G3NTX7aXuNdWHOv+QNUH6qlSRbwIHw7HAeDmmmP4z/7Wa/hzux9qexg
Xd5W4h0NtIaSqZaLBcdVcnLspG2Eby+qAZwN2vgMArFDidDd+35W8aWLR07x8M+qVqJqDVb8NUAo
uk4PjLh1j7y23iqwYQb5cjehiY74rO+AcxdRSNTnys6MKaQ9mfBzumKvsW155YFs75ja9hqRxXeN
WDrk75tccmuv1bNmQv7gJ+Gbz/EdomYLPegdN2gssgfVryMgpoMpa0DfSfyNa6mQz3CsBnkv1IoJ
McIYvgUkujjDrzU+6/MxxWCIlrFXQNHvjdwdxaexSYzaYzglgzg16XDSVOUnF58a+Zh/RsbPHCkK
tFf4cRD5DNuh2K19xMN5OXl4f6v+Z+47HDHmNSQJDRp58VICpcVOCksFO5des0/E4L2PDp48EIwh
N4PEcfgbzCFEZ+bfThivpsTIVHiWQeD6bmpgM5ZpUlYrzwFcoI5zGxTnsTWdMTVKW5tMngnO6tW7
UanbOPZ7ea7AkeqvTnEOrxxS42ZfAaH234mFs5GjYvw+mj5rxNyB7Jp4zHMMPzzgFFgBFdAnYE+A
cWWcD9F4FMwJ9oNiJFq883QaYVWcMQL4rOd2GMWAIpfHt4/Xelq91GtF47hK5KiimQnLYVhlE28i
DRIFzPrQZGUOOdtAZp+NAEUVrcd6Rh3Nsyz6bq1ATnWwtJHaYYC3frZZsv+KW6R2dDfzyYRXPIfU
qOnAsAxrGndKJa6jKwVOw/oMMMtf/58b1+2dB9vfUK0FiatvtVuAMXytmAWXlAZjg9IqMGoo40aJ
N1lWsbz8A9vk4U4vNXm8hREhIZX5VPQRmYa4oImP/HscocFdhITDAom5En+dUGqjrpgvCksAkZL/
FQqt8h3RumpKEk+bovyBXrN2+KDnzh2qagrBcBXTK+NtPW2XVhh2k9Bq9S9YFJWJEH15gXrErtxU
t4JAyyciPVya/SRd1e4zbmJ76A6/z/UrmLP+Z3uf2VEiTGCjh+VGSwS5U8GvaOLR5wFkvAdyOfF7
z/sN4YRoUNArwDn0nugI69aSr+l195PGALiEzXTifWwnyONsVxbDCEG/dh1nHotGTVqpd1R9MYGK
Yx21rVtcpttYPZgwcUCf357BVSRT5h1/QWvF7C/MjgoQKmIQ3JE8ZXtU6svTbl9xqwEd0cdzUjn+
2jPqtO3XX6uQ/aFbQ4BfENVnTVB9YLaeM6jhNXoZyeOHTbQkYAZEI6rz8yTFmXFIvZCWaAcht8EK
BIjk8muP6G0dIEfIHZsIEXq/zZQ4aKjFxcdnXnj2M2bK1siOQrWKD3S0cZtn7G1yuTzNtLsGvnzW
V+/z9yTq4gl4V/FYiNXfxKJKXtHujgcLbrX1YD3HYNCARvQyxFp6W1e3faj0Ll65YK4seJU4sbIa
4ESOzqwoH3smFLmxapsOF9iAaPX13YnCTakfxKZwhSu/HHH8BD/tl9Q55i6URZydo1eWV6pnyCuk
K9Oz6hyCZr3zh6udMl/F/4ZGpUkfDuqIxcHW0vtZ1qeSspQP/mNzn4FBC20qawZ/lwIR8ZJ3Z7xT
8vzTDGDX6Z/jWz8TuS5TNELaJtovumeEcYT3BvVGVGmuRMORWDvvzObRBsfpiRZcH+r+8A/Zj05w
Z8N1rtMJ4Se37O4XGA81BA9VDKJfJpK110WFNdoVsFaGpSieNO2rVJAATh01vl5d7K19bzmBnqaE
ibxWskADi601jn9V+oYPyVHN9GQ68XwZsLYFMyZ8T01dw+J6Fl61duWn9BLykcxDmkCwK3XBvZ1r
EP66vCxK9U/KF4cnANCCXKfw5ztI4eOS/sBEWJqxHFP6imWgF0YcTu7N1ytwFLCagQqd67lvYHpw
A8ahPR4LYGQy/bR9iXFmYB1hLoWxqLHLwnqczXMTtmVOnoTY/c/3J9glKiVes8UwJS4JKMP9f6V3
kkI4ycWQOgWERRz5Upocl/ALhStAllvAfs6uYbFQKc64wWtImPvjkgiiBB8cWFYvpUEIr33vwm8Z
HyYCpribLYEY4192JnZ+WAKiV4en88laq0BoQ0mN/EeciimlScp51ei4oiy/MxAkdJqu/QtvDDZu
v2MIQ56h3+CSDU1amsuRvYocxHOcMB+Kl0zhr5TPkHJ+0N+wkP9aF/MXh+rqg4Ueqz8/WY88cW9W
k4SlZ1bvs+6Te6qOKVN56dXK+A/TE48YOWiD4qpBULZvaHTx64FKerzNG1UBXpp6PGzcZDSdNT2I
AoSLNMiLpveKoi/cYRBfRXaymZkpcFa3vGEPgsaPDGoi4EcRcgR14zTQSLZ4erWcu91S+O5vnK2c
RuSAubkND7+orLntBLwj1EjMfZsdwSRgxglCujkvDBdVNta3XrZd+PzSoiwC0DCZak6itr55K4sZ
VY/9zL1hGilcqNcZF4hJkKaoXMkK/00Gozk+QoZUpy4hY27PPcvVTHMgrzX2Ghmx04/jbOlj+l3N
6grvlb5jM43NSZ4IEHzzxRdIj2nSh6I9U6ptcPBRKkikhUkXI2I0F/q0XohptV1KZYXQi3Eg4UCc
/ej9TYUWqaYWOw1SWWrIDYF7oWxHxlOf4h15Z7p4LkM1LsYmscS1KdSP6WC9otqXwkhz3jK3HLy/
mxry3362zTgMwKzE+v+HY5Bsx6hsWeVNgk0l+LYx687yv6TuQSLg7HgrC62C3NjRutVJksiQLdgk
Hl7MbCaInO2lp/Y8c9PgRw6jYmnGbMRKM+MFqs3o19lR3ucLkHsdS4+wtzhYukmA4EyYFjVrO3vF
Bv8vbtfz03fGR3Fk9eAyDvlzmeBlSkHnr5MgHh4flBxTVggQmcq3RrVJbJkf2k+52MjXzw/mMn8e
zVDr7VekWkLDkdXc2U1RFTCgL/ATMK3iUPKGtSvZyilw0m0YLsUmGAh1rHYNwewlo3hjZ9n8fRjF
RwaPDoHMOfvBeOm3Juu8Ar6O2g+2gRnO0gEhfTaBIqZ34MBK/Z3UJKRw7IoaxQKkidY+z58Nxta4
HPl3TYlTHrSd0N+6iiZQ/iGinwVMMQYo/Ki0oNRdIYpSYiXlIQxAYRo8wXi4baxMQy8e4q80r5yT
faNDI4DEZbzzvCuLuKVL+5ANJzAqh54vQgb7KrvBq8eDf1PCTGtrm5mzh7G4XL5s4H7lfWdEDNGu
a9pM1U6uf9eCxkO/Gc4OimPZY9KxkA1CyEPvA/NgygW/eh/Kd8s4r+NKC6Z6fbKy894BPDtj7HUD
5+YRrzjefhtAB4x6rnlzpDmVdhAUOkzZoshEDN3ookkcHtpydq/B+Fvv1SxRJEm6uL0gfbha7r5y
VcuVa4BzDP/toP+gDe0AA3JYPHw/HJhegTF5+MZ8smm/GODa4HNj9JcnIE87Wv1jwlSRfy6UoJZT
FDBOBGL21QsGIJc2CmH/GkEq+rcHo3WdnEPGZG/sQzw+FIwIDIXtKCjyf4unwkG7I8k3ZtG6zlkC
2uUPlxlNYFg7c+7i3Oxx8MY0ETi0Jh0dNnTTcL2r1GL5a+5OgX7jTpvVtMRFPW9F3pP5rVgATuXg
YmaeVknpjv7PnWg9nWwRl84E3iBrUb1P4OGVcbyYa1rI/UXb6WF6Hcxo5wowY87QcEAIlCG3IJg0
SNXKUqCGUOILTOIIvaimH0obE1VYpEBKpRpBxL5csyxKIhgZOJFzz3wdzofA/vn9+UEuri4z6SGF
Ed1dEZV4NkJlQOxzqPao4kw3QWgN9ZCl6EMcOV8CLjMDNjb/9p9nPNDAJlOYvmEff48LJrgw39Tb
piBX/23Ey7ZYvOK5fGB5kgzp00dm+hOkbNlRJoz0sXoVeq2Nsg7Gxw0OtFrVv6aREMxQN/cx0qmr
cC0NmdvARI6OkKo4Dq2lBjKu/Fz1hGvl3fFGCvoS+Ygo8ysVemetSLLV/cyH5ksxfNLrQCXipSPT
AE9vOAa8ksG2lz1j8uHCrnw1YIPZCsXFshRQb1r+X/M1y+YMxPdlcPastg1ryQZfmlCsvALa0Peo
rwW8nSiebNThjct2GtoVtC+nrWPTrADrb5/lUkRbJZ572GuyFZ04CN5hjVqQnOIr98xfH4f36JbW
pmNqGKo4CLLPLxJJSvurFocGHAYxxmG8zhYY5rWUg84IxK9xQgK+zQF9NVJd9z5/4amCQPTuiRol
XiHWDAfcSzXbOAo3iF7FdO/Yq+I/x5Ds25mVU0tt1qHrIemR9P7VJWsrMnS0YrWWw6jxbP/1weTi
qEUXJwyHYsXrIQOoPBSqTZkLm+ILHZKbh3dED9W9rC3pFO42MGJqGdu8tOx20CmkXX5DDjwLkafg
CpqxZSgjr2LHzfIjaWReBSBSAkJqarB5NuMzds+0XU2rzpvL0u6wUetchYIlhBsU8Kag2W/EWnDF
UohyYOxwoL13aeoIep0GfFYsljmDJnSbmaQly28LBIRfZt6DpHhJhMcgG7xXnX5c6LCyQXPtVKuc
a46a3ddXaXJyn8si306UxXoa/BEcjpa6QINqhd6HebSDUinyo369LmtKqGy8JdefFg7OfAy+E0kZ
goSmr1iWiRoIWroladsVYco4hpGNxtM5xqBWvBYAFd7kE/uzWdx2I+X9cyUrkOj6I5F86J+PgHVQ
HTupAWy1BGwOlxAMiHDD03x85CYuQlmhShpVkAqN1AaD2fKLSEbNoAvgl/m3VGUZ8hQU5VG9uL6e
thel0y4FIKJ/SfZuJQIJcFpmBbIkuKmMwNUo3xtV8QKSAbSnT6T1jBAysU/p8ams2Qc0FKjoU6+C
/p3Rk9KCAe4+1fusFZv6IuaJZ0E32zUGzdwW6XHYgnbqR9950XtQerFrU88z3RAj+krbcUFUDKPT
4/uuzn2e84UoISo9uVwZZR35odhzsLP27TfSkqjPuIhyUrCfORSvZZZMFpHfit7fAFxpWKcal9p0
eDcgCVeh+7PAQE8u8tRNGrwqkvakYSOrv+wt2oQxwKAcYqOBX3xFLCY48qYgpkcfT/4/Xeq/CHx8
vkTZsmartsLjCOnXbfVSVsPHQM/600HKalG7nGHhOvz59/3nByehm3UGkRDr94APTyIuyU9maIoZ
lulM+C5wamd3rsGvrmXf0Hp7f8teQLEhh0bBWyOMb5WyQPmjKvJoMB4P09xBT4D395P68Gq4jMoL
1rrSOg5JihUaUyjjATiUksMsZxi8k+81p54xn+iksnH7PZ3gxKZ/3g+Wkgroj2mjyP1Ucc+YTDcv
wdkQL3IGTxJv1IGjTrW3a5R+VRF7VEU5hBXUcCYr4jik9exBbL5ylASPapy9ItEkIBtq12dJK4QA
xWjtmAgWbP9LrlTXM1VLAW8EaYetx2uFWRZ9+1qWz6HQn0qB0LjiH5sZJ2k1lyo/uGd7yn3M6sTE
DtYvLv4tbaB0Xos27SMZ/ueIEYDQyuEMXy+DOy3q0uQpsyK46cXJ1uMsUphaFFZzYuOtxI6ACO1X
N+cX3aPf99YkeVUNd2BlWwPBabvvwQ3Z3whXlGbQWpog4hPmIFnknK0naGivfaa2pagIDUWt/H8W
PSp42lm0QVA5zChszgAuoYxO/loJBRJkz813hlng9iuiFyAjCpukCoQu2abhhy6mej5CqnCiNMe8
aon7H4ewYPUOhUUz+t4BnP4+9S/H7euGKsqykZ6wJScEChGpYoEBXdfm7XiwQZ+zVnQwco1CDDq4
iR+HaHfP9cyZT9zA0TEaoXjOYYqKwSfAAB7sfwmLMKu7W1JJTGimcX8AqM2ad1fYXr2ths0D83Z/
jpNcivu8WfNpXLpBRZqTT4L/CjTKWHwZ7yOryz7EU4EUP/C9v798/cxAFANjz3jqPD+IBCwT2Sjs
RNvVrvpWEUdrdfp+VELmo1R0c/r6j7eA/1gORAJutgHTZt8jnAA7PvDB9wqK6VLbmwiwfaHQkFyr
bdVM5g16uaNqk+VlHOPCa34NXrN/FEJ5qn1DP918DwEOleRQlYDY3BFMIBhFjbFH1wxXEnEY72ob
ereXvceEb5O403GWr1CrKE6R+G3Zh30yAVs/VQ9hLXRLe5mfeMA/c0JrnvGa5eQJ2n9G8b/msX4k
tH2eWu5aUQeBKxqpWPcKPjW7P7nrEkTQcf50G5U4embenpJFZH6TwrD9mQ3qgt3u9GRvpzMjVkR4
a8TbtproaG1k/rDv0QpJvec6lwJHLzMGoWVgFaK8XMdC+XOL28Lm6Y6umkx/GseENJZQmGfL73mZ
mbWlm9QE3+XuNMFUUYLQGxKFBhCuJCwG6KnWj07OaKRf/5T6kQMY2xfOH1peoFjjEmP/mbUpvNBR
GiKwcJOIElkMuCusFoiqj6uLzB2t9oLq8BWn0v+d+OC8OiTXczwmrCjWhOH/BAVjhKy+RSkAhf7J
MTKtufEq/srqHRjr068E+kP9erUeo9LU0vrRaUSQD3gsTHP2/OUmD76u2p59kgXfHG3KV+x0cdYz
WSsy0ygo2C1qHbwOWe5fXLCyuACSaDxGTQt3MFvOjOWn0M6KsvFFYvUyApIx3DDyUzys3hylbiN5
fsSsHj26Xi3qxXJj+T7uKmvG5fwCd6PePSxehqbWMQMNz99brcP+bJndTBS+2lYTZLAxKFS3UG2G
YwdAc3UHe0a8Cj4W2vlHm/MENFICEXUD6vgGfVOC6sfd26gtgr4cpxXkTiLMGk1xdrZzaV0Y/mRd
RqF40SfiKtT2q1Ox5hIz1YF4Fw387Qx4TvR9FiI+iE4YlkGwkoEOFRz27Dv7TAO8lbWU9gQYKa3G
nJ+lqNKEnqpKYbIInT6FCbNrtBNm3BqmckFxF7Ae7zbh6GUxiHvgZ+XUEKBDbaTOCOprjFQSTM6W
5rHv5aRGenC5N/Va0fumX0BlzXuGoOZTo0D9hjOnLopzfeWOywjG55slnrkzHAnyCbks7kYESkNZ
Tu84YzrWy7q+l/iFXb+hfEN+QoozwsF95cNOc6kBc/lvUj7D9hyJJNEFSDVG+HmMXnGtnwyj7hy4
vDhkLSPFEgn1e9xBrFsubPli558lisP7elHDxwgXypKEeDsxxcfg1S/iBOGGI5V0gfBO+PYvX0GC
1c/sRLwqDYWwXQWcn/RWxrXMxKLKzhrVzwBe331B2fjKE2PWthQGlrZPD3mS8RtdMS7iocvvsaAp
FS/4Fxt8g7FbPNfnruGIzzKaUCxGWAazrTncjbFE9Cl2cGO1TgIKevxourLfa5DLxpLeeU2lwD7A
Cd2gcZg9LPaGzWOBxJq+GigupDS2qMjJqBd30X+ZgA9pMDblQqTc0FTJZs029V7K1W7xzVkHkWW/
7H3NJJyq5EwfC8gavpt/PjO1PL+NtrP/7+M7qLFvEeqbBY4GhNdFiefMrla3N5yTyQPU8rTRug96
JOBEKXW913qVw9B1DncGNXUb2O6NKDbVpU7WDN4Jc8p9GLAS+fV3mMuk+oS6CewQsVcPea/QcD3R
xmcRgalntIjillPsCkU4U+S/wOvLflVBWEZP2CkCHgwQFRj4xMNwCqspKEnqx931vzWbFfXJ7Tdd
X3mOWCfoWbk7dd/8sOFswM279m0ckbVrurHKIRFJjGx32Fkc8xQaPXVvPuGNYa1sEtCaMy5G7/TX
va5BCL1Gpk4T1V3PFOXPc7mFBBHPENGgtzKPXKmQzbs59lpwPY3UOxKlZ6+0U47GFwtR4PWV+Yk9
WFGQAsm87yjCHwEvOCapoHKBo+yDBpT0DP05i9tkz5K2GZ2bKbwyLjghxTCLEkWj0xr7kHMZPWoU
36/fYd/j73ej1jZDoTI15YQz/hrYYLYz9MEtRFiIK7l6HplwStcYpiVmdZSD5I9EFRcHmPPSc9gA
zhkM5KoLQEEc5XQaE8Fx3AYVJRYzeZPfNbpxXh8v+UmJqjXoFKUrGXk1H/kESmHGepfXp8eV97sg
OZ/C9ApHMvFcmxPQ00W6KBiBysdxdIutCaW1Me24L0/yVkWB20hBR0sVr4XqGc2VFEY8V4e0T0uk
CxO/X7JVh78EPE2SyVDRtT5KKaHi5nOEXj/1LNTwmDH0MRcHlDxfNu0sEjrL2KGp6/GRchx7HliK
8cEaS4dsQyaOEZeV9ZI5ii6+DAlrwWQcfAOD2Kd3u5QQJMTtuOjqrRWB9vzxc5zI89Yrofml81oe
eJBUa1zmb8aF3YPuTQwUXsFJGJ7fqS/LFgTnfcRT4I/4kMvaiDvegZ6cCpfkVoH5WUOa0msazHND
mPiRwJIjDPJhFOlFxnYcZbwbeJQ2VyY0bPR0wvFtlNKmYVb2SWFDHt799s0sSSdwzfbQtLUOrvtH
+V55ZiK60ARnxDJEG7afvMvdXNyTYfAokiibGlKb55nSSXrcybhHZhL2FcBsvOoTgxeabQYDFgOn
uPBLhqu43HUxRChncZd9F2Fvy2g8isDhNrApkPSWmTx/COgUHttawntu9s6lrBfd+NcPMVa2BRoY
qggsU0+e8IkqSMuB+7uZRDmM1Fw4+9aNIFuYc5mJHqF7QA4Jcg/7Wa/YJHpq8mEe06VtnSRyTjn6
Vkzz6ksNXWkKAFI84JL4n7VP5KLQS1Jwl2TnaTD9+2h+B54t/3bIeZ82tTmQnptDUDiKVJCXAVfL
/OAU2dS3wsx4rKpnA+gd+FFN8n2APBxuW7xbicFIQnf2OHHMA0DrPJDPVMIizal//diUfMaVRKjV
ddeAwfAounLurwcyFBM+YAgsC21ZryjAGxkGRK1sHlche8yCN1qr5mgPKcA98jLaxA2T9Sq1h6Vf
fvIpnGhFHTm6Ct5Ohn6gMatrToTqQX0aN4lK6Jh3Jq/DuesjqvZZDj0fX5XYak9gkMJb9cxeVZ9V
eJ83C0nl3nrcuRxRSPBVQ0hyEfGiVC6hcuNWqd0DghDUOusJMlZTcIRJsNY74fxYpP06eN2LZiaD
6DsRi5PD8KpjWOmyTnHyfFwp5bYr10IKOVacg67uj5FTTb74CbRlf8vF6Hcfa62BfqtuCFMlpwnx
xhpLE+a21Rq6SpGjDdyjQukfmkbh7Mq0lSK11be7UwumCHd8I8exLezSxqy7AX4m9moS2uMaYNoz
/rx1fcOlSvpYoeGyJ+MlIWrqpznWU10kpPvV1d6hyol+U2TRlimNG9FSmhkv0Rx2d9fuGrxAScEb
4At08+JoiMkFG2FUFjK6756xhYGNF1GNZPAFhbjvnMAJYbTmdvWpNtUFzVuArJB7Vhs4Jn4UikNH
0HeKPRMGPRqp3q4V52snXD+ZqOlzL8cV6/eHpz5l+Ag/t9w+Qbq3rFaBqjIMKSTGCmA4rvq2UtFt
pLJijpJ904QlVxBXTHJ+szt20XecnDT7uTIbjqwkZ002+lALIf6+9sRdSnxCsIocTgrT5YB++f2E
2grHZOUI8xvryk0yZXPrgvYyz7URjyZ6bOZs6T2fbvDqJIS2nkaRbViK4qWkq5s3b/ES7fOw1AsT
YuPY3JzN4bKKRZpCooLcMmc1uWGiz8SB1CTVeHiOMaaXmJdqdVlO2NBos4CIs5zvaKyNjBSsq1FN
NqpO0JFwFxcB9hi6+dd8ERQNjTBTufsfLsfoDTGc5fp2MWckgFc7Vvl7o09+eOBSV4TbtFNnrVZK
EgamgsKDjJTM9jYKp97lOcNURffRiBNKYP9iRb8l5dGE2y/WAY4+eMO4RTkaRlk3AWz6L9BW67nD
6sab8HbUqjQRtvk9PrRxmzGbfeLdIQMlB8T8ok94I1R83xA3+2t1x8ZUAFdxDTkTjkPZSMhbJErN
Ijg8b5oSL5jEz6eKLOh77mfDn0Je2IgmUs72diyxU5UCpplpYTWKJfCaggx/FA6O6vWLU//rtW6f
0CjU6YXix8mSThtACaOh+r0FCCMZNo5wRhG5gsODVzrAZyFmYBJkxl5piA/B+DpuWD1exOQgohCR
1SjeZhL/C9Mnmieo7w4wH/xPsp66d7NifLgrExvMrcuqX1bVFW4FXdumeC8U7LyEiTG//uA9UMyQ
0awgkdI2oVv98vMNF8xkt+8ukjsv/j5dT7/YQXcLEqf6tu8NtauIo53LGZYpXrR2xkOhk2rQJGv0
fHRMKwxvpBw+oaCLPwdA8eFWtttl0iJdqyeybDaEjPHR4orWXix8+Y4CBvYqFVT0Q36wENCuTftC
+qZ21yTauKY5PylrhxjPtdUt2kaK07Xu5mjYjPptX+q3oqBtVuOkQHQyWHqzKu+zQYnCxK4sghWs
4MfTkAsscSb2smbaK3mZ2plZ+usRbk+uHyz7DuEi0LGvqXPfdsqQxCCoHwmb8/sNw2M+i3Fp59gk
0P91qKCRqC2Traczx3Jwu/4ONKkco9fgTrS6qtA4O0iljLbfc+uu3i94bt4wRXkQGRmCBwPJ9BW0
ScUN+5faMl1IWDmvoWG4fJf3OWGo2UJYrGb4gY2hNLqjHKMCtbzxIrhPEIZMAa7uba+T382Vdt8i
4Iy+pXe9iBoMA9rcC2Hgy/GPx0YSYeWQg2l6fgOyN3gqTWOdGN096BQIIVcI5F5GbYTUxDFQpr8W
z5bjwDl6wYyLh12KNxnn+KDaINXsRd0sMtd8BiwW+XRXwWcOSW2/wU/2SxbSfbz3sSqWbHxb+3Yo
GhUXI1Y2l+jFDrvzPa6AM3Y5wl2RkVQHpKW5cmbdPMusN6jLlU8MsxJ9l29NbJ9Dge3ps65DvZPv
ZWQWWc88PLTcWvZnI6Z2NCWsIZhxFv4VpFbImvg7hpAtUwZbQHqk6TACsIgLzeNiMR/A1KCstz9B
8zvCJF6Ksnymew2iT/sFXeUhg7uhuzIQBfTptwXkUn+DL37PBDlq735JX9iM1VoR/0hgqztXnTod
rsJrwYdeT+XpjzS7QRUwtFfnpcwSACGqeyAQoq1ZbpAkU000T0DaaM0kgIN5ij58nEx1pTtitl+E
3PtgS79KFtBnLMQyfMkQ24JpWVuw/IHpMbyl874/2COAPutorKX7rYY1SgllLSBFQloHVCnlzrVM
nFCYlAZPdE/ZELUHH9OymT6+MbD0s8EpxWy153LOIu0oM5FVwLEh1Mi11CcGsU+czYVYQmpMBStO
/8O2GVYZD2f4P/lBNMtsftABjq5aWeRbZb3BDuJo0GG5urd38DONRJZXZjet5ituCrUMIcS+W1EO
QZdYpksrxxiElY6twxxTs7OEEbCrUc4OmVwDRkjCiqdxBgn2zfqYzblYwjSH/W+z7jvwWdwJxmiz
Czgz2bSdzEGnCsxS/0K0ZWZWi40pp1gBPl4JrleeB1s2eVMeUCeZskv5/a0bRpRg4YiwgSV6F7iw
K065EQDQRJIiSr0042B74xtdUFPymwOvUzAcXvKZYa6+ybn1wOFoEQTk6YXnOAiZZtJXlYTpwsZd
qFT8ZRXk8cwSYzryiJgXjY2dmB3t1+HrKN6pRPSGMaIX0jSNq8wzmI5dwgByF+zeqCqKqOPQCrLN
YfnwvuCDdOUTnf6SZJE1BFlHq+IMdScPoQkCpASGvLLlTT4ZrdUEd4wQ453zng+vs19/zlSsdgjQ
mh4uk2br0+mYtbcj+2HSMSKhBiF9FAPsTJ90BLPLbyzUsV6hB/e4zDTNoLxIi11EK8hvqmP8jAPP
pF4CBb8iJk76Z0c7mqZRjwD8o8YUb+QEukaKSUqeGBJDh6y0GAY4lLK8k27grRIdJCeznMu643/O
HtidsozuyDR5FxJhtDSKUljW+yp+IMiNhEYsF8DbRQG014zP+uITcrFRYuzU65lbLQUO9ObgAyMB
Y947vLiwUbzFSVNOYiInAX6C8J1xxSAq3t+Y3ZU15kTKGlOFKiE/rCUhj6vzrDusLcFJUjxrAn8X
wqG9v8Fz9jCIiPeDDogu197FmVysD5zqB2JDW371aEq5wZugV4E47a+d1FK2XY9JL3T+ffYZTjz0
+qyebg85jeU1sNQz9iEZDFEGkv51rakdvpSHlyAnUiyWKKINNnY6A3fcx0UNehQdFRHFDtpT7KBN
VMwBiUY0t23wD38oikMxtBCcovKGl0vE5Qmj02+tN4jR1cow1KEmg4aqM3TJR2hS8DXZ3uo5UzQo
mmTnMgfm/bSdS5v2eudA2A0XytzKQ0LCpbO9xi8lrxwYdoQEE5RbO5rDH5USBSOiioycrqOeEG5N
eLczWfxX2nitOpdOtc4PCSm5UaWXuMrsnk082c5d9BIwscxyzNPDr3QAJcz9vS9B2ygEvgmINPR8
x8Iym71WHYUzsPuT1mKSmPMKLz7gUEF6kMRFNZRwKvhHGlKA8cgqd6hgrDdlkcwOwdFgVUvZoSsJ
OuRE22X7w96TxYd/gAUSg4CQlkAYzoN78abdTpLmFQf4upPhniBwOPB3UtQgbXZCCUCiIhVoqOnR
oY3JSFrHm/+pU8f+i5WAlnNOuVw7dSpNuwPOx3GsXf1YuORobzIilisxVx4mCsd005KW3YfjjnBm
SAWrvi852Idm/dxOdEY6OeeCDsp26VwGsvfF7IivNokluERYd4R/IHoXGytcadES0DcQxAVQdLda
aJgUHmDMpE/6freVrmouxOdAri2J8KneyvAUJVRK4utj+w8LKZxxud1X3VekryG49FN7nYeQwH5M
MIdDFnh56zMsKlws05cIGQtPjhgOV1LrG12+Ktu5Puy1sDMCj5NQ4/FQarGC+DePPGGqDdgg0SFE
eBErKKo35CcnqU4RDaSpy+q5uwYtKJkJYDCJODh8z3ATQNQRG2a9AQd6/hDfG1GTnTEiZ12Vly9X
iL3c5467o0NDiTNRSEgbOaplGYfwnEy4RLoArqpzFL+svhfT3FLc5Sq1JRM0KqRRALMZEvNLPsx5
FK5QKdCheQp57StNPZzyx39VRVCYHMeWIrpGvMGZY9Jd2lTlEdDvEKoQkdlzK0Vb8I+dAf8pQF6t
lCWT1PUlM1AUTRd8VgRa8kd+YXcBoNz9MShQF3M9Y1MYhd/x2m9iBlHR/s+8cNWGJEgXXB0EABSg
73aB4AEn1J4EKw+DLRYn4994vnH4GO6pmJhBICUjbRyUD3N+DQW5tzcNubTEyRfxqAEwNqy9oiDe
FLHT6Ytt1i6toI3ZKgnESkqsulEwTN4t+oJP4AGkiMZWueuexo5wnPkGnlM7XEnvt3Zhi273vfEl
dDTyJoGSbqd1UWbvH9Russ43i+raHNZWfkVIRVBe3ClK0FAP8HIw/eAx2rFMWsLCQolW5jAjEJIo
m1iLwRUzua5ge37z9bxsCxMgWpd7ZXZt1itlQDXQ7X6s60wi1y+E6X8tydROaqttZEFq4V1Zy1hO
pd7HJaU8McHbpp4MwNx1NQegRiTclaBfKvLOQWE78Nhzi02c+ajMYvW0CWKOK2G26kXv1VMu+bW/
0m/rsyuwycJQERsOrMwXTwQLlZZvKV22UGrYC+Su9l9opwbPbTZu3SPQHoUN9ntccez9yyyC4KAt
3D62EINZUqsAMyhhI0OcMwbnWV86sueGk4beW1KNWBjxz3ecTBReGirt+uwtB+kCzmoku1uOakA/
iOdUfMW32y2LvXh+E4X+bN69KT2hOjAz00cXu5pgRjx/ThQHaz+P/OPZdU3WXvyCCHInGe6Fi/UR
vACrD3GOOLUcK80fD8ie+eQC4vabEJgpLUNBUg5qs12Gd2Ot0nEHdh/2pPYebmwh/4kNJHRv6ylc
Bk9C9BW42FrSBbgDLnpepj1ryE+/LDO8hsmLHqYMKZzOCRvSTSmB3bQiOFqBt7Ebtc6nWY7dbnes
0NAk6pbSG4v2a26+22SGGSkVR78x2ltz/b9xf/LGIRi/VpraZJ33s2C5YEbjXhIUxXDtBSBNkwOU
GR/6xPoTn/9YgsyerJWmxEaVWrkhRe9d1Mzoru1xTfiwPEbfjNkGdkQFK7XLACKyCXCKUbKN+UKb
RtKJonB2RCZN9+Sjbrp+9MHebUPpKlUGiDfO2iKf0FN1vn/q80xK1y42ZianAKZVRJs/3Ojv/Nlq
cHiczId6KPCWPDr6u/yJTgd09Mls+5S5hZptLns4S5NejpLcBvWoTA2AjEXlWjmfHUH4aX+xxsiA
KZ44nTXF3YbS9EL84Pcc1oBPFb1QKLJcxxrMOPUBA+xorSt3brRrdXHxP4HrHRv+JLR+/r/FnbmX
tJoUokcOxe6ikc51UZYsNQVvVL0+x31Z5SGzlzAqNYsF8H27Vq3ortjmVH32/9cYxLwK/wIlabF0
Zy21xy9bFoA9+j6Ja9ejK6/ISsldUTgmgt4mQ7BAg0BNA5gscWA3uUeC4rqYExxVqJDubJCwZHNj
8u/nEGA6UYv57MU2j4UDNDuCitwq3+QyBbF5QOzgoLkoc6HuspHKB/O/AzO+KfY8d5OWjJk6rTvn
D8/PUXt0btR0YUhOCYdne5d1qfJd2ggLmvXRy9o4bYNdk9cWd87y8HvAAYN1NAtK4f+N8GhtYOBS
sZFyDh3g6rawReGMrwN7owpRpKGInNNn2WDU78/LidLI4Z2tTaIfYUsvvzajckjwq3GVw0YSXwxv
gvV1gNzNKjTsxuwU3aFPLH6mj3AOmDli9JngYRYioJyUB6f9Wgp/NaGF4DM0IoTP4Np6MFw7rhjo
ZSWOJ30UtdhAd6pAizdIkScb3a3PVU67eZY7r2DDRqqd/4ti1MOjRus+V1J8RBVtmHq4w9l91SUT
3U3RsgJy/So/38Cedm5axb2rvQ4DuekyBh+AVYHt2okKPpbGPLEyK57fPPiUnFCE+Iy023ITMN87
L2ZVzQpE/eSCYlkWlZwmrL3ZkpTMaMIoKPdRji6Yxhubqbx5dk0skAsQ8krkbTBpeXsmO5aSmeK1
Zvj0Yk1MqfpltkF2ZX3QyoiM9n8F+UsKgtLnw2GqSpeJk/YG3lXuI6EaJbpKUV1uYF7t+b/EZyih
jWA0WSwr5LC2PfkmCFcDwy5E94WHXfh/pLVdV6XGojLarR+tXOWDJOzoBiCFrY0GUZ39CnUPGddR
2cIIiRnFDwdr2KfqKfk6NaHXcGXqT1rF3U/85wwT+WmhXy6oVnER6m+c6NcIZ2JcB0U0lu3BoxU+
jkmo6fiSt+O7NuMwkDg9Dm4vmLKl8BCOlI8gwulJn7VUWMlB7ssu0SmS4IjeFi/MOasEfaQLJZ1J
xcI9lGTw43soyYZkrtaAp6qWUcqzHqhh64sYwIbiQl0ITz9E2TSM3phPJ6xEVs0wbaF+lqbrKMJB
t2d7ynGLvIrOjWjP1KBzux27ZAlplbMCJsPpPhQtB9oDeEVfvn+9MvXLCTuuh0c7F7J/M17zvRYH
w/S5+VlcrYr1PZ7Oad3SzeffyAd6QvTMkd52r5dV/rdghy9bskQuAQAcoAiWYbzaTrf8SfOrkanI
+dpMWDcGF9Pb8e+M0KXCnsDHbPo2AfFqCT7zFJ3+QM+mJHwR6TpdY1EH8Bc9cJpR6Em9CCp9hsNv
OZM3gpFj47rKjxiYX0nyKv0hqh4Zf9ePtAP85KuK5tlQfZpqQOPHte9ZzoN9ZCOdz3W/K2s6XiSC
zoy1xo32jUilHMA8EEpWIvI5KQROrF3BvOnbpYD/lbV2q73IVw2FjlTPELenQv0togKFOyRVRKun
CrF8iyevHOTl++zIFLPO4uSj/q1TXMa6zyyYBg5Pj2rINBMmRbtQlXWFH8AqGsum5EzH2is+vLmm
NvefDL3BusyQhW+f7Qb1KoY56FFHDYAI6G7xrMyN2/wEFm7fD8i0iIvHlKmW7tOXLbPQVvHgFJdw
dkXnfmKvShPW64Q34sHfiK5GlTyVwrtpzNc/xhTxvAbNEQQhnQXeEugZfI2pve3WpR3XdkhTO1dt
Ef12gYgoePEfwbBcWfjP8b3Mn5AQJr15oKQ1AQDM3fEZU9imdRh/HHRqpYzhuJEddvK7BirYx2UN
xiDe38tLygJm9v9eJG5GAIw1qhTngNCT8d2IdeEhg6/j+WiSi01DjGObQrVCeoHiI5AL3nz9a/PD
f/ugJirWepSQlnGqe26XFhSVigk2fsxdUEgWN/BBP6I1vWkhPGRDR5CS6bVRWKtkJhDWbzgWvTHf
L98VcBBGG56sn1u9Ps/0/3oMTqf+vLNXUe0s6+TrS/cxU+PQAR+2sr4qntzuAMKJCogBYcIqfZ2R
Y4V16ZU9AJqxUFJAgKlFedNFe3PKkc2Tdy5GPZLWyvK0rH5qDjrq1izfeq5WLcUtMHqLtbrMTWyE
R0pSV94F9+FAhF90qMxkuAl3NRrnw2kOvZQX3kRHxSETrqoA0hc8O18EWmeDXfXoGRvm0enTxBFZ
SLzdWFrNRvVxuhFnp15JRrAropdjOcFnnyABUCx9+Io6E0X4oNWWwHiscL2ay6Phzh2j6cJg0vT9
b5zrvY0IHEqEt6XcRb7uBx/ukBk44jgF5krnSyLiH4L+PEyyw+0SWN0aFQXQuBWLZhy24Ma84Lvn
dz1K6G0fY+9sWTUmh4aTO+r1n/Krvc+apB+aFcKuanUfkFkFFKrUuZsK2fjBuLmlpUAjHUEl/YHx
LUlAg0W7F6QL/LxL103tfI/lA2n5Svb/56/Qp13b87mA58P4PxrahKBZsnJmlJVmzSQcUWboHEw6
55M815nYfwxULBVqtaZQsmXhcApt54LOqb7gdLNy+1/BXKgxhIVCUSxUlSAWpBdlaPyk8OchHMgf
WQ6Fu1BkmhI1dBQtAwe5eex7tRVuLgEVJ3lCfzq4BYL4KEWtJY0DALT0bh/mBrQ66FmZJvSxilJ1
WkGi3BBV05GzyYI9Ms6uuijpBecqTpICERP363y8f2KvCjdZa+52MP4oOBywB6wjEVjQNZx/8uUi
Lt3nTGPPyB1E0J/GShNIsQGsbJtIkgLBD8NSDUQPa42Ad61FedmjIvUPqa7G2KEW5bNVtRS17ZIH
zzRJz/dMytT06o925VXFe0qzLSKZj/Vr/qSRas9ySH+AemdLEblgIhuybywWMqFxZ20pjdKhZPV+
AZg96uF/wTyFaKmi9OMpLP6xOQ/2GTEg/DJ3ogMd0RSjU19LOoXgYc+LrnvLtKLRSZSUMbE0giC0
qmajTnuBTWOYShxLF9IhGw8uMIXMTcl3OY6RmhAJZwWCUaZQhxPHc4o77RRnoqels4EA01JEcjd4
vWo3+RD9sYgUY9TwVrV61rmAoBENULTEeXfPHleKpjGRp4AytTptEv2FwT/0GLHcaO2o6hmOISUi
W66ZT0tQA2Xu9wmFJ/j1LbX/zKeWSyns7dWqsKSlG1b4uOscKCd3YsJzeHiv6qWTiZXVRyt2ZpQ3
psc6OiCft+UQlcIJ8upshbbj1iI8wBCjXHMUQfzT0PIEvoRJuCcIJC80bBr0xLXhiQJebIHnRril
PDf0YnOXnIAbzl3ny+BscIb6FvsY0pMh3ECDWr7hdSRMqMLQ8lQgWzJbkntfPupsNPUDtf0oRz3N
Qg06Bjv1Uq4jovSVCHOwfipQrQgJX1Btyd9AH/emnC529crtEnwlaueFuN+xGxXxookX9efe8E5O
1aOofON0pzv4tJM/FGAuUZHR9//I7s+9t4oJG2o+YEvr3SGC9jBB6mP3DyvbeQ8vMzVOXdboh6mh
OjmYRP0zQJZTdbTJBH+M/IZP7QhbIBWh5ECa6AYRJCf2OanAhAnnxoaPBkUkawg35UsODUUuZgrf
Mw81mWRXx4PzIkCfxoBKZm4c0yGqVmVP9o9BsDWoBUJ92livkJ+ODqCtnP3NkfovfJQZaFVApLfm
moodudH5br0tsOsV4RZTvIv/wEA1CpMwgcmYCIEoRK4BIcIEhEnvZXTYBPaUsUh2xnlujiNQ4uiA
2jZJTaMj1M05KkwULcaR/6VCFmmWsvKhLJejWJgRif6b2mtat4iZ6q3SDIxP5eSuK0IA3kIK6XqX
1n0PvmNE+P8OLMB5TuQl3ZO+mRHMYYvqVKulkpLdWASAUDyglcS96n96L9adQY16X60r/CfhIgp+
pA7OkrsU2HPDYx5XqCJ8YX3oHK2m1Ep7Zm3Z/WcS6TrV15zd4hpShdTdjpYCRIviWYBpU2ZOFiVu
+/PNmu/q2xe/PDRiOoW3cJFC5n2eSWf/gh5rsHZRZ0qI41IUwyPtq57HrMhPikCqmyOgIBGaC5y2
KwUlTc2cAvady+pWIKk54tkzHpIjeS5Eyv9WQRGEXY1RCgj/HMUpl+4m+3tN2EJ3aYl0d5O3YsqY
Mbg7j1eUeBbpKRhRxgiVkD4947+txVb0PeyzYZIYxO3bsSJRls++G3DCRu6mVvIYVcxbsCQjV1dI
TADdYkH9t+UyJzvn3TR1BqqjeK5j/rCi3Tt7+lKm/ZRZZ3041fAbt5zu2ZrS3BdyBOMWUE/4E/mC
mhZwEutDpEoKocYean16HLzvSxmBif3yiVuqHt4RGjNF+vjChYp+Tam/FnNKNNo/2Zu6iE2GR5Gw
Y9osSw74Uo75sTxRacsPAfudLBF9+WZDtPf217pBiafrmOiQ42h2YOOYO/o0dSxeX0VWBvEYz6XS
ui32mhHyM5zpFJQS+lMT5NnXw17mCAzWAGY/Ugmv1to8zz7cnoCUm3kfcJHExGaug3e65N46J0Y6
zzbaRy0G6Z3XqGSGBK7Bi0FLe55MxLrdoGBEpBw+zqLfzypx0HwVLzDaPDptGcH408be+jz0aR6y
8SweFBfB+wpssKBwM/CJOaGEmdB3W38YO+DhlPoDVLB8szi+aeuw5al1IX4dLVVVCY2/m+S27V0H
mlHyOLr9wl/+cMRIEc8WDRX4l2gEcVs5THIoMmhtz6SfpwRLj2s7o72AIygjLBLDVWnljwZCNOax
ncr9rof3aRYzcQjl69Wg0SzvJ+NmfpVEWQa28giBoR7jy46i+9PB1J6mc1mWUj3/e/r/ODUf2Rh/
I7K0ak2ahJKlFZvo4hTV66aekP3WUYpfHVD92KRGfYNCQJZ5s237adVxM4R9Ym3bCTpt+s0XydZ4
kHLHo5RPJ+AEpX4DsYVY5YMU5tV/0VJJEWZAO59D5AsF6bR6CjcMQ1UwTbrVR2jfr+sXQvHsJFoe
Ns4k7o17S0xr+PBTaCHRa0qQsErmF9yetijPnmPbi/xhCkaV7cP26bSY43UVIFiMpGCWXGtRW2bC
mCjx3AeZZ4lXDy9E83LpBix7mCcs53hsB5acJbmip+dm217X+I/RwhIGJKH9K9yUCPNnOuqHWoKL
vRhu1oisZwdojgKQUwaygNqC4Uas8oLqllRrIGRxU0b67KulU98GiMn69ShU6Y4TLskKEtnM6obI
/Lvq237+sVfah6l9iQTuyced49064ZLBqVe+5KI5h8lFmfr1rJiNWQZ037WIC5jKChp1PamDNnIg
iO0SRSfsf1mwjxYH4WoJe42ogKjGCH51LfZKCyH8JkM3mNSZV5JHKJ+C/FN8TS+dQZiPqAbrIMe+
5VSukFzAQhaAO2cvy15tA2p6Oe/eJzpOufBxp/P3xSApK1yLfLbFLIEWqIX6BFgRFtC/K7GZ6jJM
gnAQ33tooYXfJxlh1bad+zj1oYAllAQVczqA2GPJgRSF8Rht5rT1P+5dqXhcX7YMsuy4akmLAQHd
LvMwoW3NfpudHVsnQWr64C4dBeaNsQVVwA0Duc2crv3RrWZ3Cv9wMp1V9ChisK+83FVbrjWdjWxm
KulDCEvgr1I6Pohm3yLVkCQEO56rbsZZWbVqLVbyxZW74EqD5YC68LaioLNLzFAS9LmeZiS9jWfa
e/dW50pVZrvoAFQCwofwS/BVablPHXZWqFiUIPdqh+qEo3grY8CQmZHUUZ9kv3uXnrH/OeNBT4nc
zyROTCTrjQEMUOLHAV1egAHowQzkNZ1rYDLNh+Qq4Xo95jVXyduAhKXg+CXaUFK24G6rLktj07uM
2mHQIp06SIGh9cEBcj/XuHvkrq2ZFgj9s1z5L+IZ1pKA9xg7ssIpmfD/jX3pfKSXrHRZ7mTbefbk
mW3711HXYH8FwoqJ3QXKqKWZVr99MY3FlM3AGbewO6/F9bYckUhAoiEK55rXQ8gOfw50SeCNkDg6
0dS/IokA8oNz3V8pdfSzjwqzhjCGd2Wx1l9tF0j2bnI8YHgs/fMQVOOs3vQEVFBpN0gPewyIt2Ck
O+EIl9NmO1rUjA3XOcRWLf4sXipoaDDBetGUMqEVfYEKfiEIWYv04l7fGaXYFbs3TTiVj3VoD0LA
XiqL6QQj6WCAMERt+pxfCVy7dMUDm2kMnHdiTDRaD7G/hvQwTZryhIRdIw/kTO0HzyrXEOMbob5b
choqccoJ9ezPruEbArq02m3nFfAA7Tus7acHIgopQ7OqKtpa5+/insPxXx1RAxnr/w6lazpl3POW
N5Q7x5KlaAgTcCd8fqWo6n9mJIN6Fa/WPkuX0n/5Ir0iBB1EOUgoyNDfETDeAMwl6d3DwuYZ47Gl
6HVp0/+aXtd0Cq3FK1EwNYqtFdSZOcfERrxdft6FbJwC+QPl0Oy0TvHm3iK56KN8+Miadl+Kpx0s
ctBvsoTXn31nsd4qPrCgyPsI6Ok2dJPR9PqHzaDEoNdc0Pkz69D35uHr1151DpblOhbJqo0e3Ml5
epHa3RBe+NiNl1mlekLUZqx8XS43D6PjqM1TvJovL74Hki3NR+Um+LuN45g2uAbgKvnX+2gcm5VW
WHori2L1OjJHxTZdqViL7WhkZJNQzLdflBMTT6rwT5ACaNRDuyRhpSIE/iobWQ/qd4o/DDwTr36K
AkBzmJp7CrTy5MI15rwM0EUBg4/yrfC4dirkvO4xXfHB+6MtDXamr6mZu7fgIbIJs5G9NEzcyAon
BJiIr+TzT2AmDo4cCEkUAW+0ZgkEuKf4SuYCoj4e4jJXVguEHJMpmvjXGas9NLaOT06q8BN/Ymid
gV8t09Aa3sXqAppu+IgBOByVEdi4O2wYZPpp2zpMPkEfzn5Bl+duyqmgbVUc6yrqx9ffy090bNP4
grt+zFcmqNsFj97cmGvAnAii2lVuiRMPpcx6Do2x7PfDU/TC8KIG0e5jkrPgFaYNxS5aavm3NDnN
VaVauM4bYNm1CZtJmfLku04gXjf1nJQ0JmLqClgWw8F17bebIel0tEFvIT5POxd77PKQnKjCShNp
Un1cTKdt+4HjtF7fb64CYfpJ/OJ2kaBZgrXGIXYEqVf0QRfOpFRAMYx0INQzVanBf5aEllW5xrVw
cAWDY2OJsr4WAXJYUHf5yAzpUU7oySidmOvFv2k/Dswwk4CRaU5cySbGrMnB++QUIY2/rltov19+
4F9t2wFPGHpzb1bdt5qotgO5IaQSYUNAj66PfLs001yDYVghy3MpWridW3bctT8d62DKZtPJVO1N
iX5d0GJJcQaM/KtGJx799NvQFgQDVPFHYIkivs56rJHcNSSypMk/yw/Cy9K4Zn7nywKepR/k0qCJ
gvPBDfqDStLrJJfEFH+a/sgucO2iNRbh9zL4prq6rEyt9zo3aNOlOf+1PGRtfoWeNk0UoRYqVrue
sIkeKaL/XSdy8uJl5/RrZmF7pVhx/mAi49N/oVG7++DAEzOCCd0+hG0ecrBVkJ3W1DE4pQGxu7Mv
GwarR8NwknvIB9k/dlmrMgNATuck37o8QMHeK4eaejoANNDVhKYsLEf0JqCiJQcO7b24+d7SHYT2
Wfk7rqUm81Ve20ZK63DjsKhnAalmHLRHDGez+TNPwI3IN7snrtsaEzXfqbERhRUnTcIln+GHgmaS
Z6Rm10fPDM49PrQxqPOuf5wE5k/Ptj7D3DidWke3aKcUp5Yk8y+D83zeOqf0iqqmUckSl4bEfCAM
nPTG4Gr23qYCeObbDrySZKpS0ol3i0eBjj4S8zsV3sC9ET9yb2BAk0mEZaZA4Ufdh9Uto2AYrtMT
QuWjcAEE0UVTB2HnvGIET8BC9s3fjfnh2wRUB0gAE8wayg+ptpbn3jYjGDLw4NaqdrJqZdZI9kPR
MCW9d+yg7y48/P8TxXkZ/64sd0aUXwun5HNTHpFQ4h5ymIeqUlcXVIVw8qL2LnjF+Dv24Mnm7dCs
3FcVBGiN/5BC7h1FWKc62d2n3k0w/6dy5hzE+3h/NQz4/NZ+hkhQwb4A/gBZJxRNBaQszZ/Ldz8X
ZrP2LgnScr06fH6vG8iV8w/yxZue1dfua4d5wjVroJ0zPCQu3vE9q8hfQ9GiWstgAPriwTuyn5Kh
8kX8bFwGqv9vptgkcZ8TjsI7u1deM3oifcGtDRGKkEEnIwrb/BEA+vE9a4X3yM2vnJs2kb54yKP0
T118Y+X0pMY6JDDDdlFh8JPzTfRgY3Rwiu0ZY4mQu0VbHX6Z/u+LGWv9C9SpdnAz59fgT33F5gTd
Phs4aKPQTbxAhLtSoKuQWpPPuw1PeFzY7zy0Nw3tyO2mNBGiP1tUIihGw9fDutPrZ+zpVkQ8L8Rn
x49q67KFtKBwheksoImtyK9PJ6BlcD3JTklJekXVclOLid4vjW7ghX4OR328ykcoN7VPn8D2jlHC
GPt6FGWBeFZg5l7KE19MeeLeeNzLM1G2YHwRDlJMsx4qWjTQa2iK3f7p4ADXoZlbVWkGPAJiLufq
m1HwHHzUWbdD2FCo0wmn4vvfnj0CgmVhebPidqZv+XppYAw3RP9KMUCTJ2eUVd0WiYvgSM+p5Mz+
tTJJMrXvIFyQ+/8dtfJ2ivKr05BXf/Se26lllNa4xX3Diy1BwT8g1MUmpQZXZnS3g2yW6dlJmP1h
5M9GB90Qsta+A1cdDo18OlUQ0GMgpGhs3uLNSEQBdiaoMHL/Ydc6yBImspfRkZuOM/lxXHySe40o
xf32z/OvfOap5Lm5yVFlokLaxPEmGS6HPkrTmy7suN4neDHFImLReoIThY5u51R33pvNrC2FBlTO
/gBa7hqFlUxOyfGZU+UFld2K9E1Bdht/WQRFN3AIENTQrrcUJLXsOZMz/PniqH3DXs05mDCIPJFT
at1PMiZcg26KGXbQHsW6LqIPLpbk7QKMUUZoDk7jBaLGebjv44TvYph+G0x8RP+f0cB1St1iMFLt
jtdc9wYAzmA7PCym4JiDTK9o1EAjZxj38t+UI7mquJy0OimeYP649K9spS/wC9bwrk6Cx/zn1O3U
w7geb0Ff3mk44gm2s8Gh7OuRhLdNvW7qUL82BaS7y4s5xJ7D3ejLTH/PjwSVN3wlrXsj7pUSsPE/
fhbzokY55i/FRJHKA7RJPDU8+oACq/2HYwdxh3A/odcrS999dy0Hhy9AgQfTLc52LvYXoKgDsa6D
5VxO7L6agWEC17ZGtARt3ORSVzDn6i5eLNidPI6OcszSsFVagu7WEVsTSFeNgtVVDvQQfRLkOKnp
N4+AqGOJXx+vi0QLGLefSIDoolKtk6vkA5iUttI487rizfXegNvBW66+2/vfZgQ0VXczkmCcxZNT
nsi5ouESyIc9Ig6s3bRoiN9b+vOwcmAM+lZAZn6atWG1ftFA35BkkKblWIoch0xsLPCZ4UycNr2Z
VTJ9PpPXk02VGKtHdoq1BeXOOlwlG8RFgeDDc4GzTotOCcWL6qlgnvRkF+Ecx5ZpoRJ0RRST5XsV
UGBqQ0PJUE8ZIEOii6EbAOMpgntcDvAPenmc03vS17rjWf5MgnCAqsdp2M3qMqfKKcDZ2qZV3XUC
LuELzcCi2dKetKxrTliSka0zZO+jaP9VYSzC8ay7NLxdjWdvmrSnztw2xnEs3yxEu54TPJYQxRtJ
H2itMmVgTWGAio/hNZp3NPYD89fJO9AxPQH7wS4rdHxyc5Ex8eNkgWlk6Pwp+ttHybhjVqibL9qE
s9uawFLmupezgQIxJN9wpZcTlkqXZycsPsnTUJrTUpHSXBZZhCWAAIuMGphWUJNZI8HAA1UsVSPZ
Vo8AI9poGuQ2ob8ZIRpZ7/vDevsZGHjEzUp4BlfcGeVCeLKWnn8KkgOgC+sC+xuM9XFyB3s8+E1A
gFpjMMfogEjjFJFMqohkXlMETbJkjp1j5OB6r2QTCmgYamrVGhnaZXixNRwnW4E0eR0XCNjC0Lt6
Z0PkfFbZL6CVsrjFuIB67kcOq4Wm9z3ZVWKrj3v7l7phCtVoRRdJDcVc4Pfv5YKQDOr3ovQSCnHc
xoyiNJUc9ccLd6bBhyaw0YXdshLiZvHeup3tRQgvo+9GEGTloc12wbGVXku4IfxVGqK3p7l7paUH
A2PvaUuDgtZz795vCJnm7SXACIHcY4JJLha4c21AxkQmTZyymrffkokXQfBZmIS7/HyUDUNSCjZu
lAhq1pUkCKuDnIgYk6iU1Wv6lKo4X58cs3HRFO9/LNKrKLUOvm/3TtqzzsBVdXSj9cpWLR0vhXO6
WxgPMrJ9ULAzIsSE8yE+0x8rPUYPPz8Is/x9KglSMcsAuPLG4o+o8ZJUEvQJJrmSR7DGAO1YkOZ8
M/sKe1k4zfibrvOcrdmQfQMvDXasPgUUkOQqPmhskdqWAUQu13riq1MKxJYslLQEePSaxOya6X6L
jwJcxrE0qjyxVC7YulgT8ePFfXYcMTETTMsIzMbSBtOiplAyDDpTh/g+8ZZ1oLSFnMhWipOD6Noj
tBecc5c16TZ6mAS08s7wuMcMwnF9oVsDHeSeY9GtQkwubl594RaOy53a3XcfPDmKDrwC/xP6/fpc
A1d27Co6hpEDoFwPc1O/kKzXMktFxqGh26AKEZOI3GzfkQEKdw5LQjHiRnOEZK5eipqsrAkw1VJT
iDeTpr4yD9n49+NTTXsYYYaGhL7I3Kz9tIYjcbhU0KynOfDZUBLak5yMNU6jHGJ350Y+gVpHvWaH
BR5EztWk+SzNFt1AL1VnZw+moL9iFfrOl3o9u2TYD8J6c+GFamVDxRPqIuzIhAso+rnnpafs9shT
72ng6jrTSOP7HQwOw/BwQTYIifIudnKee4xh0dhyKg8541F0U6jYXVGBWrIgodNaKLN2ZeMTLFMc
S1qThK1ogdsVMmO2BRk+4vZhlLeOfrqfdIA+ZIM2cbou8DWdb4v8w41UVfedHVEiMtA8ny1CYRNc
lSqFnc1aEE+XR/wH0ySaDR+KcYW7FBHCmyanQbKdwawPkznS/ROBNzRM65WyZGSpBQa+03z5nmFr
KiIVTGAa0LitbT8ChLLlbxU8O6SiMH43EpBBEJtivN1UcO2R3xcLwF9DJAjbpHliAQfLw1ExCeGT
xAi7GvmTRmk45YbC03jAFk0xlJYOKSenaqoFUgHUIpZe+cSqbGcjQAJQ07jYPCSlQmD55TaXLZkD
hUqVUyL5rma7ylX7x2jZ9Js9NjhSZorMg23x+TcLUmmPwGEennmtqNBK2pzfJE2OkfLSatbrTtN9
p/fZ+vEREY/uZhlSfY23juLW0pKvKaZoekzSdv2YXbn3VCNAxoLJaKWkQPeMG6sQFWr+IIfPwJr4
cCR+1LQfR0fEksj7f1SNIHXEom01nmJ2ZeXOC8xwSNlldBdRlecErImH1P5nqLqDbcaqKJkQfqdV
hrdQapRYl5n1qif6mn3wH+mMfyZeEmQ5B0xN9smZNj1x2VO8VM/qcicTsTNnK3AQqSawQ4jygkwb
7OhlGC4ABkRCp7JAiLP/2QNe+B791BpKfIXLYGDffaz1FoR92FxcVtK54S+BUACjUflPoeM4UBOB
U6AjMYelno2kmAhmb2H76RyiGXhksFu7ea2TUwmdomLmMRQa1rvLwjf5diWtxLAlw4KxTM7v+DKq
HJHwVZ8H7nFv4bfWS8zJDlLmVR8FvJwDWHhF0mLZBeECNL0R4ktjoO/Y9xlP5WthUXstqF1vN4+w
JGw9rIx6D0epSHCkMtE7XNDM/6jPjwx8Jsy3t6kjgoHJ+VNKawGfQkilGHr4pc0x3b2K8zvMtRIT
DACnqO6HacFR5o5VPfkSzUbQM7Ed7KKfQ7OJJElli/IiKc9YCucI3bslQEAyC5sdwAiJUpxqBGc8
x8F5s9LFe7iV3f4j8OaePegcCJCQLuYn1rpL5BxoBRv8FQ4aHkg+dSK3zQXflHxh+HSsVatye7rj
/WqF7JHD/k60x4BYqKf9EsM3kD2nlDS8deXfz7isEYmfiEGjXgmbLeMcTEG168JsmKd4Q4T8mpy0
QEB3K1PqGJz3dPyPWI8BYJPG9GXpgX5LjTHxh11Gm7DTxji8DNIWXVJYZm4j6mA2zpKg9/A68ENQ
MBijzsAscvlqgE50JQwrWq3VvO18NVjrmyRqC/HUJLOmtAGa+SqXarRsq1983lyjB7/lUa8sHsBS
YPJGRbtW7KVOuiHFhy+8SgnK2wDmptBivG3gdzgbPR8/ZGciE9osFoYTDK3kXJZLY/2k/qbcP2xr
/7vfgY7hckk2ItevtsjCDlk0IdPqLTeNLeKR4oVlA0DOWIvACENtBicAXPlL/ZMI1OBWAmLlBGLr
aFz5UcKsWFuVIez5ce7wMJZMhcAqm8f9hJ4na8imrdixPI3wx5OfRkF83tS7eWokLYJA3mtjwxXx
+0PxvQmS4gft0/DIUQbCETqXxoe28FoeFw16L67d+4x4vdCTlt5WVhjP221cH/J/HB3lrgsOVvYP
f0Z9wfAxoci3OefhIxR2Fq5GbphBLh/4fyVF3KDQiu9i5Xra4FbzELR22Ai19vkpF6qqOKv7PN0Z
ktrIzpYsY+AIXX19Yz/zpXm9JztgtxSjv+iFUGxrb359NEhwNBvIRf08rCRjt2ZelocyaAHWzerW
r7uYoNOTAhfqLQmMZEFvXwqOUPtFy12cez/za49h2OEI2FMaBmJmZHoRBGZJkb5ks3JTPE6huUWq
SdX6HvWq1RT0ubgrIoNYPWxDlZ8OFBWHbmJzhB7WEOYVS95TqMiqwlUb3EOpe8r0X165mDIrDFoK
MZpJhEKzi8Fn5LIbBEuNXGWy5IHsUDW7dAZ7IgbxMOEQyyI5mOIt/uZ+aqyt5AyEpTXECXyuofTm
pNr3NlttwoWpr7ygOlFf7vPU4gDYOoLcnFQv3wAR26+QcYRVgmqMmsT7+vMG/05Sri1UVLYPrYA6
6Tp9xSB5mIkzqHVOPl4kNB4TacIEQvN8T9+6AaJ22QuPvnAc+PjCs3CfmO6+U72v9/2J7i+VnxfL
JPtOJ8zgCvEPqkl2i5IT4rUNam9c978czvOyH/Io90KtaIbrkxLEn2sI0p4BhlSr4eGNA7J/3pk3
4eNQPQ2pi6DcwMO+ARI8vA3sMmtCUWpoyc1gn+z19Uc91WokZFS5/ftcF9lXqZjKoHKtVdsactIj
IZoP8nErB/SqqE3g+TphT++Pd+SXBe5Gz1FJerufIeS+4AuSwzfbIN3sVfHMXy9sRbC8CgAVN6kE
7kC/BhBN1rcYbrzBh3gkrBuhv9EhP9+jrGLEbdSnDmRRbWijplAdX0hXDGp3c7QLLTMVZEORJHFx
scv8lpd/nKYl79WtnMnZO6KQZ7rfKqM1NTVy6cX60sD3L3ILzKY68pdsO5cd2EQ/PJS76pT/W7Te
FCx5Z4qWAtXQktfyu+c4EsZvIyeVe5oRW6qRltQeVHp5JHhY2TEy669qKGegW+ZSYXQpY6onJJjM
W1kA27xTVDh54fAP25pEdyAcZjr39vmuXZRMYfayZ3228rzZpuSyvTVb72GkoMJvm6c+n3zImQyH
b35cNkPzVIqyLWN+YwdkGp7+oCCgAXSqBBFm2ZOjAx8P3/MKWHfDPJ1lMdveKeDGguUG3wasSIwO
pYzvE58s8Akyfy+6koLi7Y3yic6eZFwi5Joo3NGkH+lgGVjV6XdZPywON81ZANSB7LBbq7g2cX5j
uBCJatm0oIan42YIE/J2N3ZImEsoWeXYqWJfI0cr4Uvk9k/tlgWmSCDZHvsMuxii0lnLXRgezNxs
pDqvhxs/xq2CIA9PbzZAWy4HfLxWcTcVtHfI8YeCPDkJce9n5TLqHqm/YcGPZ1rwO52RfGtnn+fx
oPDJzcxQIHT2GsL705+hgxZDkUiVrwkhYr4ihGCIS9LUUA8Np+/Q/jpclnweQ0p2L3F2NBHot94E
0r/7EmSCNTehKt6j44UdnK0zOBTnA4pMK1h/5N/NzV6gnup4NaZ70VbZ8Cib25k88YKBmqM0sdWd
9ZSvdF31J8A2qXzph1kxteAI0sRPKMDjybeUzl8YRYk4NHTJkgFmSN11brNYrbKDAdLgGvietMG2
VoUyuMFPm6F65TmEyLA2sGMyycxoiWkLoYJkVGM3Ss6bJE0MmZrz40UCesSq0qgdxdaOQyVcYrcg
kWoqWQhV4Yub3TMY1+uSHxhFVbzj2ppZeyGrTWoeChIyIZRlH2V8JhGf7ZdbnkMUyx1ETX/SaoTZ
za1JlyrEblyzoV65RrMmoQdFI1gDIlapq3DRPjOZomWnsF+JcjG4gSXzZL0VCPh30463rHrWDXPB
rF0qEj9DM6DQ3ZXXj0GXzBiSOlRqRfntNhrGUfTIscDji3SMAHoWs+/YiVGElajx9vSdBXvFTX36
SFDku8LIYnisl/4uv+VOpF9NxmGiPZAbPA6MQVtiptvWwOXeplZN45VN2OWYkKiY5JHlnw/0sR0i
zMA4kiUdL9DUSOv17DiRV1wBzOcy/dIjM4ZGQsfknm4YT+VP0W3z8Jwt1n3LoUmboKWqJIv7MLmB
2JAcJcm6mVkn7AVRNs/kzgmkMWSt4DJrd4/lBdsa1geh9JigwWRRjH7YTtsoliz9wdNBVapX3qPl
3tIrCUoAtl3O0t17izMfHHBe8QBBkuSHrAZyjYiXWmdya+WVSSvcfnrohs9EmtnSZKKJvHKbbh5m
9G9eXpvNFk5ip+AC1/6qJYCv4SZE4uW5If4Pv+B3UNex6g09ivAc+eiR8i+apdHyicRBFOCod9jP
qgbH+lNLZIyzdClWjusPCZU5ZdIB20zVE/0tCKCTxxjE7KfTSK4vXOXbUM8rQjNLhM0jyrLMJaIg
sNuwaNG+SpKbZ/gS4uuBjwCTl+ktIxQp7Xyvr0YXJF9Ay5a5jpqpia8vFsXm5wgoI12U5jh+lVR/
LHm5+In26BfYB0Xrc9b2wNy7smkpcA4jt6st2FatIjlXPEqflOtk/8v01lWDKHKDOrTwkzpnAWWH
M1mHzay/U5sVO431j68A3QX6drh96SP+uQa6N5QoRVeMd4MITNwojn/zewVfTLOmBZ/BAI0WQwad
UEskAnIO/nDJK4IpcixF5Vv2wpzOfROlwU0LGuLqHIB0M5WLuVEOHSCP2slLLOaItVxtYfxx95Bf
EhCymMRAQwvCrSnSjTMzvZgdy7g5QxppCQth1i7MDJ/rA40u/5Kiuo0ZGv5tq0VH1yi4ZK5384TW
oESgYjccaFcV2t7IX0GpN+IGOgq/jfUDQEST/g8a2ZWmHxLS7Dzq8+x0k80lTWvOwlv/DTkjQo19
5yiaRSs+T4Ot85vhGRVMi/UE+e2uDqpFkUmwssfxhBFIHzFinNJgzkY/KPgev4k8YpvXHAxWhHgT
2Mo8G7kCp0cmp6rTmb0+ZvAUXmesFeMXPJPV6CVAQvO/l2AFGxp4f5jaaQlQisVPeMrvLvvqHWth
dv8lxxYGE+e5emOWu9eS8UTnusGOhneLCYDnIYVhm5ga0Lum6KYUovK8ksMIRbDCedziPa94a0ts
f+vlQhJQMtRmTgIcOyMPvc5nsw99lkZJgCe49CPluEuiiWSmh93tRDS3ZdlvAB/pLqvcoLNRGqqY
m+GNWVLnMZk/9XCxoFzAulF3kyuDmo35LGnQoW7SXENzmPdzA4LI3BQitwCAr2wXj9WnoQdVIxJW
QBIfntnuqqEhhMlNtmKDLJ7QfJ/UQFLyVIah1FEO9i+fcUvu1st22Yxo2Krjh2kLy5w0FnYCG5xc
ToTghXWtV5GjRNi6hEpvVl/9+iOcGkaNL9PlWq+6ZAVjBchZIXP99y1XPSLIA6KxXjuBd2mg1mUV
2H0z1ujp86YlwWeT2/DRQhwvwg78RFN3mjU84L4Nv9sfh9uplxArUkO2m3F+HnI3aS/3SstSd/Eq
Y6lmW3l3t6Zpz4grOKtw8zwFVGikFb1DziieBFrhPTKkdJ7K+7fDvkSQKmWtgcgG4l4PgvgMM77s
4tWKgmnrUo4Ej2Rd/SZbIuZZLUcM6yL76o5SRscJsucs4fdtAlkXVg7L1rwnLxCY0/zM2PbsYtLi
HQ4atZ+yjZuMUI3AVugt4qN/6EP1ph1ef1XelnT2pCLqWAb6muPA5gpPnsDXkmMRm0Ts3ZbVXat6
VXW+cRQTxNECYwv/+6ywdJHp+kyZEV8KYC5dRtxjj4ESbBrpVpnbxRNrjF9mdAojbEkNqCo4HJy/
Wueg5jSjMP51EGF81wfFj3uNS8bdsNnx7qGVnIllJ8z9M5sw7UJJpmHtmwns0Ytt5R7Pag39IWyl
YtLj7hUuGmxqOTS4OMxwDNXaUHw+w/yM5T/MDJorsrqQUBcR++8AkMQqpe0HOJ7Y5cq3O7ui9dZT
X+CW+Y+IWMm0v4tDo8IjOq23y0KbM/tndU8oRIhG0HKeuAP01A90N3B8F46DO9fBTZD2F9hrbNQr
9za5vIARjKdbpt3A0MVQ1FN96Mmq3gI53tCXoHlriN56yfNnF+jSNQCHUHHgbkgZ5/TINf9RPIFZ
deO3JA8Ppglhofqd5XGqljyQfsyiA/p5dPPxczBsmyfDGD8vVRxUeLtjY+rY2HmoX7ee+o57kKgA
cjeP5iAXY2oCeTUt3eXbdoDO+fhcp9Teu+avxwUor5kvfmSRe3+MMKsA/rQwyDxDiT6052i8WiL9
F4vSdCbxNf6Mml6K9XaODlc3W33tRbhghyNl0JOWZ2P+N/d/99a+EXxHAM8qhdcj8P0EXG8q75yU
7rR+fJ9G9pHeWCX/x85pQgZeYtzYQNTGqsRAOiD5qVxFxN4Cf5il930AB8v2TpVmOQuHQBho+1/d
qqCuyOj/x0YmIfgmoh1U2s9jpFY6WTMwz4pl+TR0F/X6BggD3RFDxZaSIBacHymBCC0cfPCvlSS2
B1UEvmvVl+1PpBQnV5hRmSFt1s2Ebsnh64p7es3+OnsQDSxK2DlqqYTJQC78P50cZ+HEH91WBzKM
DyiLhi2UUXHnf+QLe4qN2iTmKLfdGGVbQtfbbfwLsQkIP8ObGLi2hvRdt/thzswdPdV+x03bz1DS
wfreBbFhCdsUCt6BWo14Oyhtbmawcip8rpfLBLHDgDF9CqmbrvhC37ol4xsWdU6/YuhqXRTfHeJ1
iCYRK50W8jPfwqgCohW7t93iQY1za+cCfgquFYZm73vBG/0ZZs6Qr0/8A5mhLyUWBtylf9LjGYwn
Y4MLES3gb8ocFPCdiyh1EA6khPdLjAz0PkTj+4c+/Wfi34dqaRRJUIBtZ6LBrm4KfX1RSLfl93rg
OiWWXRe+pesNUE4296wFjiYqQxOzEDWxb3pmv/WbO72eROs71h34X3mQV+LPH15HswpJIOXjLFBw
JbxCzlhrCdEOyNXM6LczLR7Ifm4y8YY3BslNc2R0fuo28wTrb2ECBz4UZw/A6ACM6n0LQ+LP2m0Q
jGNH8N2q6Xn7qGzLxV0AiuhjTCFA6AjKidHuccLfr3/9jmXhcx1vezbXrIgiiotduVC7ffSuPg81
lN6Vrlyq9HGdJLJTm5ywc2Flxdvoyzufls8DeXBeemC6i7GBPV3LKNuXHPc6eCWq8uZFFo6GK2LS
Ka8CF3n/dMUL5Wij33FLw8eBov9XqIzLuOWXL2TiFQhhWmLy59tdpHH2/xgqnfChQ9s4ktNDIaOl
tUMBVALvMjftbgXkbLGTr8dRKOE8iGkbid3QwzNbt6STryjnL0QE6uqIyqC+C2cZNXTFobdU/Ca+
JGmjeZ90CYRpNeMn4Q1UdaxdV18VWbyWUtjRCDMYSkqFr04ZL9BrGggNX20kokYAnCeB8/amGhQ1
E3YYI1bubP+Pcl/MKucusLvH3nOcNQzxaz7ZAyePkW6ShVkBNWtS5BfGlK5eUnUIPdl/emKnkFmf
LawUusmV1jM3djjzvpGzkc0RTXGG/BwhQrAez2qpSE43uWoabGYGe9B5UVsnBi6mpG0LBrBg7b3O
cNrgDs2bdEttoUuLUqN5CeYE3lXU6GKecMEq/WKdZpNlbn0NcwCOhLwnarUXNkVFVQ1q/j19UQqg
abiDyQ1GIjbytsFLJS10lNHMoM1kjgkk5ET4w6ShrvNSsqysbjLd7d/VjtKuA/2SIdzotzeqi7KJ
9sCzes3ysBUO3dGtHv/xzLqy7NDWrHYYOYPWiqLMyHTjVq4dkT6sTKR74h+VXxuc+UwSSVycWzJm
WWiNq3Dq6K3KTmkiLcyyUaz3KlrGrjVM5Z42sgf1ZXj+jb9BTpLbr8bLZp/7Z/AHYkxPzgyYR1iu
nbixQJUSDiLQ94NeQFTSk59lcm8z3a+lVnhrS6XILhDrn1gcYjtiSmCB2ujIcmOIfufvd57J+SSG
B8LWLycmPVAQPTWnXusE7yeK5wIL6ILZBoXfQORw0cBBBcvxIKY3uBwyOGLb1PkMWHSMgWKIY9/y
cSYM4wazE0d6q0B6hWIN9S5e65koQpQGXLQPyYONdGyPZBQDlKP/g9ZUd53iMnbNT/BkNkqGHBac
ZU8Q2gKrnQWf+2YF0riDZQNI09P4ublq6J6oqjwdyM1BS2cDXTOikPGvO9WQy2rvBsb9Il3oUiFU
l8OLdKXx12sqOXUaN2foF6U5UGyN6gWkPbsyLh1C73+TegZVzDd7C1xsIYWxTExP+yaUCTI/TXKZ
sSRbEHMcMDuZU3aPfZLi4ARujsroBals1prhJ+FgDmMaEGdOLY8AJPPyLjWC0UHZb4oLYc5Wz7Zk
Z2O1yOaoyiCXekMuvbibIIHMigbSf0SwYdyQnpy8iYXYwfH0tpwBy4YVypiMDXnPUBS1+oWNtknM
btflIKQOptfge5yVFvu4RUW9uY40IvW/xcjVhltJco7RtT+mWE9vRWeTKJZwXsOA2Ry6QLoQHZ4n
Dp8Ug7oc2N+U0uLbwDD2U96ubXrCwtJmoxnsmjG6A7cawDpi41csH3RkVzxybPe5H6EDlIA2lqR/
RrO0yxYR/vTWeTb576QsI6WlGsGle9aQW8aLtPhx+Vp/2GJPNj7m8I2VihYJXmFNwi3HlWM3n6Qp
i7YJrYJB0XxHwcg8WE05JKualsBONYwLotJxyacmDO9rTieH1dUYRvG/jPb02uIf+v2RTpQJXbyf
meFCMuFvdqkbhXVd2eQLo6Zmt35inQsQJAORPgtkXrzvuouBY6Db5ATVhkxBFj7IOijZyDdyPeKL
R/kHkUUa5p1oHcI4+2qU61OO15IQgHT5KuyaA135JBhyDFjtv2bkmvL1qBU7nkyIvgFE3i/luH+i
nKsc4L7IAyjwUgijAFKF+je/VPc7i+Kz4zzOatGPaoAs6vohc0YOghCDug+rviP1URTjCIRqPscR
P07pcf/MIqY7Vhre6l3QlkOwsLguGu3gkw+OJexSmc7bGYKVHUsI7zE3KMtGav/biJ6Nov+9Iv3Z
94SFgygPewMJHT/sQdqFuz62jyR7hzz96yntKxjpfE+pzAzraOO6Jsbs+tP4xSAGoRJw3dPYMhuV
QIOd592A0amuWjPfAzKuQdWO4m/VtAvA7G584lg8q6NCgblfSEUp9cuXCnHHd+vp/TfcsMro/xQD
sJdVDabGsTMSBb/jq6ISPGoUrrggNgLiQ0grJPyUCBHy9eNtaVmVElrMBZkEJXOYe3WGpQwXTLyd
oL1i+6aOKtPpZQnQzwt4ennkMLVQv9LkTnkgu+Nm541aCN9jeKJnBPNCZUac3nZIt4zuthwi9JsZ
x3MYDCsBV1ydOYEGEI6Ln2TePrH3WiFQrF9IudZRMcofQB0MaeLqXqHGuu4QghTjgaMH2GKlQ7h1
pOxI4sz0NgrTnVkEG21ijiSl4rujnM1v0Mexn/hua+mg2UHy6O8g6rL5dOFYIFYw5pfw8toFLG67
70HRukQSy6qyLdr4GXHJn3GBvvHlYKO24LCvSKPK7Nu3HmjN/udjXIFIBxudr4jrgjkDncqPZPWJ
bf53w0GqMt02DSgCd436AK3PQdzvPUg7m7Cpwvd5uOIB4pUzRpzzCV8Zlt/VAIDrHvpl/FfdlddH
XpDmhflKaq3tX5aCwo8IIBYec7xDlh7LN/R3ts9lBHwSzc/gwDJFvColmEu9hCraPwcf7Q4cLbI2
NMHTXqYcHhX0bkYXF048O2wWW6ezMlGI51AIumYS1XAe5VTbM4NUB+N2JUAN84odb6+5bt6neSWI
wRIu9LDp4Vir0Uz1odmmhL0St7ElDvQELDtFyd6X10J9uuU9R4yCuHznYiAmaQ8JznE06uulf24L
anED7D5W8ESj/D4BuZ/0YEfIfFYErJsd2CIvcdKN/I/q5Mw5IbDdh6MaP+uqYyFyfAMWHqyfVkNM
xvIqCXS2m69An1nOZRku3D6SRhzx8uVqt15pvTOoXx3G+NkAZ4ZeoxTMxO+jiRMIS75nNNZNa248
7Ph/jQkzl21d/MNN8GbCWR/61suVgCJrIsJBMsOpRClJgkDMRpZwlAu9ls+PJp/qZIE1uOlmqfGm
Cen3dqYTyYeAGLXgAXlw/zkrb7RnXbavYUOGVsU9arEVYig29OYijLAbEZjqwWG1qmlpXeqtmc1J
DqrbzAzPyoqa2Nc0KaMtBmQ9FApXuLIP0iXNKy4o9XN8pFakUkO4Hw3WnmjpfMZzENImyPZwyc9+
kk9N/jCopnFMfRJ3DQk7N+zwRI0Qzw99M3dXShWE/2eK1GAXHHcoq2jyDZyEKQzndgnznOM6CgZp
t8Sl2SPpyLUxXDCuXY4X7zoof/AR33tRcTHGQWvJ6V4bq3d7yho7IfLr32q/JPw2G9aLxIo6/Oba
q8FkWDzuq8sAoazTKzAw0Aio7HX7JQ3BvqsPX+y0oSg8UlyIDK2v/o2UhsyiCegXnofOC1MGwqOS
Ip3sVoxxm/Sk0ie+s074+NupAU+Yhc4gMpO9XJb0Tp0i+xb+iNknqoVRAy57KA8akDS74TZUu1c5
smyQ60K0caomNf2xjuKgzRI/4VPwnrBY7rPLBXgUdNV7fJLz3PA9NZDnHaiF/Qq2HpgDa0wQk/9v
Yf1K86T+2LHRDYHFMmvTM1TiiOBMrDgXwrnlUt+gEykSQndLTMcNDzNEUIxz+ADGDskpKsJNpINs
nkxoekvpbVHuXFXkVOC8tr7OE1q2sDLAyOjlBU1DVOUkgBXBWdlULYKhBCfYfvR9jglR+haCezVW
2KcGkQQdRsIeKSCdSN9+oEnz9S7EhL1TiaDOazb3KyeY0THcANOmFA2dKtrdAMMuPZjTzmzvcXa0
eIrSH67JfMdA6iX9eO2403hnMeO+q/etO7ubU9CikxCitAGeux7oi25n9RAAxU4okNEWneyb9m6w
lanZuZI4lwZaMCaI6VUejOStLe/yT56l8gTdVsFf+YlafLDgHg3r1fSAoadS6MnhQ+uZe0xdPyb0
RMO8kADf8VFpTIG0nsMDorQSMAxIfycOJnRjLtFGpNQaDfvanQwhPMaKZxRAkM7o+VJPsaTWyzD+
m0nGgfX0rRb2Mq8v+m6hLB29nh1qmfQOOlkl+nVvjwcVZxISQK/nrUVaDnn9f+3YqGrE24Aaqd/u
8648MTyv+LYUfnfTi5wnpWAdLFdN21sJXXFY/0APWUCI3QxJyw8qu3j9YqvJq6Djcf/DEqwLjVc7
Gz5FzLP5Mz/817zHR/76JBW2bL3/q5ZBdBqO5Ks2xaOkaqQiug7i8iJT9VL/9W4neJKix4XzTSUz
Z08kcwAhXmwnSHb2tEIp4XLVsJxZYarzpbrefeVzaQY8IWBtRIMVlXNDwbZuuhFsK68Q4h8hdbeB
69qjo8ZNOE+jo7QEHatN6lEBKzVjxPq0fqIB+ZvUg9WIqNMuN6QKi7yK1B8buagNfRZHI4UN6pHb
Fb2O2qBBbJ9NFtCV3mTKsivPjxz5aPOBHM2RJ8QrGMplj9N23ibBXGfUL573YIjsZ+Wi+reRhNMF
mWNvAs/1v2Axo/7BpsUkonXZVk2AkYIg2QehunGetDM6vLkc5h2PGGr7VckedO8huK/QRh6j1YFJ
LAmT3thFyhVXCzNHiT6L46sS5E8HSey0yWhu4up93tyLKHAtNEI7/nrUkWnSEV3ge/p5fE+/gddW
BGuVX9UFSK8VKvtCVpKxNjQ/KQo/KidpVce3E6q45D8slxmjNTxczyF3Qnmizd8eEzHpgASRexL6
yghZTTwy0N1FspeSYkdNw5DpoK4jTAiPaaZuzAltx5TF66QXOlsUI1Qb34zgtsdc56TLKbYnlV5/
XKsUh4a9Rnwowfh0bkqxQnSYN4aFEWfege+7KF0frG6AGPbs/2zRKR/VvQX+J9JgQnFEku8KNwKx
BMimxeUCTQcPZNuVD8spuOzqqpOT0JQY/nPqPFhl99Gk829BN+30kveZ+KBZgt0Ebcoj0wwf2vVC
GgHXo47HDNrF6hBd6bHKG3JofnJoMekUozGfZLkx7w2gZNagozIcEs7uWRy9AtkpgjcHnrx2rUVz
rhrG5rOwnVt0BHoDwIiFt/+tjXQla7bfvtThXXlcdqysJs5u9P8fZLjQcYytXezAEA5x4iUVppRi
cg2gntAnyEmIFB7Zf+wmXXHbogSc1Ip4SqY7lsIUcOEq6uVVfmSSLlkqCosgpjk9byhVgPtPuR1U
7c6w4SA1oBUMJtZVOm7DlF/ixTEp7QNhWwit3P7wB8F1jf5zZ/FJdM79kwj5VKMxO9BpGnq+VP9u
C1+5Hy9rxqu8QpQoTmMiRxm5IWICDrhmnjqpTezWgG+OP6LniUbrm6xK/FlvL0IKJNVGHO0J9IOY
MK/1LZw3vgeo27KIn7C3zsR0MJFjSqHuPXrjLfOhtz8WPid/SQe4Hf+Wu+ge7CoAK0tF8oQUW7HC
pr4Beq57kzXfzEA/zTTQObwIlUJINA/ZjPOOYTpTaL+/EBw0v3931YPVL/3bRr+dPe3SZw0IRLY6
ZDEZq2QA13VRpB39gw0DzNXbxIsnEGj9qBlt4oceFKpVcKsgpTbKi+IdPhx3sZ2RJtF59mNJlFsG
AetV9nmlcFqYbVDhkfZPVh8jVkjPJBbPl6ocrETUQrTgGk8aPp5XCFRA/vG27+9FJ3mDWjv4eC5M
t6szUG1LxA4cXGibePYt9ky7YGhPkR2Y/I3G9qn/0vpNwjwQXxDi7yBfsKezDTmlU0dayaM4L57a
Lh1Hy4SYmM/OJdLvYW9vN5fFWw0YRoxHdDobx+Q7KWR0K2/r50s+crrnHDD4YqQorPxOadHWwMe9
QezCYv7E3jjfwEW7ApxD2imV//0kpwEO3fYtcHxOEk+xoPfoJOWn/G9cJKpi1VU+JNOccPY6XvVO
vPxogSb6pioTXancYf77l/enbLZsx+DHvwVukn3NXAlAqLbmDcJ9oRJjosxqRrKBDPRaRbTkponm
di6RZ7Tk/hbGaOXK+zkE8z8rxicv+oqiQQRQhH+Q5j8rjcC94/E51NsTMSON3VSb7DF1UNuG5z8V
ZYVeMt3w+u4zkAo1MABHCg9sLm+y2j00pVp7zgnMAimBjfocvnBB6geLf8l+WCSJ1RyxUKwYSnHu
N+eJbmsMCWi+FBPB1Auo8gt8IGqEkoJoH7JST2prsEfStUTlwKJ3H98QIBTsPUj959Gn39ASNazs
xNIhnd4RjVi8PviYl2pdOSXxPMT4cy+j0g+v6qPfMQiUtzhnjglIxPkSekkf5Px9mF9wyI+E6jBz
U9JnRHxumN0r+IsT31t9l3QS/3gCoDACER2CFqs8KiJ+r9FicClOx0edclpSIZfJfZItF0l+Sa5g
2EpS7B3uEvYpSKTWaOoOHxiCtcTsQfk2hwk782ulbFN5NuEt/GDV4Zl9vSCPNm3BIwvxPkfpUlCK
1qN66XifQhvBj3SOg1JVL73mILMW+EON/0eiUFvNlqp0LXgPAoSUt3YR69bgGtzo52vh1ahsDCQR
amr3h160MaeSXingW7PsnvmyZzmUoSVbwSkuVA9XHbTWEbMQKK2hwHBtO4pubbRJqF6NVEA0cfVt
ZyUxch2cRwvG8UclbtGR+17NOCGzGljjzhUeB58F9VqboWYDImRTA2bfPaVQYsV8vzzhtsgrDuwx
Eb04vVoPz4OPKtXlwBkkCw2lYcK2EkGtpd2ULUKhuUiYwhUYPL/qoJfTtqIcn7cxoPLX8vifk7dc
neLvRihj2/B8uShzpMCIkykDdj2Vh8baht7brSd90p1p26gSuta2VKrvo2FrZFDHp1+8wozSjWSH
VnPBqwMc9xAu5WW93vNQcwW2pWWsHgdnyN2rMMLuS+zLyHWb5xDZxkD5pMK21pjE+FTat0GBa1K5
Mj866RcgOCVHbz7DQe/OT6tw5YdG6gneFRft+v+LpCVTbtEEnvIRFQgVq6NI6TZqc0eisDA6bw7d
pHtMrLxKuEKhHOw2Bvb0emkXXYGx3hmnq3c35NBWdppfZ5XwzMCvm+fL70PJCSMDGQYxfGSAnzPp
4Ww/ge5FQPdYxpVqYueL4Df17ID5mT00cBuDvUXq1H5En1QDxJyktcv2pkm35+PhF1sE1GeZPham
w9VTaz3GYK/n5Eht37aw21f7A9pO3KD08zssNPfkguZght3sIojcshdiGiH8aCm0SKq2KXrqDDR2
jOLXMJY68zua+Rwh+tQmBBlE65Tf2eG3MQ3EgH5pIW5X6DHNyDriG3wqDklKNCuunNcYiWHfuVZj
DJwj6rww8t0hfz380/09E+JE9VPyE/QH4Eqqo8S8UXu6w5cg6eAQKszLkjdrvgN/pkKYPzSCpkeU
+KOk23sJqEo9/pEaTslZWX9Rp9kiUG070MXmJEFqiehnFfzPluI4ob0eTR16TYQxWzfQDBMWeqD+
X09m3haIvgzHQwT8N61Lo+xWeVCTJekZvPrbwpnWjsKvXs6ygQA17IkfooWEX5wp/vTh89D5IZud
JyDZY0dkIiAhiyYx/T4+zz1t3z6MQLm5HT2MYtsyYIjo7UZwGri/xfMfualAs7EJwz6lAniH457F
29BddIIVlZtftHS9Xje6N3at6pKXu6EM+V7tWRuAyUShAUIkQ/P052njLXCaVqAbSXLc0Bqs8fbr
Oty6I5iZ6uZ7oHx98B1RPdAn1EsSkq3o+6WlhYZl1w0ZfbHSC3+kW2SngS1OQLN8R7jF0U4H6s1N
IDkZ7PPAiggFYSktMabRCcDwTcAoKDz5hYEOWJVPFXByDU8QVeRKiMPrdRIK5aIKsEciFMyQYNLC
BPFWSmeEZrshJ0y4ncGqABIkKwbHEAQ1kRZvEr2sbV5O2a0sF/bUctf4I7PujjF4hW+7Hp7voDcK
X0mfhz6sPVWblZA4MnEJzqz/fzbOMon7BUcJzPn2mmfsH/LqbK9pq9rBQgF8t8oVehD+ffyW0ejB
t7rOD3xfU6rvLh168pwb6lJtU9Q1ZNCgmv2QSwO1Vngh47F459Aggbg1s/ViciZGwL8bqul3UQ14
DVsa5qx7aAOTXvkJtp3PLDrAfhrTqlpIEn4uw/OcLdTUuS6KtPFuGMLLAId6Txjh/LHKmCfhVBEK
gvkREcXfoZWFr9tw41pcME25+XBXwd/zP44eA/mTXWviPba7BwYZzA1+Ap+jueQm/ne5MTGaQNhy
LGl4OQNFiGB0FKdsZJd8+SKEz4t1ywl6ayWe7lw6qqdGHtN3i2NN3ik5T/0TxHWqszLTjwhOuPO0
L/Uj0u3QQJqjsS0d5X14xvKWcuRyBXSjkbF3R6nIfaA0LdHSJb26ur3SiGmL0s85IXvCpgsE7fIs
4Rlhsdscu65AazwFsBTvWngNaj0+FxF+XTCOYnSyFP7MUTnAMoIXO6MhLELIkglSo10S9Jaq582C
/dg5m8IaKgoVvPgOo4nGE+WrQpUd81SQ8phSqk5bk8gf3mOMNBhklF7mPLDjDSWUNCjohdaIQNma
zs0WCX92aM/V/4hy7B3sKOynu2jnihHMCU0oPE31+KMGfGFFeQ4ntkTq8ZzWCNajTqF6ooOLdlOm
OnWymT7hu0FdGHnfDDKjBBofNWQ8MdYwp7gXJNhpsudYZHomAjSkHwhPIkFsINMbRXYT6YbNx7cb
8ugPAcagJiGJytrDf/fv9lttN9vE/sgW4YeosJAPNfnqrnpR+S98Ng3P9neD9j3q0vA0nBlNoXIH
Yvsh7sowaQFM7W/x3UTiSQp7bFPhw+/2Vj2GQ3jRTfUmS7wKwkEtiEA90M0FrWaOaQ4hY7YA9IiK
XDZ9aQzensOM77Xtme2txuy8DiOXOXcd5ak6TlAGvma7nxDYqpZeSEi6/OOcR9RPUVObLHVRhPQ3
w/HsabwJdxY1bMfypxGJwObNL978YVwGjSu87jNaYuEju8zWNHqn+yM/94aXTe1t+2rxmVmPMQvU
v9RLT5mSw5Uu4M4mWY2vqdekhQHLICgKhjmWio9grWoyfGXw9/68J6NjVa8cBzYdu5/eSAmoBRpz
7o/DkY5fGYS8ikeKnBjQrWIHCYa1e2q42pPd2Kq3m2sUS3pS8zvjBlDSDdvfHxAAACLCjHohgpGB
7LhymWuH35jRIJ5Jrr55hDW/W8jXiAIhaVZX2JW4rSS92TLx3GhWU9kEmK0eNQin00+jzHW1P/4A
D5T+kf3DuSv1kFzKXiZ3/xBTFEsmAK5qO9Xwc/KLJZt41pCBGJPry6bnXEyRtrZhzFwvUwApZFYA
Ehku04oDuxWlZXrVV2ohpzNXPoElYbt+m2/LCojG0lEKWhBygCsLrrmRruCeHLCRIWyJ+RuW4BMi
/izFCyH9DsiCfOS8wBymX44KuSswcCnFPBExUtpNFi7sCbfdM4IkoDxPssjiMnpWIP81DoCwk0zm
5M6lLHDKSTm6jZfUUgwt1IMFTgnYll8pvAgOCl3YoQ5oAnrrUd12SZNYdVwtZAmpAAzdNJMDjuJF
R78XAc1eOkU+HBNSXbIbPRhhMQD9LlGCLuaXNGKFMSrBXx7QvrQoWrn72LIOSYNR//4GbxRjXkCR
vrU8PdztLiRZBd669wujMguyrOtf6wmfK67rH/G8GEf1BESi+OkSwLZtj0gFmoYe8As4GmJo4myQ
RfAAaSl3C9JVQalBel6WgqS/ss8PYBMlXBPssohxcRMS7yVNciEHqvgP+55uyd7gBWQx5nddD7m+
mzrEqjRHtGjCCsr5b5v6rMEA081vdh/pZXW9E1z7B4LCsYElI3u+aMs61o56iJBKgxh21T19ms+O
WQzzKR4rA4wu3HH0/64fDCF6q7Vap3gCP9mhGpm6FoOjqhXoBAusuhSLoxmSqa/AkyaOOJaJMoH2
Lse6eKGoi2SIrpx2he/oLpebJIY/H80xI597Fqsu907aIkapvOEb1cxIyeZU64OP0FLRjeo174nk
8QUSqnKA8PlykrMAg1PrMekyZ2J22Kemds+KzKMlNF/OJRcxu9XV7KfSM/NahP4kUiA26EXPRcUM
toR4aQ3Xobh+rNYeaC7nOec4/B/1Zq/929Jsdlt5LHo5BblIdtKB0KMV6/BqqcTguxqoibWDYeEZ
QUNI1mjC2vrRrHAntoUq1Zfqwrd99FGPA+1EMjIjNiKCKkU64AC+ZirNISi+A42jjqZlMzdC2ikm
Zhrgk6SCphKtuP4aIoHUPUjOp/OgqoPct+q+M2iaN8cX8cugPRixGA52OpBz+LUFkFf+Bv7uKAzg
c+UHdq9iSTlk5HkREVgR9HbWu4X8a5ZZEJvsRev2ml+yCj5h3ZXaAGBkave7jT3Ww0a8Bkr49OLy
WkC2BSwWr6RNqTKEOnVKiTTNPgjMfSLwuNOMXz3qaf/Hzs1GsgAlzxMGR3UcOATk2vupcKeED5R4
eGcCDbr0zZsfuuBlBec/7jLW8+voN5xrHki6Wgr9g44ktn/2gED6ebL+tSnBWH+kyNlWxd1f5IXO
GKloZ1nnU4IvINkxa9231AaQl7tSCr/AyXGIG+aUPNEm1e5gYO+H4yl1kXkNLCtkyCvH6LoXf2Rh
fbpyeJZEi1FF3QJ5quEeHZRVmVY4kFdz8ipH1MSRSunAadHx0sg7ZuyAzGQNUPWAMbw+aW5AJQVk
qQcESH5zpVKpm2VWmUZ3HztVsgnd54OevcFOTAXzJDy9FSSOfcvo5gf3xl2XnnBlVIc12Wdr4lzO
RDb7hRBDioWSp0czblvpteHJ4gSi3sdbHZLTXOR5i5rm8jzMVq7bnB06gDR1DLOD3jWAk44ti012
ZlT6EPXn6oRgE7Zelzc1124qGmPWSPc2vMn+kl9R3/g72LgDvOXsjejVK5VF5J7ufkhv6Mtsa70q
1Ck5zxpcY6OM2Q9e+2ow0x94xg4RJRpdu+5vXH7G5aOZ+cLYZqpLQUMxviSrnfIgRp10M3yZoV0Z
oUFmTugpTtoPUawfoxFk6Kbm/CDePzkuXbD0J93CYfXpuOJ0SQBA/+CLQtVTBwhviLR8u90UEcgs
Z6JidQJ9pRN+1rhkz3xormP7Y9sD8lF4pIx84v2OSnxPBU4BknCqlQChRY7ycKbxF03MM9ADjdk9
Zty/UUsHS2gvptTHvZvsYqUBZmAiYvYyJAU6fQsOj1mmi6SjJRLfU8PzTNTR1GmL64aOj562QLJJ
UW08ZdQ/s7NJHKM5yYw3PYcVSkwoy7ap3Qvw0GelWEmW4OGSP+IDwaC7f6eMuM81uaNxESMuapzO
CUvuvfFw3mS+DZ6fcRhkpCCcVAl2LiGNQdL0Aw3FZSXCudRwbJug/oiKetETjFTaCOxriQWiJqAI
L4myWsheAI4ST0miEeoiK5ie9kp1docrrBs4oDUovzyj9LXeVRd6wDTbhuS4Z613009Ie8c4vmwK
7cNYdl04vgOJguCDuloVaz8SzuofbaS1IRufNw0YgaNwfCoIuETt45QzMEjs7ziVhdRVnCuzunRV
HEU8wXFF/fzw3HzONu/qGd/GQrjamOF/i9V5qFEBtFc+2mvqUCVtKG0xi43sfabGL+5cCiow1Hn2
lNqQ91fbJ3/g4y8zvhpCjiusxn6rUeJWJnwCqP0dK4b8QslxXEWc4aJDmUMCwOfz/mXSMwU3uZ1b
IZ3pB28HGKH6TXTJKAPXrLxIxGgTRT+NNDnmct232n8DF/kIbKRHEKZJ1tWz+7ea2fLWyOjNjekE
iToDNIJtB2xYckCrg8lTl9RKgjGvbge4bcB3dIl7ebHqRXER8Xc4Tk4i7zZlM8hnZPV+X01H0SEn
B7bsIfHYiiE/qP8JjASB/tYftHTMa1ze9lMNOSLDcar/Y2bfJeL/7Y3FJuNvma5VseswSRUC0GKr
Mdcg/AU5Ouq89L/Fxg8dJx15/fT/RQhV6UDEMXgP6D4M1AS9gd8wPYHRdUSHfcN5a3IKoFrEWdIM
BJSxoc8xNZQbRuwse1WrmvZCQXfEewtPYDNJDeNjPw9A88Q6f+kVpeFHAucjLN0zAv1hFhmz8Bv1
URrC0hjYPsQstX+MX/pPj2txfn2W50Vl3uf7d46dwI+/E5f2Qo0rnuLzkXbAYCLyRaTNFQTCJrR0
DTX3OzTpu+G9k7UKow+WtgwbTGuFHdGdOwwfxZLmAaelTKlbN15mG5KVXkKAODfOQjL+OL94vW0C
oiM8E6gfn9tBWxj/cAh+uLUs+2Uedy3R/m4IBMj9hOlJcBzqsq6g9AQeTFyXWb+T43NeaYT8yi+0
PT8Fx0nS/TKGML5/gcLnjog3ojU6D91xrHyEcu88jLtxi4pMXQpRe8oymwVpCOBswgCriVt2uMoH
Ca6aXcp2nrkLwVbOKDrdBjUK8Jq5/6UbN+4tNsGJx966mAKNUdOcCUGxk3AsQD0/kj2AFN9jkaQb
gf1Su1W++pjzCY7H70HQYlNXN6+ru8H38Z8Ce7fjtjs/l2sa7UvIRNqixpGai+VeOuB02FFIw/g4
y7Hg5pWr9/+9JExzfL0OovjegECH2NKeEBpNrZ/tSRobjFSrpW3YySyxmhONElFNBUffNaG4L9wT
c+/TFOsOuvITUqx1i9J5bCY4iKhDkZ/7JVkMxPoA9n06PIDLQc5g511FNL8sCwzOVSziLqdUwzyS
rQTcv4NAHYqpOvkerW6dvOtz4p8SeqlfHL3rL8Tac6fRT4AJXBKozNYPQYu37mZBjurfEU5QofF1
QwxMidzY4v4+FzHJ0Do7fEeN42C7Q4g5icAUiy9gimanVdWH69LCYjGJqdoRkb8RruY4ztXVB7JV
SrUkFgmnXh9M2TAKRzB76KrUlSAtBl6wezJMUpQgiF13VcQte77U9tsMVJTDzVWE7sj7e2hJZB2d
mx5faDV9T7qSIw9En5ksHfh69WROoeeeEaK1LUNEtbfDbgjhF/TrtOMpWO1KQrHhHIp3cjqKUyZB
xGNSotvsW5LyQjAZw87DPdblUhnvQ5N6frPSxyVfmTQ0B78uwLdVggeJAJbzXdtmMIQeI7bcNP8q
WF93D9HMxXYuzKP+L+QPGMcqjUaUb2bjDWG4AL7Z+P83oXt9S3aJ/d2ow2/K8cSAoyvanho/RxjC
+ESzfhYrPdpYsAnJ2obSc018zgODjIR1fmysfi1dE94VweL7GrJW7mohXLWidEteAwTsfNDpacIF
58v8Z8B1ZASUbaVNXXEsudnTFR0V7pDeeOsZhPd7oHQfN741c/dIEwxmZD9tOYNqXRJ+MUN32IIf
OFGG8O2hasarY7cXpCMWrVEK4e+gwgNHueptjAHz8qzRTgkLY0MhI/w8ZPIpzKkIrZPPctzDIJrd
baY+siiVmy1v+bUzd0Pj+FdRlp4QnvIJBv9rjXNBmZtr6dgaAQWRs1bnuzjawmG0QE4TGdDHQ8y0
UJQL0bZ7SBByKYe/sTvcCW3hbNDBBpkGp9w0phWvXyO30aRTKCjXC4Ib2T3heZE4P8F7RzCU34o9
b+Lc3bW6CjONK+lzpaR9v+aSYAbLcc6iI2PZfQIUwZ7EsKRhcMrbuxoJz4HYU8KEM56DUsp9A6Qa
1EhiEGNknrLvnCSDhv4NduMaZa19j5tiBlAYBRIvEugYSf2UYmcEtlmYRhQKqvws3uIMeZ8qqsUF
2i5NBopVOTaagSqKODHsfLARNR9H+HYcnhMzt9+4kpZ10yzBb+4b2BtDXsffv83fyl7QzDF9YHxi
HjPTW6iqdK67qQBC2FPvg0rMO+1ZJvXuqWv064ovylgUDCTiJfkfbL2M6ftgBcsZsU5pH2RjorB5
J8dk7vdgo/slB6CpLspNYMcjo5fua8RIysJAzd+apMC0vSkoKb/iKS603C64u8wOY0zi20vwTIw0
9UyzXDhuqswIB+hya2ez1vYeJvYproOlstDLRPPS2g+8FKVbNRSEfVrur81l3gg/U9InWgWz+/rS
4iTGxmYYWh68/ib2KhFe48n24lbKDoWl8oUVeLALRFXNexTU+0U4g916zLZwp0dDaHW0GoELYMuR
3VB3+cXgwfro88IfqTcgKygUWGD+M/eQLcn9gv2Bfiw0fSLfp6p4Z7Qxu7ldS4MLRPxQxzz0FhFk
vtICp6/zT9Gjz8f1WLT0ty4wfPVNburvfbAFm8eGvFF5hNcDeaYi5wxnW5NbvdixPOauMsVZ5iAR
3bGTBps90qK1TVlNhKjN5JYGFqFW7Xy1KpN8AyxXyupIOwzJaKwRSpQABWUY5ib4fAWREUg0lyVv
OqJ5gHW13ujJyG6IOfdtmYLq/dAC7cMn2g2oGOP6GPq3wI4NatdoD4FHtTQonxTi3loqtwi0GfoK
p+hCcJkKimSrVycG2zLQJ5oIPfHVDCyOwuhREMRk2iYJCdos/Lvkc2tMAQEZDVFWFBt95R57uBGx
OVC64N/Uzv4KP+5si62i51OU+GuAsGsbpsL8/laMgGXBMscacTyOg6CmK14t3EBx/dxcQiBe46Ew
8HZfkBHng3qdQQwxV8J9v9EOCSCTUOwO1ZU0NMOSAn2jBcv08m4qq81Xx/bpYx4vfNn20cG2/s5y
ecJRaibC4Sk/8NeoVzA4UpM9ElfzrbAGv/mit5SuByij++/h6clX76cyHQZSNZ6AAhxxzwfa6XcB
Yk6miKl/rgk/CRz25WKQe3jiP2sgaSP7+UCJ7COpmQ5KYq2JL2Q8jfKGQsDec7eKoZlcS9s0GfW2
p3Ec6MyjTicNL7dRlfdcdJRogdmBAuHI8Nxrl8a6HDsTDkJBhdaW4Kqt+DQMh1vKwlI0aue90EvR
roIps9W/qCrkAwTo4K4ssOzvk2hILFoC4qIiO0Y3dmDZLON7gjNINQPMlphwdOW60vIzxJodliQ+
ASpBeH4zFT5TL37O4PZj6rdw7R4vtISDWzu5qYEOOq0hrC7LCyXXcjl0OGSeEFcUuO5/qHuZq56Q
XqNFJJP2/Xvtw91oeejo9MPL8ypSMvP4Ir/uA1IK9XcmafzbNP0XIpqIdfT8YQgGfOIkoIiRxSnJ
OWc1imnl+1uHUmZu3mJxkblT2o1/2TwbgYM5qeXMB/+BR+WbrBfYnqhWNn8lx373SAOggvyIy8kC
hXwY02kPdM22v6IRiZb0OfXGtw5SOzq+e4IdggHrXX0xn7gIB1JvGa9wKzJml6mriHzt19K7Uq2r
+UJpk8LJ1++Iv0OR36Vqq6J0rrcG3tXG8l/A1F5XbAkgTonDXNYMFFBbvzsduMkDd6548WIqzALu
w7lMAyVpEzV1oLYGw3bBUqaDrN6qeD8xwO0P45Vl9ua0hEfSRot5lGxkJfF133+7jXW5hdc6kqVM
cTb8bR6lpuCxHzpoXgnRT7uaMzoGNk1gOntBp0TFcgAAEv1s1FVk7lJwMIJ7NBQ5fjqf9my9wjSg
U+4rIEAFWT3VuwSQ72K3jW4ydOUZiMJJtfZ+aXgsu12fFkb2SyDHyfQQUpoqivwK7P/5mSbJW0s9
EjBriueeoibvr6v70zklZYx8Y1lvyMfADxsy2W5KpCrcV2zmRAmoolROxn8oSaysgzushfPu2kah
3T20oki4yPc1Zado3UedlVkUF2Qz2fUAjR1J08gtRsJyIejZHWkYftDwBmAIP9ERlo5/Szj6rm0r
ndaB6UwKMGu0wOtvKaO0UBgZC0nbLfapWk+t3bYc7mkuVt8iJP8vE93+c0MFQmgcQvMyDnFdZLMk
OhYKQk84D3MSEP+cWjmgZRziOIqBH8mCNvdlbHYKHCBpFvDQ2k5CwzhzuENotFmDMqLG4nrn4+i2
4ytyL3IkTCECNTVj3jfbGTlPkkF8c803Cp966aUCpl71G22ipNBi4Ir+dGkPrb+BE3vccnf4IjO5
PF2tS0gbjQwdrqfleQX6g6gH/7PEA+LE8zMQ/3NJ9q6h3+s/7doHgUQpqupWTao1mAMSltvgOteQ
TKDvyrEWmuQZBK8H4d3Y8+W9ab4mFlsiI4nQYKssDELtM/QSGGdfmUAoC8V/xD6IOyAhb0ZMaods
TrqyszCyQrXmT5dTmlwSvDifsDnya0RDH4VdTMbOeUe6FazV8gD41diLAtRheHl5PkfjzttZa3wD
TyHrk1MBP5+jw4LmFUkQtn/KvMARTGNHsy6iCmh90ip1KN7Q71lCXJ9p4r8+VTEji1T7yVvHQUxa
PYz4KC0jMdfgnc7GlKNrOwwWAe2Jv21/tWtNRFvEB6QxoaJYorAuzfKhmew5gpTmPxi7h48Gjz7F
OituehFCOu08WZcux9g/tZ5/QKUR4nbyoZNMoyVl3SNr7Sd/tzH3si7YjYOWj1c1hC6TJGGkhyL3
wndkuuHCx84kMwejSI00y4EnlmOJs35UlgKcT+w0ecNI7C8eX4yU6fwOAggpEeQRkCUvnYF/kTz+
L9xa5M9qen1I2ZcdGe/GWeXaDK8/BPP2MVM9DovLLkxpbxtkVxwOSV29L59PKGuQUizJ6jhOXx+T
ghGaiL+OneMsCTgBHhDBXPxoaTHL3XxmUFa1cHCr2QV93qaCDqYIwpxl+qysBN7oRLKiuCbdvsyx
sKUv6qzM3hRqgpXA7lpzqB7ld7EzEvgeO8LPKJTv2y+sGCj3rODMSSuxwhNGcKrB9yCwM13OdFdE
iX89zT0UKgPKe6rvQV6NGgM5JMTtKoyihgtXiP1oSE23Zv/WcuSmB++RlxOG2rjHeHqzPzG301Tb
8RdwcIzYMGuWbgJvk5zkMSQbQtrsW/MuNLgx0KESjr0jm2IRQGwIPRE9vanxtsLZp60Eb91tQYp3
2P6Zj67Ig2c9svNmjRtcYn4QkyJBCgLJrWFcfM389MPIjO1R3Sld404G1APSUkahlL+RAVDJo5p0
brN/TfuuiTioFz+IkAV+5dHv6wtcuA1vEs0aUJ7V/khcXF47DqEXxcAuvabF1itvjANpJkWzB/P8
82l3xlznSvuLG6ZOYXNs9YUlB0a8skDDB2yyM4UTe7PGxZjIr2QY1+log/L1Ci3xK9xjLXb5z7k1
ctJ9n82RHq7hqSCV5gP5P9C2sRy3dmnHn+9+vuAQ8XR8JYzwh/keXSDnHLXe6r9S3s6659nJQCxD
kpWFGF52YPHEfTg1hkRhlDCxP/uLFcXm2tMHgqj/w3lyIr5+7mnHb/U/yFyesgh4mh7AinvJVuIY
deYyEchMGKxiSGsK6hSNye+BcOxR9RZsTJ31/eVQSWgATdP6ppPJkhCPJezwwOGo/3DdfZX722Y6
DpZcye9E2sBe6jeMB1zE73j9MOpWD3JB68YNGmbsqBooclqkxjBqy3MG5Ov3XtWdMA/QeHdbmk1N
Vw8b1z+8hsW3stJNTq5jEqQimtqG7dOXofG+Qg9SouztZ/sje9r/muo1Zdkm86Mk8YNuhZoiApxY
mZrnMjlEaexs1YNIdhb2x0qBRekevDAmVHDbIGwVNlOn5Q6Q3jvpeenhQFyioHncR3us8VSvhzqq
6JfA0WaIHNlseCksMhmNeceDmEZIw1cQson43YQQQDlWc4VMZcDGWzulpiOozDpxDG4n3lI0hZtX
9ZCnNcFFfyNUSo7dmpWjMkpcXBgLxIKoG/eIcat9YhkquisOkIi+3NHfGq6F4c40p1Swf4qFfzsW
hWHvJmz9gmgputXnC+AxqZGN6g/8bXXBzCTAf5SfuGtq4Ndk3Mi1HltShWQPeHTpgpJbxihQGmUJ
OM95KohQ3D/nlf2cQF02r771DUr/DfRdVjejXCuvocoBGNgUlwGk/H3/+YxN87AoKnqXABRcGoDK
wA9NqEzj43Bh18yqlcZD4uNhRlqj2YUJgv148mnVTxD1EzuBs4qJcvZInDpdbqlL5SOYMI65y73T
e0eHezXD5hlHdlg13oHwA7JUnpXLuhHNdzeF3aI+1PdOjRSjrvrtJpjtwUq7C44DTeSpKyFBiuGD
W+B3RUx2S9FmjrLrBybqwpLaiHNbev19uzcbOOMbFQAalY+91xfBnuPbD8/q76kj1GLAYgX7xnsI
xzdJRkZK4P9jZvOrBm27EbVHaCMYM2ybPZ8VzpI9n0aDJFUnt5dP9cgE5N/bWuH113+wEP+ylN0e
lCWSOomudhvYN6LC3wZhX9/pHjhUPOzsGDIIxP6X3a5mr+KGyjJqZJE4GPAJfqqiCK3T1YR9ESmW
mr37XYZGS64093mbCyw1Mj2BbdLIDZ0XDW1X61UREY2E8KqT7qXoGOpa3HE/maOFKLbkhQ7GKWDr
sCPvr7t7BUwhMFTvu6OCrVOEjsKe6PkVhHe79kVBVXOUizmAETFQoZIinDRGFa05WOAQrNKm/Xcg
qLYErdkuwe6jVG3WmOmyE/RMM2uYtugSOcZmt1i7wRHvYEZeflZGy2H5sIkMDuskuqkF33QHLPyf
tbmzcS3ExC+QaWrapXlVCPgtPIzvoveVQAWyyXN455TW/BQGb2j4rERjvZ65DI/pM2Ium296UQlS
ryPj4bUXT1nzcIylCfsfGIrffcmfJHAMW5kcRqOaxjkSDhP/62OvFMJkRrWHTIVz22D0/CftjZ/Z
lKPAL/7JRjY46gAPSXD9taXCSwlzFigMAuwb0G1BPDWZ4CNcY92fTKWHVB6SGIPXVzCfKW6PfxI3
BdrX/T77U+WJzfod6kNaBSJ1BLYoAgaTM7gOrPHUceLuXy6hlWiCBfOnAQgkzvwjTXeknOtWLvMs
qhSK1WO/JxuGQ9armSC+GcFartilEjC6TCSS4W+JH8YnfIdjMWFZ9bG9KQDGbSk/70YoL08YqN6I
7SY3wSiVjZ4GrROWMVZhQ7OYZj8UraN564x3OVN70gfi1K9RmYSLcG4lVNM9qppdPvB8bixAMzhy
ExgnwRPLHABgj3cFu57cwX0Oo4ai/0QiVi9BgR0TlbazCm4tlEP77i5ITtRl4d8XBMC0L3iJdCha
EplM7wkk9l3i6wVZpkDk+oARQrEeLBFPTGNE3Y3hI5d/DuFXjpg+JNc9oA3AoM6zrk26J12p2JqN
yaiV0x6yODUqba/P6STvIAmammq/YnPUvMRBJS92o+0NE07OZCodG80yOR+Agvf3cefVPRMITU5T
o7iLHv6EZ/5VbKJq4+2La8N4pJRHkWLmGr7LYDfyjJTQkSAT72EllS3dOUfZHD/1vhPzKKrPTFvn
mzCZf+v2HZ7dEkm7VTcJ08pQxRzs1jFuCM+lRHRQkgFGZk3JdLZLx1WsMfU2Kck4DAnOtClrs5VT
uXoGQdtS5uhkqxCpfd7PhydVD4EHXmJCqS89jmY/QS7hx8Dgh+z9qv968wLK2KavGRLaCFOIZig8
x+BMK4XRyVJYpOCr3zZGjczNvT8JUzIrslRTY7DOaezrXfH0+1lQi4XlEUdM/ZkfPw9KqC1jX//G
x9/DE0wmGh3tw6speJRDiTrXlIzQgVwFA5u9uz8+/Nyt0KT1EaFQDFMRanOvNauBU/bDsIlox1R4
XjERY291Drnuik8jchhp7uwg/afYDf1Ho97eUP1xk0Phe2+vf8NUCd0Lm+ozSla4yMt+uUhA7O22
WX/lbM2dylKK5tQlZmN7BPDwuiXNVbsNjIfSfkVcQFLjIh6D74Uw2pdicdqbP3m5ee8P9f+YiHRc
ROPHtC+pLtbXBLHahtmD9MY8sb9sVQBcpZo1qq79LFk7xpenAO48zMYHt/XJz9vhXSHJEzWrsSOh
oLqKLo+4/Gc/npwZ4u/H6eM//V46dzZ3lt00ifEVqe/gPV+gMCtA+tv/R4YjTH+mwwoWcA2HmSQC
jhuLJkTP5T0wEw4cPKwjhRugu6Qf/SAaOZhf1AFrIuwzn1tlJ06se3CSGeuzj6ZbA3whii4I3j+R
/HOwh0CZZzdNsK47XNUWrQVIGLKGcBbC/CKb0+MOMIhYS4dlifRDvJPK1uE/3DoPx4+1r0z8CleB
H+v8DFht2wH/rSKLe16ZKQcf0sbE8ti818UDbBAFK1/AIdLq9EFp+gxd1KzhnLOZlB2pzT8hp1d3
Hk51e5dEA0uuTQNHDtvRCqECWpOpD5wzbUHk5/trAm0bU+6QjXKpgHxLUmrqn+77BBZRo3cDGIN3
tjU2LjZgpQy3SLOFLEkgtM8WIb/6DlRE+alONzsYKzrYWgoQsDLSnt9yDOUj4BwJ7Bc5FZt4BYAW
mrJKXNfCvJ0Ry1lWYdgIY9PUHQ6wSAwpXO6yO0hrFDogjUyUbjtpIHjweiKTi4oN6tRV9sV7M7OQ
FrLVEIKXOfUIpF1B7NZ+HpVsQQvCGFdfRo0O86ryyRQiwNZLK3h+PUUoSY14slTai2WtOqhA/nD7
v9pQBS3m+7A7UCM3JPALILn6z4fAZ5/Rr4/D/bczmiEHG2mPg1k/CbWfdMlKoYA4FvGBEswHrCTL
6q962G7DOeWzXnFagcuh/lx3NbiCWS6zI2wHXudz000fd65nCRLjh54RBGczRE1VnfVb4BhonGRU
kyLdeknbXjafhc518QT70UzTQ0MnGPmrCc6duJv6KMJPZ+tna1gNdBF/ky+IoMpGkU4atiAmxCuM
tqXnDCsbnsslCmXeoEF8Wxi5++yTvCUCmsuw0Jl6RHYp+CS28zhCpKqxXpZvLe+prhzsKzo2tn4N
bK6+uAuSz8e8HAioCx/VV/MQ44c4mDTpM9wg4HgZiQnukRwgd+GTeS1Gwxcgnhge/bcnn8vknxxK
U6ze3c0/Zb/k1TiYenSTpZ/YhrtNUnbUSO/Ruq0ylbkrHdx7IWwZYhhvzGy4lSUNqk/9Qr7Ez/0Y
yab8o9libu7+Ir6oqgSpoGJiA1clmqk+Ca+gxyBLNI0yozFF0ZfdXUU+Jc0qMi0RFziB5J7aM1eV
I89yI08xG3vc4MRb54Y+XFyPxcEFcgzxYdHwzeuxb88Z07c/UpgArnrvuerPCZTovq614lbA2rgX
ZEplUeqbOTZbEIytmaeJJwP+PB0KBjgSHpWXX//xdYUpr2o37QQe4xKG6uc5aVaqTrbMXJ5EQ+yz
mZCf1wYQQCF2QskinIDYoovSEpfAYuRTJBuRlqlJj2VAxEDixxY3Hz2jkVxjs5lDJuFP0eYkX3lt
YbQl/LYHKAzvUGJIiI3C7aD5AZ1/nBE5NxqBJRTjbGH16kgiQuJA6dlMoViljjFyc9eSB6sMgmJL
4QXeuM4n717C1qU/MjRpUZXWk7pggbNlbI9IVJwTAqt+TlBwJTE6xpgW+WMlUbJYhzfnWxzDRadC
3uN2FwTaMr1dJE2QDPgy2xFQxyXNwzSnz8IGt+nPBq6Yk8nPkIEAHs6j8SebtXAq1gA4wK27GRxt
iYdd1dOcRVTdjxEmp5qDy9K5V5kv7hxcbE4A3DYuME5I+JBDsjK/eCQ2egNxnBa54LHIh0x+edbh
PuWRpcG7Sd3LE9/XXw0vHt3GEKpAtZJAvame9tCxaDZZF12OTzduWhkXNyMm+nWQQWIHKsbfNdh2
NpY+gvystYf/SklYlZ5vhWffjgBJ3SUayb3qPBmIau7kVL/1AxI25oewW4TebQNB20Y56aXXAm5n
y5/ZK7J8xA+KzV+XWfWJKEkml5orj1VnaFZ0VHfFLXYXQuh29wkrg/FctVwzNSxu9HrLjomq5tyU
GYm+NfK2MltWua+jCd7nGO2bdnlCk0X1E4qQWCQydlwHY/83b3BF7F58ODyk2mcgoXtDAlGTmiyv
aEsrSz9Erp8VIOY2TJobapLQhXY8n7m8Kkr2yNC5iHIxVQQYDLjqPu6jmMfEqfscwXuufpwk/WhQ
MG9RSkXYPYBUsj6SAI0EQSKK9BC+jxs8JTqZeyTwT74ksbKAI0fvNBzyizYthSYQpipQx9L8oTKv
gy7sPX8drRNkB+Djp1zn9zVq8/fejMtVILGHQFAQCMGXzHNKWJUyQXo+IdFJ9VvWO+oBam4rOw/A
jcDSH+R7J4qIqtnpBaS3TUYUfdQQaKC51iEZgm1Pv/o6jK5Dk+Dl9tyks78J5ubuOJTj2NPE8Zs2
1kK6qK0sUXvJ/UDUtm3rrDTxKrewLadhDYLWWoHYkJdDo7ioFM6plnGMO6Om/jXTKt06XXgTa0Hd
rSnnf5T1ZVGlL7ppk8F5Hr3a2PG5qMLx0Sc37PQzse+UhS4qWH92pEG9PaLviLFbGfvI/ijtzNZK
rdSrluy94BvDCcq1ZESiSf2zqqgxv0HAaiR08nUhQOLmV89WkqMlT6UGBZJya77OLaoZHCMo8j6W
aa4/vuQewj6AhMPPrSrHz5R+y3j8aXTH6KkX1NOSoOAXoGvrVVUBTDB41jGBJbp/5FXLbLHDGDq3
Jzoadkbr9WDBqM3BAHwyFnhqmfMXn/+21/5pmyzp9e2wUWM3Bx7D44SYs1k7J64s2JtzMlMmU6aB
AK+TX+x12LltCFNGbG/U3BeRsP6u29iJd/SZBj+AWgdf+4U1qMgr02sGW0y0btXqQTB8ZwtDRhmM
uh9xjXpimAHFThJAAF2Rja2McGoL+nWoBJJ9txGDIX0IRHcIXHC/CU6V84JdulmuDdkUv7Yolg4p
+vmYUfZrWt7QNWhHf2Kq205m0yZkBCVuUgFGnUnzz4p+oinZGbHhYDpT/WHHaR3Vo1Id6cMbiSCY
+8QZ8CLubArEcw8IpdGzP86EptMRJ2GbkZjZyj8HKm6rImVnvTL2FW+NnUZQYgyXA9H7tg2ojttB
dO01IjI3V46TCmy9K7vhZyMCTPwoSblWvZ06wgJ0kdI88ME07VNYuaaDhjX26Z6//RK/rUEcgAG6
BnRH2K82O/KycKxat5T8GzXu3FsTP7jEQ6p6KyJ1FZwEIeMESXE/KwPLYfjYVu0ohgkAEMp4R5SO
Lwa41zr+CfB9Z/idHs/FKBBfU/B0v6IKn/En99z+yF9uZNZjJoC3ToXPkvHHbPrPL8j1sfNu/yTx
C0qkmWVUbRLGihJMWrgFqcJ5CtGU3pHP00PX5G9JoUKcwkcU1Ey87uWFAvaXkSswTY0Bd6yLaL3b
BKmTdzuWpP7CAXJ34bP0iB0K+X62R+W1+27V/3IUn9/c7OpNNqETQgcRQ2BTGdsbEPsQpxD8Tbdt
Q9SXnhVCVRgRGnjyawzXjtaHNFgrwD8lJ4EmO99tw4hBfECuMyQh7lXvTHriXthGeO+OKZfN6d9F
TuSRJj5y5DWhbNTtWfX+mSugToDDUKnUnLD+IfvXC4L+0CdqwOeg4We7rOMKVr0FKlgm8sBbVqoI
rx8Z5nnWHr6BkRnuyavQZxSK3ca0z8UQRuvsbxrL1jc2RNGD2fJlOPQqI73lvEN/GCfXJ7HNLlNg
IWdr5R9v8nFk3KZPnCh10WINJd/gg64cJBkFqYNBCeRk2guq75xVIEc+14W9xfvQC5Dw3eRqDl0u
4yhNuoYPDc+arpcmv6NOCcRLrqRCldZ6JLbJALwVxU4Gfu8Hb+fZdZGuM93YxgAmpRuKJhgHuKCh
4QBgFw75egO/a/peOVH0L9VicZaNLIFeJ/usMmnqojArrhB0cNaJ79Thx0Foca4x3nCNTwGNqhpg
hW9Y39KMxu+97gtsSItgt/DfiCsD68hL/ZzzRWYwHqID3qm2rhBn35VkC9SKLR0Ad3SlZjhiedWc
VedLJXa3jEeHLoDWTkMZzCEa12r0zfH4ogMYSNu6ei26kF2M5075YIRvRgBroKWsz5UvRdM3BBfW
dfYLvQFhyWStSOtkGsGCLPDDwjn4hI6ZiC8rRhjL+QaIZiLUwTZisA/EmYidZoibv7PJIXdiWBhH
un6YOYtA+2x06tFd2bCbsdlVwPjPO9EagSRD1aqNB2RiGvhAWVl+v/3+BsG4Q1paZ4PqHdk5x6bf
nkRNC8DQI7Ysl3JraWGrn/fJdJ1hND/BP9AXrmu4k6y4j3RcoJGXsAkUTwyheNl54dZOJ/vTqrLK
63UwXcXeRmiAX23r8UjneHmQZVCGuymi0ieixorAHdjKEJksHuh+mFHln0nFL/eaZBZ06R/CFHAp
M1LyF/t3aB14BVqJew2KPYU33ald2956sv3jmPJnSOO/8N08Uc/ddi/9geHN/X/aaCSPi0kmUEwj
AUD5TxbNaQcj3+ZK2Zpckryge62MIlrhbUXAwyX0cMnxuKbl68I7XYBhCv/vQ6v6AwO/oafjDmQu
YrAfyl5A0L3beNwiIJtZTpl50gQf+pc1k4Bh8/F//GkZKcLdxK5PpzMgTy1T4L/rXKvn9mAHlLm0
ERqPqZ5OYUIls4IpTA4ZsZ5ohl3Bt8I5Tgb0gtNwi8q4Dhe9lAwN0I3AsR6BOPJVpXqV+zWI+H6Y
oyvzHZ/9bNjmIPjgyeTxcvpVxloE0ZBae8YGFJQEBt5qBH+GxohN6vIJ/GxLLhjXRX8n9XQe9OHt
NZq5xV2zG4E7Bzgdrt8NL/wsOxFX7vGG8yes7PGatiJOjBgJImgEor84+o3Viw4b8jN8TpQR4CrI
t/XvLPvr1s7WC2Hzb5sf7CW6XSp2CCeOpLsv/LKGeEHNER+nCUHpSdmqFhYwK2L2zeYgCe2I5QEy
GdbsRZgnO0aBGyb1mG0mavP4GRAMo5eQNx7IVG3SMwOVKnfBTWoTYEQVMUHAo8pTrB/c9E75NY5w
5Bln47OIY8cyDlzm5+xN/+ZH6j7aXESmKpiArX6F0F0GPisEw6VokUyZGsl3HZB1OQCz3ergym3V
tdzQDwjzt9uVZiRp3gNpMGpgnaHDzbGGkkdQ7lABfGTXIN7CVdOxaEVZxYeXm+pLFTR8Hx1fdGEs
2smk8p1JDyGb0zuOZVE9id6X/UwWFpTm6pXuVlTgCk0aMLUfyml/zhGUnpvM1dqSscz0vCW3ckPe
EFo45U8C5M9c8YQwSGKEjuSWGi8SqFpKsG+kt0PS7YzY95jWizZvbtjKjJHc7xPwDWjmMm156aUg
2lrhdWG/eEeRxMoyF/ztkd5HiZj4WYldUaWu9Sc+pHVI521UfAQDJaUO7iPuhU7yrI78nKhaDzUl
ay8cPGbAUhwJoDy/AkUkeSRh4CYfHdS9VCoj/YZAVqJU/G57ZX6zFlWgSw4AOviOulZCnEp4eNKS
wUQjoF0pqcGI7afiUwevqH+T5MfAU2l6o5YypSBHtbk40lkg/s2zDN7f6S5zUbTY3+rJTjmXOcpM
o1wxU3P55Y0uAXq9PxmkgHVQnPHQzqF8jYcx7wVijUJOiwv54tjQ00N/gxqSlo2V2MECNCLfmntv
QEEubZCvZqO9A6Ir8EvC0xv2OTS8V3FjsmKxqMj66pRBPsUP379LSSKZmzf539IujhjWkQokLBW0
6t9gK//HqFQGMubu0XnSk0XAV5ki5+9DLY+jgQHsd5gNeRms6BV5RfZ8hIcdGMaqzIa41lkyLpCF
bb7GdXino/dRuof9GBPzwAbWwapigIhSrLBebOBwh2ErqJYEb2Bjbx9IwLWdXILGER+UryuEthnN
0O74zHoP94tktGExaavjMCF0aoFYPlPHMIUHUf9qAXm+pmE5t2Xqjrwlc0FaRpSNsx3PZV4lV+sn
58WWWgr0+IYANbqTrKntiPyLtpRQbaHoLdzgT7Fqyi5vwjmaig7dFocOkP/zFlW841AUzfwdVw5I
EZ1h3Q+/y3LkZSTKx/05SKjxBNkj1bgcqyTbPpgTazEF4x+inATTtDS7r9NEWc3e8w31dB3pq7Cd
YjH9n1yEq7ZdogLu4Qt5CVC89LAYpyIQfuLk01WBRmrWnC42hblo2SXcLQ7Ac+CQUAkmk0149ihl
uv9nD/O67q6DoWbElmnUhB5uFRdtfYv6UgO/46sXgGqkQmbhJh4OlRkNDUpnHlppGNXdhV9O77oF
EvwNDAIkIvdXOoQoTp66j5MvAGu7hSu1VSGKf4baFdk8jptlI86XXMhLle7q5BA3tTnp10aNeHUZ
hzG6O5RJ5h8ehck5aWI50B5ucv/44UnRf8QHquliTEOkqefH5tUpV8qyMD61IurbU52qtPLsA7nW
DAj+HHlhtbDXCL0GfGHznCo8PMuSgRKGenCfN0p03Kx1APOExr/uMySfYVosWCG0zsH3QNGhNBsB
3wmseV6BfoPd0CzsCCnLDhB5avXb9oYn+DpM7kAfIZXVMjUA0fzIxoySgF0+EUl6V7/TG3bDKgPU
KSFPoHYzjvtV78L6b5q5v06fhGYTavy18pg5aikkDsjcUMu5dTCAGG5QXrhNArr/+l5HA+Lcozgo
CXUqEric1wOQzljKUhvSgvV48fIGEo9KKgePeiA7XKPS8Ke5eocuMy41XejGADCfmUEJIClsKJ63
0n0D0la+KJ7WpRKHPEF6vujbU80nsfC5JUozXtJJNoek38abnRj9msjOzITdjGAitVSrnO+U1iSq
tgtJ/FfaqdSXX2fjN/jkk0xio5T/EDyPuHCZ3roxfGUFki2+EHwmeILG+skYjBUtZGF8hEempPE5
2Frcv7NNUNeyBtqS6w9YFZtHe4bVmdlrHDNdkwQY2l+pzS25g5dB+9c9cHRRm78BGny/rR1j0Nnq
2uKXLkxPl0uswRppEFUvFk2EDMSx7cyLZ1JyXmEqk5x2E0tACjAnsidxa8d2DdHuWFRhwhrMYKAh
oJ/xTqJ2ZXHIp7uZ4xPM88uaBzeCmVffHi95NDBd5AwytKtYwmPYPnhlPkvrRYKO3/Muwt3c6LbB
b+NNtIYfpwkJTb3m18Q+xAzrCDmUTHM+biQlQQuv3JYNI2OwcfTAV4PXztTT/b0Kf8utggudIhMz
cbEgkqGFySdI0qBGd0rVFw4TUr2J2e/Zpan9m0UT1N8SfNXS8vYG+ouVcGryEnz/GoOvhn10RNal
AuWm5L1cJLwG4FhEOLfGyK1yRIw6mTyqO/n9C5JpE6s9iw8eHZKm8zlK9edvT091SQ77VNu/+hko
O0mkVWQOE98Nx7U/mmkItNBjlByRQfKXj21eXl6NUxLR6WhHhQuKHriIzP7/MQtnbty63sxtL5iL
VTo0I5/UrihAp3HQRYBQwuys2XvaQu81vZWjJmewPj+U83AIlTgpELDX0jDxbNVTQpufIQtBg/4r
+uWp40OcYiOxKE/fGZddU5lXQsofKGwO7mDI9PhrBMHP0p+LFseyxt+iuEJ+5/Oiq1JoCWB2CBK+
RYge46/OffqLtpRledt0fXx3OVTl2qc9RqInaL4+nINNU4ylPBy8wVhylC1kuXPsGgwVtoMjO/Lk
Aw6fud/L93Vf+8U55V5eY1u7Wgi2a5jh75j8ct0j8Ov4h0VLg3JzzdOAz+SItOakn2pHkLIH7C57
yumyn8+OpJipNDzUoKfswPh7qjhGCQk2iNRfRN+vgZ1gtCE6G3K7Hlr+AhFcuBAz+0OLreYUnaK1
CRr+YG/QIONZqlVzRo6ozha77nYQ/1WNGxZIg2nRjn7Mw0b3dhuXTC4TbBanRDi5Wq8NejCmKci6
gMzXSyT8OvJnYNwGaQbEYLGfi7ohAVCdrlpJTuvbI0fHNcBIl3oZWPpl1A4uNPh2/HaJxzf4Qevh
oiOY5MiN+qhGHuXioLubRI9b3dyl691QiayavILEf/utdGvUijbF9dz5DeQsipfg0V7lF76+NuGJ
cn60Kd+xLGeM3r4xgxKJqhWa7RnvvjaYHzgPB6aZp9coe7TJbvNPDtm5I9KhzUQp8TK0GPm/RWm0
s88WHi+gHhNLPdAElfWLrbyEBnWfVLOaNucG+tDJb/gFRCammbQvmR/X6deHgfZSxtEivO6GL0rw
EBtN97YTPeElr3MdCPN2rzSKHz6NYtnOigu9q2YWIm+hooV6kR6iyRUdAcHOod+ohkJSIsLvgveE
tuVpPCzSAaA21gy4OCw4zM2fZdRahc0NaQXRqYQyWKomeSO7MeyDOyyp1Tb0ZgGlS7Zu+riRUQQE
21cWuGy9OEpAUdHcphZzBlgm7BX0dHiiLEBFUkcq2mJ6KO5a83heM31p+I33mc9Bl93tD/TPMVPw
0Xt7wl/mFTHBdI0DlCgTtxc5O5Tx2NSU2q+V0OKoaNK+TO6q3Fphwu8qXXKnUL7GacxkzAbiocFy
ZXOTObi/FeBpIn8GFr+DSD9GmquV9k3ePb68L87+D1/wQ+7eiwsBEj2w2+aKcAzsqXiA7r+lrZIW
IKsnkYCZhGusvGAkAErmjU6o7PXmf+T1xXfdUsE5BeLepCtlsE+KRFu1H9LPtsyMv8B2CfxqXkAA
PgMOK/C+XT7YRXwyIXsG3db0y1KNqqcQ6od96pPmT6OoQ476E7Hif3fGbhJnlh5AjxhYE/PU031e
vGtCp9GM2muSqmMsF4iXwkKZHT947b99qUldfnEvHvhgQr92U72aFP8fktN2SeKVEgREk97eiP+G
5inpZWZdItMrUFNsEQfdzFuPgmUHNoyfSBuMLramXFtIfUne3djm0rRF9j+ltu8X0tjHcB57pvHE
qODVzDYAAjcPhzQGaH62w8athtQ7v4WqKpWW//h4StTw1YLNna1oWkWkvV4Bz6Sh4FzpNjFNn4jF
mfODA67h8FB7u3L/oGpirnUxmHMRjwW0PJ3lOS/vzXOb8DRUiNVBz6Ez5cFPLi1eFDQiroYuEsZk
lLAjCqF/WY+lDFHZFdcZWA363g9P1OQpfVXnZVGy/ZQ/kLBz5+svEl0nH4DpfpkAJ4nukoi3ckE0
Jm0kt9+Wo7CPaLgURrXjRWDV+sooV1PtfKNh6b/0XOBtug4r2bIk5ZTuH54w6XDdv5XwnamzNj77
Z0ciWHUK2jJocUf0qFjvMz7psqcmndJke0rnvmrKsg8Rd5q8jF5TpWsPgBxj7YlA+Ck6tyvAlfom
mHechPFp9nQt6uXg/WJ/uZANGEtnc0lkzr8FfWKCMkdhn7loxIC9rrTno9aJYYufvQLXpG0ZmD+C
A8Z49SGrIhw5sBNR8fcEJy00ECyhezZaWsgrLKmF+E6t29zMYO/ejDtZJrNbTlNyTkP1Ou6weM/5
2zAnmeWfIkzTfV6KsGZrV4wJEjXeKYfxB1rKr9keSpyPenmWVxyR5hN49lOndYFRkdx8A4ZIQA2U
7yik9w5/Eoh+3GZxRyn+x8aLDDKuLzjUg2iDGAaqQ9Gs8cu5mzp933wXYmM0SfHl3/IOchaPHWaf
iTS6sW5+N7v/zZMu1Fhol+2hfVou5i6nLpc0S8INGY7jbs41NaGHBxm7mblzLwJH+5aYG5OKgGrH
qiKBxrZINvMb8VyryJmohRl8Bs4BnrEaW9+yT8lm1EsJOLBn/+5n/8povIun+MakDN4cljTO0b1c
xmpKZfzU+bHecK8TXuNzFiZRQL2v18nlwklQHor0IW+sKPcCojI2ma97Y7Pz21bHDcuBnL7xmafX
kppSIhO+B9DvcYcpzwnqr7SWOeXpKiJHb/mF5unWiQrqO/ybxI1n040rLqKtPTMfBBtgmnmHlEog
Doz6fpPPcag5BhX9F5aze34TEbkytc/GUL1GwrgG55vLsECaK2RMbLW51i6GXmOcn2LhnWPapak1
gsyWoF+jgd2EYVolfFQv9NFjLHzoIXlkhETcvFJcjPjI4FX8o3f9NyZziWxnO0gW+oCrjmQNg382
A5Ybk5v8fhsetx330xMUi4dTYTwEzqDBVSCR2VrL1Ww94LR5eFtiWYlw3jtMNkTEBA3MaAEtN4ve
ygxkUKXkFXHY4P51zMB/Fda6/EYJD0Wzh/ArEOEsKzJNcsynSff4MRidmBjp6CDE7GXtBAiMeSKM
m7qNAdpBalx8YBj/iZiEBCTqhRiLMdKB3PoOiSeCCMoRgCUNQZHlPZ3CtgJzkgh8ss0yiKDzQbYU
VFWhzjstrCr/yD3gAMjfpg9hWkPdB1TJ6J7hBG4dc9+C75HOdX5fyXyMMAF3BHzr9EZQ1YVYiAla
semC4OssHZTpQGlQs1a9j9Nk1wGBcowJ1D72uvkFnAnr4zvINoGLUEo2NODT9gIZnX5pKgVVAZ2E
28LAVG+ADEeIkCgMzUgt1xJES+fWkNOWO957jQF8KiFf6iNsIGoACcmmp0dBF0uFxWNXvs3DlLP7
NaRPZQmAP8SMBT/eCPBmBhDw0S4NcrykB+JheFTHqY6zRPq0GlYrWQaLPAvf7GobiL+XTyN7gnq4
uDJ2B3G9+jriwCvpFrGEnOn8EeFvZBO3mbuxiAKSLsaZb4yxn2qTyYe7QyoQDdJwFURehcnktbE2
GMjcLI/iAalG5Kc9EdxOIoMRhcUTnf3nMCOCW/V/hkN2fjFWZ3wIvILhwjh1EE4+SpQmFrDqi7vD
ob/AFyxGiT9++wO2nSqeqSZw1Xy7w9sSYKub9LpGRKgM5mntNjWsmOcoZhn8vRtLVS3UUUuuGfa9
SIO6Bstr0KD+I3m610ROBMur3GHyMRJPvlkhOJzd1U1QVKVXuqb5Kwqad3Shj2WdA+5sICvw6vpC
Eb+DWN4onwXC7/5CoAoo7T374s28rboVLy2NugIFYNAar3NElRo4D8u6Q8k8LAOsi4r8g4hf9/eB
DQFhQDSoBqVxPQhSuyYTPLVxPmU4iOhvbt/etvpQd3gwi/0hZ1S5DifShhFRF+3Ax4vvhhcqkv98
y9HawQX22go/qsqjsush1WrL8Wuar8qQbW/8SQ4Y6+W/y2/SyWwm/1IBKAZmyTKnjVlk0KGRWZve
UEQm1Z2gPLz4QGnb+wB89okMl5cjTxY/NGq2ksAEUoCYKPZdjHlc9F1W0EnhvCp2cXS7VgokQ0Dl
OLOi7mzZZhXerILK5urRb6XcfY3Uj0uNwcYRv8kbxZU1VRtlR5RZ1no+dB3/QuQbkogpf8TvNSG1
rhL5sOiTMMnTLQ+jlb/ZSOPpdsEBE9Ie7O060uAHoqt07A7H0IFiFwrW4zYrhI6hlJP2wQ2L+7F7
5xOpKsQ8HyC2SODfm4NXxAWYh6ZSXhaG4ofFKuRwmmWZrAYHhMRld3Tzs7jbCwE2AFE+0fqaArJh
jJGDDbUcMBHlXZQn4GazGZGGE3I2uO4qhlL//kT/z63HVt1seaCykrYFQgsblPnvWI48K8RYTiEW
8u7qpZh5RQ6OeQOf/0faYt4Z56l5ZEl+3TVX9Ou3n00V0iMErjvjQcfxEGTye8nh35Ad2fS3nvjT
KsQRO7fxAFlTv48MRSu9GdXFLzO4JQjiYiVINWCcI6OGcsvKS7wMoyWAH+I9dFLD/M0PdMUJnTJm
tPTKodbz1WhaPtJgiidx1+jrxusUa5L/q3yD0WEnzu0NOYs99pktbBSRd9IUoZBDzaJXRR7fYVnd
+guLOjZEgq4HTw79ve+e/JeKKBXX0hoqa44mexwS4d1r068quRZ63foTbU3i91Jeo1MM5FjNFsPs
bHreqXUVLVpybgOQYWf2FXm4sU2ob//NKwE6QFvraVlEsVfJ1IM32/fzlu6GBOvkypc0m7inEkWy
HLGooapBTY1Mx1n93T8Y5Rd5z4BfWcHDZzEn1En2d4sWITSSbvKsFCAMpLGwCahZJ2DcS6mQtN2C
DTvw+qmWVXS1tM6JkG9BKLSGI6FQOTYXSG27+ICkDVEBU0Py/BL7i3bIg7mT+ragoRkSu0VmNGVn
e/zbKluspqYoTgYIEr+A8DznOzQ0IEH8SS/zXYvdlpJN0WAl5KSBHY6w+kRD2F23Kw0vzNvJB5yW
RU6DRgYn3Xb7uWlS2q0Miis9ccYK52/oalPas9/0qX6twSlmdUtG67w0OM3jpR32djAeiwHudhu5
JtADI0cmL7LcnkT0wKzcd0j1Hp6KyI28O8Mn/Pgx4c6Z8a4prXDSna/CtHuBvD0l84AbiwndqyQe
h4HVkQ9c1d3gr7190/+9f4oXUVrpwD2wWUL1RygQsRRmLiUYmlCEhXMh+04bk9npEUJxi82lXI5+
69JYHicLXI+kp0iZEhZ8CNL3KO6zrbIC6uLg2j3AgYTfPPTpx0MIQZXgSAAxIpY10ksTblo5iHGF
qyv1ghVXfMy7NXQ8DvpoiTw569vrNSOagy1itUxPAXLp1ptmGT7E9DFyKWrVzrT3SNrqFo6io85X
ky02pyz1TtYsEumtVT9BN8dMleaktTWnq5Iosl+c9tZYYoQ+KLD9nRfxUpLMsv0AxlipbvpC2SUs
pOjQDV1uluV/NLLZ5jDSbL3EryaXm3dCDRO5B0ouzhQmgN5L1jIUiH5bIupKppqsLsXwadne4iTY
cJKhfGG1mYq4/Q8I4VbgoKIXf/7byrmNi8GrCatYdVK2tTmOmo1uGikyBdGDUYxuYlPd3sKE6mjh
M/0YbcWa5JRAcbdDwVce7BSfeQ7GFtWM6bxG8EdQrk6juL8w7v1qyH2vkMbwomvE1308RblCkt2L
YTgvn39Jjuj2WBoqZaKvh4T5osA8/bZZQQK2PRw4B1+3rcJlt/xSqaYeUZyDQopVwyxPfVNZUfDI
89qypheUQxMbKXHbCcSPCSWs/r48tsqzceLgFG18ou96iGY9TXC9RWq6PB20Thuh4xfb9brxcfJI
mnI6ybbDKBMGDQYDmSEcwZT/jNaF61hrM68Vrbnp0KuUc85eX8qKjVFT4Um32GItNothxRo0RgQi
0EaUspc3AtEvfMYH9ONH25FdW7S6XNedaAHjZZdQ7+Q2bGJt4xgmBlXDotoOXc0lSZU9p+n4yweK
iQKCgIX78OqqEYmJ/1nKtwnUp5IULzoOcp12jsIk5aNMk36arVOsNrTjsXsenyhLhM30sSYFX9ex
psvL9p6a2IXFxPyGhXlgh9jbYQMUR2W9K3tZpJDxOR7wnjwxPAFRajA+7tlGx1mMqLSXGk4ICa5O
dKwT09eRQgYiEOIy7o+kilTKba91Hh10h+FfdYed7WNP7q3QpRLCLjU7X12MSa/Q7ExrL2n5XrzR
iOatDzZo64w4uYpcwDcH9l7KqIz8x5mf5XIHM7xolqWEdkOkQ8zt4v0rMmbKgXXf4SXxLNx78ypI
AEPdLSp+uRntMBvHUyl8bWAgitR6CMacv3whJd1nsaNyl1wgLiN8b4Vu9Ev/Ji2o+VLlvkEDXvym
auOZjgtAxciBoe7h7OEqjcEb7QZOmkJgHelQfiO+glhSv0uaZe4UH7Er925arHEXNSzD15KBcO6F
iBzV5UJWue2TquR/xm/YTWRON/5rW6oJWho1jrW7XWqDy+vYFxWjnDMcc+v3zDx0EvUpOjKYj8vP
lYXZN55sdbyqZKoA1jHtnEYkbUYwX9VE6oiuUNLGNuZV7ltwCJW+BiORYO+C4pq69W0f7O5hDkuv
Nrw4ekS3ljxVYJoMSxGzQLKNYGMSO7V35HvVrsS6mEV1dOfJp5owG1DSCU+fW/A+RIv6/BApbhha
SRc3aBHT8ogEZJ26w6b0wRTutCMGk90J59fGoXvhhNrpLsJ9+1N9d9STOV9axsL1b9B3TS5zk759
cSntfWe+VXD79+Q2qhJzktmoys8UU4ugJyDSC6lGds2AacBSvE4ch2zeIapo8kyWhvJxpue8unGi
6ta+CE3gqMByHNjhCu4YE03xQFQ2H2XdtYwd4B/KtcOpSBRjU88Y+45hNFSrQrke3zJtCVE4fChO
p/9dz28wVzq/zKQjctw4g3Xs27nLu1tGsMVt2oo1kVXjpeD8TgqbH1CBsVK139fFOYpMOJYdJG4I
vtIA8yZAbdzxJxVDAN8fBGNupiX2oQHIkh1onzSPILnNHXRZYia0Qa6a8yBWyziJZzwFo+nC2Mrl
UkWxezVsJeXcWjTMBhiCpEoadSzXUwVr9OkOCzi57KCr6AWWe/6SBGInWgkhHxh7RjMZZfnPN3Xs
Lu5fCWWskW2FP8YZhP3eI+CZsZxD2ZJIeYslgAlKYnCrLyT4q0Vy5GQIS+JGytsMCFq9Ys0H+wXG
Bn8D8FGd2M8cYjLn/pXUNPXMV8+m8nX71rLbQ5SCuk38c8zYRssc1dDx/ihMgjsFp6o+VMKbwGoz
+3HzvgGYlYAFDB6cOhwT7GUz8rAQRKAvg1tbjSQRhu/s7uc8khcQMMfaNk0bw8Ya04wkSLslENYn
kzCkCYSFQjkuTKgoNjLLMt4zyTD+Mg4FKhtaSpIPeMvrSPO6Nh6aItHlD2iY3reKnzPLg9MJttZd
+rPOTxAN3I/h1lhFlLnTQEXQNuQx+vsYE+IZZy2vmsUMZtV8SOUpQxtwDdtQMPmyGDnZbcft9lk4
muwKLJYk35OEVsnVVQ9aDfyY3Btos9xC3kbQxmkIo11vrfNBsboIo0s8a2ap8L7wRnEQsdQJcuhv
vZ7+NxwslAEDrHNqDU3193mcviyDIIKgsABNZ0DxjtW8P+A61xu7ery8mDGgCc8W2uCgmZYJcNin
k0hjZ9Xp4OwGBuMx3RVbuhvjSbgMbtf2wJSk3R8o0Q07oHUKfSK73dR2Q6TZk/GXtCBdMlsfsDab
pNo/T36lyb1KJTdnvB7637IGyYLxVw5SxfIWGAuwFyu64hhHWl51O6nq6Miq+TI7nGkk4k2JN4qb
CyDKfvIVYbcfxFuA+WH/BEEwwmjpRuXMAOKxAfddS8gSFpugiTS/01hGiXmNVazIBbvEJQSo1HsB
RdVvPrYqMwFuKr9qfP3DlafGhzVbU5i4NWdgD6uVV/N8kbxA3mMquESuNIsNXFUaTAzgPvoO+XIf
Ir9UngiL6Ex1SJRzd9xlrOPUYVwM3sSZod3csI5Yf5VDIGZ61NDo+2QIsuP98yc0wWnUV7nTm8bN
4G6v0X1NmOn5M8x33jAm91gFb2XjBlXWYOjZVED1zTJUOElm95WIEsgsB9ix219l/RLeniJgGZoe
kbkkpdqGXvoofx3eVAsKDnQBkNK8BKNjLRyu92cQYo3i1v3hG596R4/I5mABnjbN+eG86zpP6+3H
fpYYPzyjfPxfi/Yj4Clzx+CK2n9quiYVfcRcpl6hmezvojm0CtMgvuLfQT43t1c3qRjp6CDKxKJY
qR0QFANKCZC76K3DIpaGKi7fJed+E39AoL3vc3cBW+mVNM61jlPYBi+NEvn86SYia6eg1cfsXkHX
QtTpj43Roqqzhwk2rHu58ygzyO61HXOhM5e3Bzi6Vp1pmVnAamVO4JV6aIN+wfTR0TDO8LU1SUiA
dk5yW5pJaW/g+0B8/fBlG95k06WwV8H5dSBJ0Tm9k0jPwgGIIPAY33tPSbdxLWILQlmFL+empK3m
N05lJvg6YXDT6kgMIwoCDFl9wNFMfbkd1mZ88/P/RgR5oY+TaL3pZlwm4BBDd+FnLOGnd/6Tzd6n
oxQFk12DDrhvAkql/PtguCVRnhvmLSZKvTDrNK0loixnl3mrb2ilUlo3TRgmGaDdcqpcfCetKHdw
JFhEfwz7H8BqKOEcg6JcUFxe1DAxUMbXksxJxPH04+UvNOvSP3RXDXoVrFmGbTHgjrS721VtFc+g
lNOn1ZEzS06NIBgEABEJOPck8YePlouUn9UQXx6Ercu2W2n6PAK59YiF5lUm/EYcutumbU0gSi2+
s6JsrEEHxRJR+if7QirlxLnONfnornzBoIx2yWHJxr0NuG85//bwfx/4ZtGGIswyI9CPtvBu7t6E
FeecfKMwmCxWQ3N1qDzF3SPtYUB9nWYI07K/1+lFYXkLscOt+OPjcNs638E+r0lCxpgo2lEQZh3g
QWj5zudx5C2pqJ80q4NC5PRdK1zI0Fzd9ftzJKzKDfZjtKr2XO6F1WTuqhHE+y2iZZTbFKAVnLvJ
K8yCbajtpsfqjrrafgRuE61m9JU/Z8AM4M4cGqVIuAaHuHbjK5NBkNRBFqpcG/EielW302T7cFkH
u4X9lJ8bxun0vIwpH8V39nh5drYKI3ylwwFLvCIT+ws3hcPqMaRxjwj+hRPPlndwyd/djfZYU33o
g7i+gYvWMeGRnevt4sSQrc3Sx0qde6J1agOGqxnAWJGd5lO93VIUoYFBvpsDnaj6HklrXmY+KfwW
pHufviExuMwdMcQLBZwzLTFFn5EIM0CdF/e+3paotU+QYVt10pgFTTWsH8lxgZjeprI+8D28HJIC
8W/+68fpLN85O/9t8CVkpAredPer1m5BkyBsmR3fIiV6/FJfhLvqr2ihZLPAqfLBOYaTPsnBvdpV
92XzhgP02gT9wJNIkxRHobqvjVaem0+uTZBdySTi96nCJ1iQyzvyIQQ2OxaDzDMww2qZKib7p7r+
exF2H8z+cz5ISri0lfNyOlD4YgB8bswIbzp9zKN8zFuSU7+wbFeBSMawfB0HSMzOdRL+FTMFxWjw
UIPs3QaH1OOzqH6d3XibcOqNSmLgaRbojx+fQYHF+iPF45K6ZaruCoJCTig9/T5KDXjO5seLUrbk
qsyqbAtqDSs7gMZg5ypgTO7+lvayhXEMmcw4765nvatCAv8FHwXsb/Dm/NGIkljN9cxVz2tI+JS5
DLgh69z6Ov346ZlE7Q+E/WYU1C6tBkVmOHl2ktZvF834Ib9FjbwnjYs9H1D6I1o67axzNNxTjN8X
jVtJ70E9oSXMC3O57rWUZISb2uvnaHNUPKxHehltCpEYIvMPg1ZrPRJzYTk/qVdhhf3PEYAUOYO2
6g6GLLFu6H1jVP+R9pnE8vEZydyJ30f1/CPWNfZcLlhr33o40vD0XOdHNUoYl4+T3sZA1n9V0gzW
nJDG2DpB7XHg7ALnP61TGLEmItgNjrUlU3U5UnAA28bOa9/AS4Ul1pY3SkyVdQUwTmH1TC920j79
zGCHu53EYrT56prr+o8i55jr+RomdfA69IdBUv0+ht/raNIu6xQJ27sYlgx6OHnhgQ+HERv/XW73
Wr8sZ2eyA1yrOaQyJMsj4S8bkcZMANP/1cMENQt11F11ebmxoYYU6E+J/84vN0dT2qNR99qCU2Dv
IOmKL8jvbOy2QVoy4BVKUI/9VWkYLksyQU6AYnDthhOX/8pi6kRvgTHHJgVwHZNtPqJeOMasE/zF
ZweK3j7xTkaLyWjlcF/uEWuBZfozuDoobeXV+CAjfmgzVLctWLl/UrlMQrYWr3b/FS6Op8zKVLdL
Rj6co76B0WOFUr71MFQ/ve4EBiX0gHp/2cawfvE6nz9ztYoeyTow9Uh6qEGK2/ayrx0BTGvxXncA
nNGEVM+mvX0Y1t2XV37wZIZj6adAVLIo7eic3ArlLRNsbkL9EcdPIHQ7ak4NXmzKQo0LTUzsbha5
PvRMB4LnPlkLrBmkscfGC7K39Yaz3zaVmbUVTqjZUFkZN1KxIw6GsROU9sWo0qdN/9GznxrRinIO
b+kD+FJj1kkdBQyXocWjaC4ctACnG536vcO0a6qG+GCjM0VvFV0W0ct5LPjUDncUNSWG8En3+HMi
hu0tbyYqrj2lDQvwwx6Ewepzynd9AklEx79k3REzlBcjduM1zMEun5svpC71Gb7j3LjFBSiMZjAu
Gd9TBzILDPyVp+HXM77daZc+LOHDFszMykuhHdakJLGRMXieyfJuIhNxZIHzSl6+QxRHUbqqOdjC
AXyXfm6pj25PZKxOH3rghvp/WieussJRQfVLt7JGzbQAYFMCqdeHQ3P5vNpYHyq2XPMTlUNCOlfy
3Gi7O4T0jDv2wEoxixkXIAYHOY0OpZZbHdQgu5nnBQrHyjJ33gTdaPqTCxJ1AHhwT/WWxGd7QlEV
o9sSfX32d3QQgwPUjMrrSs614HrTGJ45e2Vh0HH1tefd28EbgW60w8hUe1ZaDDKPtlc10fBdywi0
O22N9c5W3f5M7BPZdYLB1tEFhUIAE1d2Kp3G95YCU1eudxynZszWLHDsWhbJaXAZaxA9Vy+tQfy2
+l03MuWYBMZafqArwsXQhBBYKspF5y2rERa565i/wWeQ1ZuxGC7yAO6Y212ONlozqp1e2bkrljTW
ccN3E/XSSMHL/bR5o25Rg+PtDbUvwxe8OdgBAye0vS3DUh/g9AfJif4C/ivEJwlWWCd/t0LrfhKU
bc5rjAqPh+sJt3pLrbQm0FdV055rgRlHAeO9aGWKH1wti3Xg1Ps1Hn8Yt0jR07TT4ZNFH0c2g5/q
905RrIuZaF6jJ3kXaDRpqSfNHw+Heu6u0DDPWltJWDM/6XgfYWc6OAzQpQ7kZJNtsKM9+1Mwo8/X
/3RTCpMgKREFyaeKBBwkCWv2t9Z5mvecRLS6F7oDArRSIu+iNoQm3OuoKFJGdsXb/6JTiqwNhwKX
TdXFuhSzS/G7eeso8Lrje7eOUL1jKiYy4ZaufWLNjrlXaxqi9y60mAIoTrNEqop2IJ97uBJ/H2xQ
b52AeAq1x2naVq01LGB72QazvsyfxoZa+Z+6c7r5dpS9KMLNI1L2sY3C8zIhjlYmeZougsN/dXni
bQg77aUTvXKbCVpROoSHr2KW3vfjb3scCNP6OYkUUOuqNYm+TQlzcRtBFzuw8ss7Wl+EfMVzSE0G
FM4AWJ5m7vtZ6PrWup+2KZn+5n2kpP9NdTbbYdaVbmRre9QbVgF9bFUHzRvTBqcWOdUI2RsRwSLa
Bq73C012VJ4eRRlxV25i8t4ufHCpIKw/cXdMFMkM13/YjMKT35lrMUXhBiK3lloz66x8TSImKi7M
QG6wuOEYJe5JCooMxtqSMHF65NJhYoylbbjXGeGHpRJqtPcrKqwPIoSMS0JYBkP9uxg9cnD6svqo
H3bNrIs6kYaJPtkTh8fWRr4oo7kR5Ao1ZDP0B6yuR92K5KSE665ildwCI5osje8zOBITkAYmLdGW
rkytHAtg1s9w0XkurFWOw3o5g337NiNTX1SnqRvcfIPHtdU7PqFVd24emaOj/UrbuseGE/O+D4gg
ptRKMpxEYY8Z58QT5ScCgb9+r4ZB/AsdOfL2TR+2OOFiZSCZTT2ddvhosji5SCRBQPsWzpBGDgVH
N78rrmkjWJewvFrSldVhG7wukbas49k8dITzze794P4cNOoIAgW36YkIPNQ3lLa6fNRbNPcdFZ7h
bHEDPoq0R30DAUXngpqiY0O7s//sF/QWD9yKJmMA6mTbHPT1mXJnO+JA08DDDozH+hZeo8WJH8DT
YEMXrX/j582TfB7r1bcDCP1QZOnGcUAkXP1JdVCZ7hMOTdIE18jSsM1iZ+aRMgQ7s2Pzv4IB3kCb
KQnR/GerHKsjJliCREMg6OnOLB9obMoXzOmUuh1eCs9ek6PI+V43/kPxh23H5INGjWsTU0MQiVhs
dHKxXj+7YSLwFWguoBzHMyReqmoqIP3FcDW3Ztqf9QwLz6NiK5LjDF+E2kTr4cY8vA4bymwyEd2q
zd9KsfZmAAl/ycLYvmK/DrvDa2GscM8Ny1AS8P1c1+8gt+27Yyqg9vHvLn54UPZJrjshmie4JKid
mownUQeEt7NX2kMJOUhLGfYhlCF3QeJzqnxTQFnKIUwbBNMyJ8jKBZEeiBcvGHpbO5uUJjgX3r5o
5/aPzCCX2I17MGWWmVMpno+To7rJ3IcaW88whuceOVCM4tPYC2rZVwrZjDgQFdmtQVBk+bdHbTRC
yWz6mULG8ei1HaN0M4FdIa2bwFkqMgRM2J/z1w9UuS89hpTwUA/YIEycJswhtm0hl3S7529my+1O
XVphh1Py5gUQKVf6PVrCFwOpJ5eru2rL8CUd913n2O+ZUSvWWbTDmMcNf3yQwgLJ7Jebz6kk7h3H
PvpJCEgjg58jX3HTz+NbUeg+qDR8d1asNmpYGob9l+kTeHW4RFpPcBnwZ5xG7o5kf05+CT/qb28O
YhInqY/ISTYysc4Vyz58gmGTXcSTTphwl3D+js1M5Tc/ey35GFGkvzNgOS5CIBH4fgfs0ErHgEtF
tzdX1/swMVfdst5XOqJimZesASK4eIWhspWOX6CO5eHtO77VG0eFdhPlvVQdQOR6q5Xif8nO6AbY
iWZUVQmBppfL+xp6Sxddf8nTFE5cT5jZ1Rq0FFK0ptmuO/doL6vPB29CkuEtCjvgphzrXuxSHTu2
hxytrqFhh0cdeiML0Ok94xPmaOlHGh0h/mSy7CR1P2aPzq4Egv+gwJ6JBEQoljoBQ+nlq+rEL6ud
q/mGWuDjcqyw7Cdl3CWFN0VMEnUUHm3FOYq35kQU+xhvwmkhNVswmQY9v4rD8ePDTTk0Y1ytyUaR
4ca1Z6//X5CUSS4YG9Au8Lb+oMHO9hBJq0Jr50K1I18Yp66JOCeBPCKgMz0klh2X+lTetq5jzvaD
Ab8f0eBOSze5nyU5kBtP6PkVWgC4VGzx3iji/ZRQ/d1ju4TbkXbBBpdsdDlt3UFpqF4J5gbW4UsU
u/J1GpU0M683C56Ukl+xqY1TZ3+72tkGM0/EAAWf1Oqxxv9Ai7pWTIsmFVrWD5YY/p7UFQ4lCRns
u3OAKwLxTZBoHN8fFnnKBYsgyiKyrSbCFoIbNxBP1Ghv1fbcbwhKqe9NJQ1R5LrPRKB1bADPiD8L
OkdlT2jeXVnyWleKBiG66ZBuQrx//MOexVaUZrsXen8rXgy5w1MWFH56PyvvWfDrestFN9KJp0xF
YqxsaJr12myF/L+7O2/vtE5SSKbw+hK+60cCqqSCE8WwD+rTRrQZ1jiGWnsfX9Ilp+zMQJHVXynC
2Eax8S0nwb12ac5wLcKUf7fyUQSxxv2mYQLtWekFs27rktbQMB97IxzjQJHbdrt3On+faD7C8tfZ
MtAj4Fl9ADP2ioybES8fUfYaQYBiyn11DHx8lZ8JIPdQ99UdX4JiSNzM2yWLj+Wt+zA/JBtB2PEM
NB0uP/bzKA0r2RryXgtH3+EZIgI0OhhqxCcwdp/ZKAoTGhEJUenE+teyZTbEdm7g6MPr7NVceG68
MJ5zmlsK3LMrWE8EY2HUqKf7X9RQVY0iaEw7fjfZmgmYcpr40lubNvaDF7Y7Y+8SpzFvNUii+SRK
SmmzrWTWfBFlv9b6/bYKYE+jwl5EuqvjaCN4LrYt71iOQ64egC/wm8p00IWtxuY8PRzW35uTGe/q
NNTwlUroZhd34T3TjGonB4V2gAVntvJdxkm8m1s7mLF+7NbEsqFGvHCXv0QyJEWseJi8BrvXkp96
hjyQJdowwZ7yvQYd72SDNmc8Jo71ghfXS7NDLGogt4Z0JyshSavzp5trM6UfesY1Sbyx9Q2jtJ3w
nD+/JilVRbSnsE9+IgJiZuYiuJq3aBFlqYYVFCFK0hixIOfUYkRyK2g7+RZPy+GwFcqKkF4j9S1Z
UpvvQbQciqLgq6bXO04yI0pLL0V30qvf1Aq/Q2ZRhS0qCSRvQu2BPLmOBjortuc2UekTv14yRS7D
QPrVAcdGaNZCAQW6dldXapqb1Jx/A7/ub/Y0P39NEwPbRaUN5Oqic+QIjeFeRfEu+bFAPbncKv9o
LS2V+IyYty7sR2r6uXJxkitI7/Zpe4boN9n7wJnOQ8EMRuY06qJfiFgCI/EnhHY/NT7S+k8JCYuJ
2/qRCsUsI05Ydednf09mZSaPRCcEZeaMfYoKp6UTOnQ+OzDWoaWoIqu3hUv4jEMZNVf7Q31uARQh
PB60nwP2fnp/bJKqtE5y+4m3gBwawV2pPqcQPGAJ1pV8utrXS4boRVXR6qep4kdZs2oVzEzOlAHL
bokFjkZjxzX7GiKBHuI1WKvQMatrhtdAJM3J1sUEhK7SVN5UCYrbAK359LlKugXWyUAhGPPdenmD
k8fU33Huhj3t5QysblUbmElt+7SKthAmb2aB9s2IaoP6WgNrOkBZQzgjL28JvFez/oczjglpYssf
FjCto9MUJekaA7jA4V6q7aFaFUTq+zOWr36IK5I1SUT6ywVtVT6uoc3YAu/gQ5V2Ew5GNhVQaIDZ
asAACJjvEw309qbUYsflB9edTHS9NZeYPS6cx1ChCz+EdVtweZg+H1qeBh5+hCzkUk80aAr+0Bhn
fZGJ2i87rHiePBkMBwiSdK4F1LQSqHs8ZdyWY3BjUoeg8pubCsSUz+yeiUh3qWBZjsMQuXKxImjC
6xJ4gBWlyDeS98n6w7rcFecbzPWz0CA/iSjaLRWBTIL1oDu405kMpAbcFVqxHSTHM2mADiFx46S/
mgxtxd6YgKwKJ0XDn81UxvbQJfsmW81wOLeXiFsMtRL1sBqQQzsF4m7wRmGS4CAVmxW+QQgLAnYW
9zdOBfQcUkkGqWWLBBGFfGnujIPgwZnWk1uvAYOKDzrzvwiO9/xnbAJyhN3mmxYNbtdiSrMsC5D8
O163PmjyXdFs5fkBmH7LS57zH/T4DIVQ/xNcydJnGLF6lOOaPsPfXitsBINuBFMF0GwcctR6bvsG
udYyWGc9Ug33jq8Sj0LK7O3bDbub+28W6DqYlmiPke0IMNn6gQMfbxHgJPyz/4TXFFQBi1C22Oth
ZPux18/DhV9bQH84TUR/AkP3Eqg1yqF036J4W8n85XMBX+to27KrC7AKsCLF1CpG/rzNhbC26SAw
GGVMP8x10zrJZfPj9UcT/N42WuuQxmoV4KhN7D9EUQ/2sMeLlEORxT22EXDFtPKupZ49pTPggFxd
5u2WrU+R9pNfE5kTOtPpAaP9sd65J4zdT1pC7+0qOSqK32X0/o0DkNEMphjvlvQGoI++lSSoWOic
lueBo36kgSLd8+K0SOqqjKtFqCSCMAP4l8UP/oA4MtdLj+HbEWBG5oqWVQibj0iu2Ug8UT+52h2+
zO28quumH9exIhn2ymks+dxRdg2WB7YqYYQbyPD2X0/NK9yvP3flDUavla7AAMAYzT4XNGzBfEeQ
Y/TSCRh1FDTn6Pw+Af7BwJ4KhNqq2sEZrb0r6V+Tl7j/oCGmNTFNiLUmM4sJomW1Wm3yYiXAkkxz
01n3tsnEOqXaoxD11zR+ANzwzoEqqztY3Yne0b60qtaWsGfeP54j42+jfsaK7p7/sYztzWLEw/T3
M+Mj/0V15b2z/1R/dSh57uVk4fiCrjNYrsra682peAQlSQfKbANxEkP2nBcDXHIJ/x2FvDPalkxq
K6QdEhTFl844gmYj48LtRlyCHDs5i+oo0+eh/hKmnDE3BTWgdKN1SBBBkpiX7tI5imqqt+MomxuU
tF67qMK/mj9GYA5T8hCtEmbdNBWCDPGI/DvC8wnqqyk3gvGj1WKAQ0MQS/eHEpnsjIg+shWl9v+g
/vst/n/LLFczqpeihmRNEg8fmPPrSR/LOl8w2bQrhZv0Y33WHDMk9p/rsF86sG4rIvHgZgUnLaL5
5SxCzhDHe1XoCy/ZHmKwVWGv7T6gdG/pVvynzc7Ob9PM9KIXa25BFAnTuElF8M1pllb0wkB5XmEu
aQ6L+rWKRjHa9z6TX9+MvqaO4sMz5AHr/MpCLQX63hWpRZ9kDkq+2ZHOP1U6Y8U2nmbRUbFP7prH
h/XOqZGgYUUjtjgK8PNZ3K284tfAFzNwgIsAZgfd/uqKlm1b3VQUAcuyCbyTgR2YCVe0/U6ZELrV
2N2f+IEVFtcireC6yIdxTvI3wnAbZNj+/Xg8qQ9U7SsWeMjbKi70q7i2FEEmPO3wAjbKYjb5WNte
fF7iHMk83DVAuXwcC3BL15u5unBg0vx/qqc86rCWjl8Eev+lBIedXTF+tfrWDzObI6+bAAbm2utf
3FxSQFiditEAeqcKGvebnfJ/jNulKJHn+iLBEMjNA7Xg3VkC50nHl51/TV+T61c7rucoTO2jnH71
KBaOponGaYECh5srQ99/e7YRs9vFl7uXnN1lbFGlwfceyYXDdKOb0AwKbDIKyezZH4TBTp6N5zKt
YW1LwVaLha+UMuxl0EKJN0XOrzbVsN5W+JzfrEkMhRjhMoQybbNBPq7cr+R6WDuJuksa7hvNiiJi
k4p70YXhjfhtbjkuo0vMF7KuVrGSb8OGxYHbzhowiqm9JLHFmiQsO8wmS4sN60cMRUwLT+wX6KsX
R+VcQb8qg5dqbn5RRJZuiBsUCnyeGxkiGWzBPHPsabxrD9AlnksFB/8/ZnJ6zsPRbsLP31Hk5uwI
KCX+rINiyqO6sRoneahTmaQ+VGARQ0vkubWIo9tJcPxPQ5rfr2iDIRcUbL4KTdhIZ14O9mRBvozq
PKiTteA3g8jmq4GEFaAleryzc5Ca/CzinLt2CvcbG/KqtSN//uJimSafGpi3v1zsxh+u4kqzXoPo
ARJ1Tta/ZLByBUNGjRCj15EO6yW4hfu96KOp+VJVFYjOwfoikt6DkfS5Tj2EEq3Y3+AbAnD8OLeV
yPK23kKx2KwNWj2PZo9MssqONdvdhZx5v78Z2fp0PbZEX+b+43L043NCkQedGv3gxiehGM50Cq3/
wQh1u1ZOetaU2bjlBqK8Ez8XUImcXCNXNKz0GJu4zLZmmZUcOSHWEdt4qNf9MpClB58XI0rRrFLS
ijHs/gDrF0LeQPlIxaZW5E/jbBAVYSskSOwyMymn1yiXyv88nIy+w/jX3jTMOg6v7NOPY3gOVyFb
nzDDDWrUd4Yu08izjSkMgcEYCCeSzhkooBrC9q6R7HHhOgJCQ5wgNcj5utf+LMiUFnPnPACJnZil
L/lRhGsgaDbR7qOmAxIo0KFeHPaILJOwli2kTaMnN+ePvSEg1NVafDsAI5x+zGkvM5f40uP15U4J
WqBw7on9KyC9T4J9Mu8cqXCWxOnrzasYBND8ul4ZJhfvOMwprEJalJOGsnM/ETJum6+l02unpQYC
mkLn16IOxvdZweHtkxzjChZ9ivzcptsA/uDdjJxuT6GfX7J1I06WjY7lWU7Jrl7Xk7F52QJEfWOl
fQknWOKMLNS45hyKHpF+80Tk4KutkYEdtkNELbLWHDBknZGyXkKaK+KpM+76wZ61UrfcEN4G8gCT
q4mcOA8UrrRxsXSii0xMXGqInALKZAx+oPQpV5E6oXafDsZqyr9o55pIqns5DRvopf1wXuFZOTAg
wnY04G9N7zvrP/cvfvTcHzMgCDfk06JmaKMsfdfvGGTQn6cAZFk8cz7bOyRY8hAt8ge3BtQZS1nt
2UkjiPJDd7JoIMAPL4jf1nbcF7hObEvqTHegBtpbRmOYW0m49anYxew9vQHVVUkkG9YsaJlhJtYJ
ue9WMgH+KSzy+b5hBQsc9RFmlpRj1rHhOCS0ssD4TcMTYeyT1w2qEv5XyzbC2AX7qMA3OwMuMt4j
0fuh2rHtUI0vZ0tcf3T4drfv2K2sw2SY93eSK0q1o5Y9iwe9NXkRoCDExIbuuO77SLgbH6pdcpH+
sWFzCxNZg5sGgJpSqgZ94PRs1tlbis2vcv5uJMCxHPh6zpqoNZY9keSZg3oKlVZp3wBMmMQa0Y3T
K9TLUjhsYPyv8z/fiDVuY1sU1ZMFzDr0armJiCjZ/BWM165sWsjwgw2Q/DgdXjznfhTt4/M3gzD7
wotNOR81q6YpxlELGKLiCE/4+iy886zYwI+oPbNDpMwtBYPOQ88equDNcZi+qDeYwdj/03IrW53o
iDhXW2k6VcjQ4yLfGlAjzZcYOg0oBdHML7xqqHz+sb+brcGW6CBUMUXmFvlm7RaMcCPBVCQxRJhd
j/qq1zELwuxF7CCRNeABuGg0mdtbIxDnOTSdgMfxBo0IQQTudBwmnXLZe50O5OIU9/sZqpxexcK0
WjbI0fV3z+oUyssNoKc8b5av11QND717GLLLZR/YwchgL8/US2N06XF7IBhGizmb0oAUlGPVGiEi
r7lpiCXVH/bxFwnOZbK8RnqjgwCbXsKYyl7ifTmbsMZXmfyIitcE35KT1lGW4abrYZzms2FD30eg
rwjktmRHOnVquGgdoUd3mYGZcMwAcQqvlgp4LkH5YpYUO3BtUFvZ28zjoiMML2UId9z9Sf4Mq1SX
HYkr5+O3Eio68dp2bxTgJ8OMflkX0oyvaS1OYAKRow8ioXS0L3h0DoveLwoHW2ErHFnjuVc092ek
+Ep8ppbnMYLo1NtEQkP5JjjFdsaSRNuI+b4DDxixXjTutGF3CFXuYfcf1KHuOYwyDMMF2h2jLfcK
Ine2X0mYmzrjpMHXtdhVDb0oN7FpEHF0KMZd5I0dNZerf0zssUrHosdiOnvJm0f8jFI9oPgRrP3B
awcfHpmW1RCHaw5CcbqY/JUIQQ3h3Co+jollw08o9DQ73bGmDhVzxrFGZypQ0u2EdkKdvh5CD+HW
DdPc340sJVOb917K3OzRChMgGn3KUEBnzbXmGtlhR6WpYlq4LQVY0wy6qYXZWxZA5gcu6ZBbYUfn
/1iAIzyQaJKBfvVXirdWHR5EakAc6UzysGzDCu0029Bb8H46Oqc5XPvToHEbeOv7d2ZWTGCZmQFW
+2nNohg3GHQmKhV3/zEzZ5ZbMJem41CnqsFHkzTpxKrhldSlpp9bhWJjP/WyU0VmLS3xrFU13HXx
t1KaFGt+u5+jMihtbJ+KIvZ0E50gq8Jto2vN0JALVmSBXChrQSlNAeo5VUp2bkKsbxBA/T6j7Wbd
rZMeE+xbn2vrmDUuYj3kTzAnUfLsO5uKIzJN0Iv7OC5o2rnXzUmVMNajCySMUY6g95F6mRfmHFte
xhgsWNQ33ZE830cLq47mI6VZOb0TPx43L/GPsPSeB9yuAIIJkmtnjGpPjhiMwY1uBFtMMH7vfet/
ebBUM2JQpAnI+riswgOiqB06wNXB49IPhYbs1MBBnGttI4ipW9q5K73Ec5RhkpYN3s16BZL0ovcO
cF5EZ7PG9qS8KeJKUzRRNTJL+BMzRLV051fjkiLoGlHhiFVlqztX/TG35Dseq+r8baoq33yGpHCg
DeMVNySpbsOeJXK+1SBEfJpasJKSZOr8r5YXsDAMyuvgXXydPTpDrDLwMI7HGQZjTAsAUMSFAvQ3
hXP2ZQG2fHe7C2S8ZL5b+QanhrfyhQD3jCTYKP62WWox0dkfPE1bopAT0iUrq7u4v+Ed/1j5yW3f
SGrkR+I7kybgGndGpfhNe2laAZzHFQ49RnFrfKwCQjgBwmEkIoAlmjkf81cpNwCveEHiZASaBwpM
PLuP//KUnB+o4Yq/Em5gFrdlustqgF36Vn+B6uQmaG0R5byr0QVIEzQB8xWC5UIrSZuFqYUgAfH2
s1+5RNnSuiTxc/1MO+6SgF0hr+ip9pEusenqCVk5uRhaY/HTA4EvxovcvJc3abNCocbWvMky1G8m
uM+0hP5nsZxOWi5MSgFMjvVbJmDcOh6hZ9P48EmQYHOfOm74MxH+HeFgYD0M+v4iptTemTGFovd3
3vSs9W+/EO3G/NTE4ZxaEKHXvoS0Jr0k+V7fPpr8q8vutp071FvUKkyFv02REVi5yeMDMVH6avvg
CaxlVWyIoBlmd/1CPq3J80aJlMzTBEnznueMIabecjTbWVJy/K2lFsRcyDLB6ROMvDBQ5vyPm40w
iVy2JeuHaBXWOfbDhh/xkZ8LkNzTMwRY13mVky/X4rjlwE0qxzbVnPMSrXeDLAm8KpiZDa+0nIc5
P652MtPkwdoqScCkjhQd+WJqhkwmqw3cqbFvd3mfU8IfwsnrVmrUrjLf8V3qV+5Id/iQChHl7R7M
gA9yfclYK0GlXya0FG4xvaxn96hvTcr9e5Tfz9G/Mj04DYah0FMoZW+9w1oirJWuj8O47g/ksBgD
PwJuiEm8FCN8VZJaetXOa7eyVuN2Z6mgn7mSS0TrUPpJd93B8koCyobgeY1Zc57+8PuWR8G9C6sl
r0I2Vl0Z/PdDbod44RNREKskKodRPWQan8K47He8XNMnN1ZYvZMVf5ZAiRN50Txvcxf0cktssz2h
mwQandptbnjMjCvuu145CZOGNy4BSM7dvWceTmP9zEqHezIiYgzMTFbpF2g5PPGdY10FbGtQQsoJ
xTh9wlwJsPhD07ZHtgylcej3M1Ysr9ji69/ReN063rT+9CT+PjCuUxtWIJYg4DyqqhqVLCFs8Z14
/JUcEyfc9axwq6im5z49C1DB0w3yiw3nLOEwSpQCQQkn0fec5zpslixIhyzbxgTWYV/ZNN2FXuae
/LanLhqDjZQFGQagq3c/ch2FSj1x5cYzmUDMSljkwsjJXcuAKV0jPWU2Belc6cKN8M2A2DVTD4xn
OFpwJ9WJLWV6JD/Of1fqTFacOEyj0h7+RyTFB4oNgjd7OWQuon5YC1831Cn4jKQKkSvZqPQI/hY0
Y9bHiTMpNJ9LxzTtwnbFGN9iSbsZaDdQgqQx9jfOHTIlDIuXKMFf0wxXrLTrJsZhg6lwzUt4I8iA
T7xFbVYQLwkH0mx3oqQWlpYas5EYr3cjeTLlpuq/eawRXutEh32uMJipK+g6oHufpGIexqevmhoC
tTKPvtsyPAsni1w5vDlH92ZoZ/evZupSSTYtabUw55lg5ksUWUFkR1nX+OKIKAqGqDLv2a6X7nKi
Aq+aUJcqNJWAfLlfv0Mnb0/KzuSHU8nL5mX1gtz3dIazijbOBnNjI9trYJubF27Lt0o+h6j6WEHT
fsV4ffQj110IoDdR86tQMj9B4RHu0gC7Y5SpbWIxJni4Joa95a4VeWQJ7CezxJyzqe5OrGw9Lppq
0agcLNMVP6ZCg3MXyoXG5NMMUxmD2Ts7gxi52Y0BVWcS4cnbHc2IVHkSfVGB0jhtiaROIgZKUpl/
s5PTht4qA3FQcXXOKeKrNMaYW3Pv8LtsUV/5spZ8IGvtMO4QJc3CxohM/bFqODq1YTlDw/IvJisl
9EVefE+Hcyjyvfg6ugh5bEBjb9uqPDjoiDguyQMk+l4mTx8558uirbkdT6KfZivMYAEqQzkdTIAZ
UqU5uRhR7R6IyjXRC3O7X0nbHFxYEEK/AAGug+aG1ONmCjHe12xzXk/7aWc9LBqC7iSyNeIQ8XMc
bhPYbHKrk5GEIUFzLoROCZpAvmHIfjWNOjyIgkgXGv6pM+6+Z8ohepD/v0hxtYOgKnMzrUo1/CUm
hn/5Yh0pGtaLGU5+iTdlNkRLXg8LaZ5iLMx2lOyS6YHhzxZ94Jv/jjU9uaQH3YDtmsAr+DWHh74A
HeSl0CvVGemIn59fSu/JBkZb1vEZhVoBUGMOYwPEgjTv+viB9GCogiT23u7U09uXLCzXtNA4sVsv
vliqW2LKMDQaxYUWYlehYbFQ4g3htBAcYkQ5OOip4Noezca69NlB6DanFzXHYiAXi3IZWX3SqDdx
apne/jLDoCXsazLyfN5nyF01bdWlPAw/zZe7U0V3PyyRzJrJTSnCEoceS4lNfL6GiaiFnuDyi7Cw
ohGcsAs5lW8TiydCfZIHzblXsbxwEISsfNarmKJ6ROITW4J7G962K1GDX8HOR+CBKB2b6Dx3kyCw
/BNvWn/p3rqQlxb5WptBAZlQ5o3/QyPZEWsIlsFqEKnEWh0KMRUwAaYq85M4X7gFRYAo8X5ByKHt
8lmi2RL6NK5/2XslWf0x8/NaKNy4hGCxElSjeKfSgKMg1o3FCnomtIUdn84/wdYfHdMh+XS8aw0E
XtQZdnHqgH+tkc3MKjTQMt8m0LRX68PHS2fXVu5/PRi5xxD8B0vaJ0BleKNbuZqcTXH0lm47mYYw
t1tY0ubEkLVVY9f/78EdsC2tK/pjMDRF56H8jm+ZVqlXyubfnCcq3aO9ZIs6HyDQbPl7GfbzuK4W
uPvVtXYz3RiGQ/+CLRVannRNsgsjt/3f0esrjbKqbcbxqk5IrJ5KCsUGDtYujPCm0TDBH994mBsA
I5+btSbb/EJCT1NoLNP/xtC0btXKPO0A0RzcYQkT9jwPH40HCd5Qg8PY33z4Nl+2QfmJuZ0YOa9+
T6itetYWkiPqOfvY5ukoqpt0pRNNkUmeDpnU/4s2hl8B/IZZ3slorUQ2/0noUEHtIQpOoWhAfjf3
Qmzd3kqEN18jTU176KEkW+lMH5Qm6VVkuf6TB7t/9gURm2opMuCG62+q7gTy1exrf5M7Y6yGi0TC
QA1Pkctajl0agAki61Yz1Onl6MC0sfVtoGy1x5hzESiEEFwEUltx3Lqu7jF1H2Mc+XJL+06rkm/g
vHs+Ddlb253rpc1ly8cwGn9HR7lk78St2clEj/rg/1JoTj7m5zd1xmjfMiyVOLtRl5XDXFKh6Wig
n+Il3HbCO2tpxdrqvvsLoEDD9UN0T0ZkUtj6suXsCaWN8eKo1w1vVNLUCrc5J8t9KbF7IW/l14+6
fq5HCc/KtluZh7a0jt8XEzBtvnc5Y5SB24FsHjwrt44Lg/9MMGvCjghAGj2NFAJhEgufOFtqtLnR
WM+E77VfTDYs2agiMB0LVN0yCYBBIM6cEUZtHSsG7euTbNsFVfeKM8nQE3w9k8sAw784V2eWzOZb
IJujp403mpT7FwIFVnAABPjtVOzwGAOayxyndXSKWJjVc8pOhDOMnz3q31SeoCylNevzU+B8eXcj
dtj8Z5JLOarfiuQlujoH396tLXOdQY6ludJjuqrwbYLDn2S7vKKZrNlqqSS4F9wRrwEBubTjRNgh
oxeocN1p1yz+KC5yP40XwgZCc80BJXFN8X6klJ6RThdL5jFxlbCrkbzm5ExQwWi/9RjOuaVeS6ur
IQDJrgF27BwezQbIC1i4DefcPSRSGcquEyt1soObzNTlE+d144q2poGdF+b0X2YS0aA0UdLIq1zP
IvT/1Da8TlGsADZy0qFknUWKnJbOiYRd8sIcwlrChMB8qXwgfJfnPfaP/p3cmyIrx0KcNvPADCbr
TJuuPyIyYiANJP1emGp3mxVJvdsVNs7aLHMc5gJ6f583k14Oezi2ErvkjAoA+YfsYV6ZlCPGyEVM
f6atllucKuOKcdQ0G26+Z/Mgj39SODmsAV30yYEH6F4g3gUZ+/r9D1kJ2APMhPj0Q41uh2Xn0/LT
wBLzjIGJC0Hg2wXcw3PC6jXw9VoicGiYLrks0JeaX0HAiBemBSARCI7bhkQwJqCCIM6m01nVUEhV
637AAPAJDDw/lLUJpQ7YsPWvX0hPEdfqhY06enFistrbGXVWwmGcldMRTZHmIPvYiPa6SAWasRS9
xkW1yAM51UHzogGPzSBcQ4Mv5a2IM2iQwqPiKFKif4KoUrqzJ+80XuT4bp2n1Jlsf1IrJxpnPgb+
F/JWpO2qj9T2jM22UQrm2FOQ6fsCNkM1zGTygvgviqv8C75oWNcX8+5/s5P6BsKy6q9HsWDYD1e3
NHs0BCC9qHcQO2EdpG2zW/Fa485Pqt8SIYjihvmPpvj3gmeSbWfvlNGEj2iIjm/sfjGo11IswqBd
PScepvLqAx7m7RWQwjUX9ebc/JVJTlgikkEBcLDHa05kgf5OMd2dKDAPJ+jOtMrb1f7jG/Eh+suN
kUgvSSZxR5TDjGPJLRF+d3S7N9LgRWxx9/QHeSaXi6ruvFScN0KrEpPRpzxAWxue0RDuGQlOQ70B
GTyTHLeswYLZnH8AcFvMhpT3e0ijo/LnHgyJR9bNsI6S0Oh/kaO8oEQjRK1RmDmt6olDF7Cl6UnA
/GngLW1tD/QaVMn4sR41rodVMOoirgzk2da0bZoLVzdaM2kEq0Vv36J8NdjraNu/elUigpyZ7DW+
chrsBV0e5MA76rc75WbfJhtdCSNt5QtY9HmAeqhKQ29BlogmtZo7LqJcW3KEgQ0yv0PaQZCyth/7
pllCQ0vyv28drx5mHyRlANq1sBE4VI9Fd7kSvigdGtMvMAtciBPZ1V+dl5D5gTToDWjFAH+NZgxt
tybSbh/rva40o0h6aousCq/eqF5FwGRyun2lFLwNQfQ/lvAiXN3ctmeOcHGBYlu0gKddrWIu7K4j
PlpipdsvUEyzdwCG3A5duv2xGOfX2R26ndTTc/8/9mpztzhvonZbLYuRx33MaCs6fTWX7xNoiOGc
APGeTgz+vH0ZnzA3bebX6eqJoSzm+LAuoT4+IvChFlCJYmaOBK3KDgzs7UTjqmklQQvJpAxeDndJ
oEHWDQeHjk1jsrQfDruwVepEx94dqfXjEJNLzTHAQYXeI4I7wfTYZutqjB4sKWSx6nGgmp3ljy7g
tE0FJmcY/ZGrx2jRCPWxAb1lW/5XdkpsevjLFZBPMf0okiHACyz19PAR5ak7+Xb/oZhqlP67XqWb
S5Nm+BxcWQHp5BXnbLAOfRW3V5MLZpixgSnD7JjQ+8k3AEfYqnLO+8Kf+zJxcnwDnyfydVkdx/6p
CTvNCKZyPUtQkxqxJ3HVsWulX1U9I7zoovQqqr12I/5+0SUue3CsYv+Wq4KbIL60o0q3aO6LY5QD
z2Dddo3o3SNkQsoNFJNXWMXr9v6LamTgNYHN1Oeu3rGxmvc1PAXeMiwoBVH4IScr8afDK1s42bfB
YQdR6xH0DTbHMLmjgyX61v6Shl4M4cljfkUNs6fHbB/hDyDCF8CCIcl3BzzVbx7H8KVbShpE4ehP
TB9gXlprDooOU1eoiqHccEWJm+C5Xxxs0P/Qg9PuJEx6aNsKfrtZzR0+oHqfCFFND0gOM/ey0Wis
FodZk4KkQVPjsxonOeO/eA7ZnfWYLjJuZRG+f0TThX6qjm1EP0mLBJLZcsk16Ig9mS5GEtXnX8/Y
0zSIIV4xGTTvLaWPr8MMlDXd9gUntOWKjeojXC/Rfsx6/QT9GWN3IWATNPXg34C1vypOKSuvX0I8
D7G+5QhnRbNCpXHGora45xlqb577xlXADcuVc1+JEWDgPMsfC5Pyx1SEmzeIiBNFqpup6i187msE
2TWoxVY6Uk7Xl5F9tYVi3cWtUJ8oOKBhNSd9MW8ygcJhM0cS+qtmDEcdMf8qOr7Ol8Q4jb9UxsU6
rSpnxu8eAqeC5H8H7E07xs/q/HNLDNgvVOx+4QHmvufIoeeNQxdPhp0yKjuA8xVZAaSdWqmDU6OU
S62TNfkKT5fM663LgV1dnGI90WZT1EUpuLy8UJK4K2gdCHW+6pJgo7AYLdz7W3G1lxxlfZPhutJh
dPaoWrzNTTOKrnqhJN/HsnVYexDYR1vgu/alp5f2wPXvjninOwGOOrfZ9zGIxdaiCUvs88TVeCGC
3ngffFHn/hRocgcm8YuORrZ+Bm81CfPGHa0YhPko/x8TNnInKghiGYrHinmL/1RRhDu6PsR+Gxbh
gJRiaL5PFKph0HGX3dVMIpSSfr+wCNrOp4H/eTv2hvmN8AJ9YAXq6iJFFMIoeLQ710OqU9jSh81T
HAaMaZWPmVKBDdimUqfn19lbqZoNJLfj/MzBMLFi7yUXa9HiVOxgf4F/Sb8D92mMmKQmNFfcNQX7
J03uW9KMNe5o4NkerXTuVlB+H57wI9eOOtHX88grZ/QkyND99mhxNVUCN3NUthAOFCaCGH0EnYdO
i6iAHG/5rgg0KwJagn5eqNW6Zw0rYHW81ONetxaErSMYffimdfiY8fOa2BeqdnzpNpL7BvX8MdU2
WPU49F1kp3X2vUlJlAgTnCksBt47E4iEpU1vEJ0mPDHbaK2mHRBwyhsgDdTBXAgylz9Y5jSqKKJR
wV56nxq/pqB13lEjPNx8eLDFyIcB9uaH0I8hJ5VAiRKi83CP51Kb2aVTcYe8MprJi1/feFgNQNlD
JJ3xtJqsHIK6j/tGzl2o2ky6gIJvkqcjjWrPNoMVI77zhLrAYA9EVBVNonuGM3xxmKjLsStDDCWX
c/XwCvjzEUXelD7rIHsmHjD8+UCOC2O32xKDRQ0H23YEDquLJXmTHiRHwvxUXhGBJVi4+XogNEQs
Y4OxgAGefm8OLLZfykvPCayi3eObUrABbz6Ws1OZXzAufhA4AyF6sSrqQ10WWQVq8xatZgirmH5J
4d0+eUqGyV5uRc9iEc09mWXTm7k3oYTEhX4Hs/Z94t9vOIRRJwinZHqKTVzvKa1Rg9O6JiQpCFbg
updidhkc7dD08bfcZPVBJM9Pki96hxTZnhzk3WM2I0ReO+givqJZiiRdqKkHEQyfdKGlAYODym9K
DLrjJTCSY/Fbf3Qjl4Rp26TJcoJkn0v1OXux5ML9WRDYThZLv8NaG6nTpn/TAZ57n9CL0LdoHXd4
z7splNcXViXVu+OOtc5FK/B3khfIf07knnr3nw+X7aBITD95W6En8z/3ceZtEeevw1nj5Sbd6YdT
zY1UgVVRhWivOqJsi+yokFmxqQWA7clmLGennhm33k1sJTsCejRwO01am+3ZA0yNkXLkazDmTo5g
nnriAnPe2D69e4is0Xat2hZgFVJAHtunskyXwc/n4jd9RiLfJrSv9FWVkPBSaowHlB6hEcvK1/20
B5et2LAFteQJqvkWbrdw8EXvERzFUgZyrA7AKp3Fi3hdNcARX/4ZFGxQVSPpcmaY2GY12+7wytSp
zvgT+b2UTeHQPZHX8ewinKPrMb2F1MNsQcYFIHIrg8y55YL6KTEVHUDwvE23PnmYl6u8sexYOog0
mC/Flu1OyThSjZC8P3XlMZcM89vc+6bATNI67DMUK6vKQGhVSl7CR26rpZRfHsL2gY1ApwqSqk74
G/TC3YODZxbZvoPFPDG8SN9IDUJc1Ug+pXvHfQD/O5B9YayltGGNM9qr6zwhjAbw+ezC0kbNjx2G
YQFVUjuwEpnAoH9MuQNh7Wtpr7cgnFCfvqWjZfHGTB69OdAbr04ArWmx9TE+oReNmwY9y4QTWnil
Eg9XVFIR3Bm9/KBo/YFPOTd7Y6YRUBHDW06upZcJs2d75edQfzEG+umE7ppWAQ7gokY78cQr6wzm
tAW7Pq/i2IRXUiSuCRlHAy154GPds69MnBcBfkKmSOMV5VsPHU7TzzblZ7+DyQ0FnQeODwCQ9gE3
c3Fs9+CYT9vHYhP/dgxm9q103bBNtYAgolFDcsgbDrvI6Tzv2GRW8loYhWfs73xRoOtg39jRjE3m
DCO5eKCsLkJPk7/7fGrawKqOAJleies7INRsZieA/NkTQkXknpfkgVUAKiXMcq8bWGcvPBwh5PJ0
L2gwuadzl1LXbzKsIifhtZN1OqJZzsAilE0OMkWgsx9d/CHyN8+n6RFMfoFB4Uh6OfRSlWht6IsV
bRwS4xard+bBQ0qKrdfXCPSiU4LwE/z7ypyAFXnV4xZHgN/MxPGbeCgx88z4XQX2KQl4fz+KiIYx
sNbBmp1WvYPBYHLAVdFp2ZvZCdCdZy/vz0ifrEmSIyObkuk9kfz8qk/wnJPTWjrUY/3Q/PZoi2g5
YUx4q7zyZz9kYJFRT4NpKcclZYgJn0UMsoH55L9t0ruBUrRa2/hsdtHRhdqHGmWaquu7d4fDY4b1
ufd8sBLuGdwQXN9E9rQl6pOOb660GBhIkHHngeGLFyhzWmhMs3Q8AOXGhlCmNkqvgUsw6xv35P7Z
xEunyoIzyZIkPPK/pk5tT4oOfBToRoe9exHEq1PObfn9MGs2kTDAi4/VhpGYDRWnQxLU7KmGpARh
lO/15i5dvubeeeWfj+AbueXZcR+cQPs5xrSKCKRCBpgRJsKDxX4W4Vfxt9I/e7n5T178xM3ih4t9
tWpqJwsbcjeY1RLn2tt1gGIJeAkgcbELmZoj4D7XoRn98FUBgXX1lRCohLWVpb7fsItzmX0uRlUm
VW8eqTL7OKfzxDfx1ciE1BoMYeeHRIGPJ9ve+/jC2FI8ToaMGTDgWmDDClurVBl+XlyVg7OtzYba
sATNI7jIfGnnUSNdG97H5k7qg1fthLNDyeyE6A90MEHWBrZaehNBke7F6jOQP+p9ARcV1Y/2sE2U
3ySngjdi0VMUEgUOvlu0D4C5sf4kncmTAaLhFtz3objMOiPKwXQZQuIJDtrA+YfF8Q4DS4Ga7cIe
jB/0G3/K8HJxvASg7YSuSSsmq4wk7YRX5+hH98DZOYzk3oHkEq3jW8rEQY1OSXqsyhJeFmBk4j9D
7mJ4Du7Srm9OU3VVP3onfpO8WtYpnncpwu5CG2uWQVf2u38eK0wV74iwxmXucLXyqNkd+0Xata1g
PW+o4Eu4u+gbI4u5YQm/S/z2Aasvii68MYgIZdydK177v5+0aj3TOzoo4VUlewkH5utJqfwZzyTj
GUnwAs0wp61r5RDtkojz49DZl3W1/TaYYpLU3YwhjtwLGoLDRZSDgUJdSbme+3oRlRZ20D0iPoK6
Tgmd2/zGEIkQah9/fDTWuuoPrF3tH3NTCi5XPqzikxhH0XGyPlKRIKU50c/zrlEHruxrFnO41a+6
e9fRpS9K6wO6huI73t6un3wNUl6QxbCf3l5Y3exRphhICXvU+exniMq5dZ7sSG8JoYnKFhmDZ7+W
wux3GvDX5+s3T2KO+kUEbmeczLr0cMMmZLCN/Y+JkyUi6vuSv94/OmDJIFNpjkmwd3q/432U9AzQ
8oYIQf3DAZ91SFdw6z2Ni+ok5b7W4Cyjc2VWmz7NZ6vkLpikreq19nNmBine2TWQB9dwIB/Et38K
SWLfmaUfuvCi97tLNdLDFDlHKU4gA01l1kOiwKAbeXucLRUCJONbrR6N1ku2C8vHVJMVOCIUotok
MLBB3gOrj0gKrP5yFBF6Liorb5LNJxxbFtOfKN9sPE6Ou6uBUpaKWxmvwdF3l62e+Vju/Hb7odVZ
pwbMT90sPCs6/PfjSpleO+EMVtqYZKr2IHKMjQ2UmIbNgKB38PAKxH+G87KEOFlW+MKbalssEcs9
MgguFYB/ka2Y7m+ufrZCppWPMq+nO0ifxQqqpfA1eCJLMSIHcrQ+z87sub+eeN+1eIMhmOX03Nez
fo/2S3XbV/lRtzLm1ksLzFaP8Ss7Y12cD1Sch2NMC0HfcrXpS6V7lMukugQkdjrrdAfM9F8ml0X6
dsVW8YPRPXSRsEkaG9wqiT+s3iEkxZjOw4K8ycNZjHKwal5uOyZ8Ykh6XFL+HtRmKNGvmlORLht4
NBJyO1W/qcBCXdqoxdB+6mBXhX7TIb6zT8zpHAoWLGwrhlhv5khWT16LpOOsSZr5An9y11aWTp+q
ccXoHbaBSWxdpTyisMeawlbrIQJhiAU/fDHLsoCBBaavWWRY9aGGb3j5CqIBFXEzpV9Wcp3FlPjv
LZjrq1zMLc4MBAb4Wjj1SPPo7S8J8jSimmCmk0HOwl0jMg9iYs3ewdJpMrXZ9/sAqrS8ptG+xUvT
MKL0zi1TZhRNMVXiDB7n5ciLDufYomXDz9em1GTMgQilk5setKaHwrTwEfyfXc+jurt2cBlqgTXG
3XfzH20VDdVu5XoNrmmKQGIqtp6Z8iTpVnXNNZvGhrNaOW5dOeIgmIi8WymfJc25OKb4iy3J7wI5
rluT3ylGK0EV30vWsj5mHuZA9k0vBuw7Nzjh1GaoV6KZNGS9mrDhTPwH1l9hJhYIGlYRTARgheld
2MVTkHZmp1+2t5bBI9v7xgkYysAsk7Fv3CqQBblRF6VXuF7AC+noP11mE/bOh18uo/tK8k/X+ilo
Xp4AfTOmUA5qdqah13Tp4zCPDw9xoAw+p++HYEDTS/FWTKHDJdW/w+MwWlwejZNGjRA+LJO+FEuy
SMtad6qRIZAvTa2LSH6xvHqC7w831jCThwgMTxY3doVdtj4S/yNdsLKjOg2ORIENQuRLXGsvZRps
I0Q9UOHIarBzdXW+b29xccz1CVzTO/WHt7PvTbe59ib8l4vsb8ufNUqzqeVL2VxOqVes/55B9CsI
MEfbAq0SByiooRgaiNirGm8I/evlVLJDdPk7QLr1KyzhQ3BTlutUx1dqvlXnEdHB5J26zfLN3NC9
s2XzfIe4fPDwcvErthUFMNEr4ms6WPwBdY/z3XSbb5iKWpiNLGUIFPD9Qxro6XcXtScNBnazmicq
tqT+mvp5X9/UbHAB79eM1DNCrvq2yihGo1MdSuy+EivXLXV5lony9O92rnCb8LMGhp3yFB98ojbo
a4JmPZZo4mtDTxLNfDKhvKGe9txhOtzkGRqCrZ1UzbD76Q2ozR6lZ6OpF/TTVZCj4MEgBzPZ22V4
vB6KuL6v1n8+P6vDz5WBy2JREru4l2+3eWOAgI3+PCK9QAojmpLUctQoDVBgvaQfFAFWlthyKSg3
LHRbfwGx2JWhbeOU5pufq52M/3Zw6L9Do+1byShZTxzTYXcHlGkIKalhRPq9oLFFyf5OF1ItvWOC
AGU5QbZwEmRW9SewylrKur7V3MieRnwpTMlwAnYKC+DyuWdN8GFWhJQvQ1y7negLq8SDqt2Kpyh8
4e95RsXunH4HPukQh5A0ikky8kIvmD/uXRuYP0Idy4vgerCOmhmWdezr5R6JU5uBiBGxqzWYPG3n
jm9xDhQoiWtgJbFtmvZoPBJ2m8ALIR3+FR9ezFFrCT6LUhAQ54bihz+iuG30RSrsgdZMpIaGKPt2
N6Mj6QponRencR5bByHgRJZ4T445aBtd2Gi6WKxNWfLlGUsPtXMki63tJtcUBprLZilm81PZqY7K
NUjhLJG4YnUgcS13h9oX0PejXh3oomzm0X1E8nPj9XAcpbQklFG3ruOmh3dufBa22zghmaQpJ1UY
CBq9BOnEL+TeXkQVJNZDV7zO+NCMQUKit1FwNAeiKpu1C+qnr2YLATMQ/YX7LQPra9AMHtTJIU7R
mYQ8pUiGYHPAfIRiHe7DkmEKzhSDW/sdCP8N3Xb0+aPAej2hEafuk6hrFbcwQUv5D8hx3PkZUjGW
z1+d7D1to91V6fXK6RVMYykcebgHukzDQJtJ0M99NQIXuj0WUkIgLdI3tIwluAAv8mDI6/AHxLiz
IMRKieRfHWD/ysp98wXGtwVpu8R4xrVdX8bZGqa0/lY3TqTdQUGp6M9xrBV04FiqPg/SDw6aTUzm
H9Vx2rV6K5TXSk1PENnQxsp/uLARnNK2QpvnZGLDqq0OJ8Uw3k7TAqz49+ohvCaTEUw3Z0ih+Dij
0/p1LsxdxbnyvoLAXnf0GJez0SlNWd2oV/JRk+63aSB7YHSu9toNoylHKZNlytKdX4olnuVvnf0M
qFMzYJSst8i14lGMZKiB76zoscNgP7jCkiRTKgNon6lR4NKoHjhjx5ED/xz8NM+dDKotYxW2nr8X
8+ycI27b9MbLmEXgX3BCE/xUQIcqzl277l0Q/5PFb0YPvm/67i9fzlsK1dXmQMDTnVXTaKYpBHWw
Kdw//2q4VAWDkzzkx1GrOshUDRnmiJnOnFwKjw92ICUZ4jBk0C26VQYiRgtxQWQC7fYt9c7xfR1u
/4BwdV6Bz8awP2MiNHFVYb0XXDVs4MjpmFoT4yHSPc7xfkekIj2qJbqJymtfDqtHK8unhFsIQmV2
MPwLzGW4xqB8yA+kL4SNHHzGUe+k8vORmjKgu60LpVttWbgOK4QUhLMn2pBbAUeMMCLkKJFj3R7I
XiYgH3vv+T75pv3lRkRyYCvzCbLtf+b61nRM0/M830CzyDEWEcbXkF+RG7hRg8AVg/ZgpkDWRa+d
XI8i4/WUGbf0GoQAFlLPMOku/0r6x7QHJSon4PU3p0+Tpc3rsO6nl+OcwdhjbO85csS8cinKImf8
IIzBltWvr0r3zN231KuwMhnAoBACNfcOakwECPZfCksUY97KYG97KLXy4k00UMfTTnQra5np8BbP
skqfQhDGGo2s6bdBtzXdu4S9V6E3rWBDRG+XJsbylQDD7wqh1hVlsikjP7BlPm6rabc7TUIHIlHj
5TIFXRB/j5tmncJtcZbv/GH4UZkPmaz8hpGQcicdv2tRc/GRz8gu7udHiaUWkCMaagW3bZ+dIu68
NWXdyEQPpvULT010cb7LNgDTIrDh0VxINL7G3Ks00HRGjPOfeoExH9qsRQJF1JXTJ0frnocPyIwG
FZP3Zd1ua2Vq87BWN3RGsYi27YB0ilEwcASB2eDZEt17KdRFquC/gC05HcxK+Jnqnw++QtK2l2Y9
kPMYq9tHEs9a+9c7RC6QQXyasXBhpZvxVCNSuEySy70GEiFIoK4SOn+2ErBE22wKRuOBlRFScTcC
1FqmCOdN8cDr+Nq4LtVgQ4BEGfTqUqsN/uWKWb6m2xxeq9JQnlVkuP+z0eqMa5an7vEJc59stFdt
dl5MuqLGhVPLTVE5F0noczCecXPnX20sIGg8mMLOcetxcnlGOcfqHTzG5UJMqxm3seiDxW8ANFGr
//WUgiOhAhlvbUOrMHHUoAs47IPsTGziT+IsMRYSSu/AvuAmPaEe218FsHYDuWq5Y7OESujzpPj0
HJ8zZPIvLpcibf5lwu3BdLM+gHfBxkgrjWDuivJZnuYAaJIjixaS5QZS9jGmWD7Sdm9Qm2IcjpmN
W2Rc2B1moFrVuwfg0mDy5s5s681ydea3ESETKADrsTCdu9eFy0rBt/V14zu7GeRmFAjAi8jIADpb
RCVekaLZIZIXBv1rZu7XN0REyfM6hObpO3FCUl3zD0lCtvtwKAs5WnTqg7moTrV0oR7L3Q73iYzX
i81TzOut4SGsIdLPdZhyodaLgSk45LwG1Hi8OA5uyIf9Q240bHPGPTnWdvnzG12fBHEo+X7P7cRE
Ypff/PEedwjNg6rMY6BbuKj8es20dCe6zVnFM38ovaW7sjukgeknrn3llefVcDmYagsvycol8Ggx
K/Ris7S3I9j7v6x9zE9q+FZu14ntjsC4gJEzF2Y7A5x+vx2yPeIF0TJwipV7WzGLy7QE9Rjk7FzL
s7kCS7YFx9UXvXefA5NbxgR/u5c0arOlVTvrOWfVYm2WfJJ8/sv7Fo0cEFmNvHz/UzzP/SpyWode
nryqXsfxFcrLyhQfw79T28fYOi8ZOze52b8ix4RjrPZ6cfMdlSN+XokG8L7i3I8TtreBzNsepMhw
PiKjorFUoNZLEoylj1f2EMnk7ed4f9UJrXh8kok0attZo4KbnVBt+eLH8QDrPLu98ESPO8f3iDmx
J+w410Owzrf56Rl0UrH5KTA328yBZ6qPco8ZJb0quiFTy3om1tsVOuZrivrfOFYhUGtMM3tAOjXY
EKUSnm3GSxbFMWNBW58+tCpQYC7brl3u9scp+R/eWNUbyNGsWRDiqg3RZMUBwJF+38AzYm8nQY6P
xSJ917cUfb4tkAtylmevpmJpOV/NYvOGNP/YzESIHNLL3w329wWk47/Ms4Qz2tJnGvg4lP8jUs3/
itjE8/UPA/jxLT5878vJi4jmBHY4f8SBzO4huWtij9Ff4f34HBfnZzkf4suS6yoEXjZfbpKCauIq
CUnfjImoUeKo/A+QLU843aygsA4+uuMcG5gcDx32LGRwCyc6okamLz9JphelbCNA1X3FxOiUDTqc
JUURwQRXPbaEkIhuGmSKO7Jh8lrP6FYtHzOB9vNR0AnCvA1TaGLfvyXAyF5oZJBRUXjirNw3jhsA
XDQEKfdAgJK4DpDZIEiR7tMy5Uhi96vjGyNyi9cIjnXc0E+HjAu6Jx3xS0Ovy6Tjyg3m6I/v+Jcc
1ygeTz0ujkcZYuLpGIiNyUaYb9f+5tixHTxXgpbegcbo/jhw8iq/gxa26VF213I2QMSlSAuoDxL8
krp45GSUYaI/PN0LDumzhhm2hrlFFBaTGUMA3eWMFsS+kg7/HPlMB/aaWb2rc72spl60QRO3ma/j
zq+RNyR1CZy1gZPazmjXkGr7GoQQqZB+QgWUgOmu1TRlb8sLJak5JVVDu3rLJSdy12Ame5HgBXwH
I+/YFYyB43c/CmrUnbkmSXSwfOZeFchx86y+mLQlsb3jWbWiBIyVgT0siZ6WYogSfO2jnCXHUIjJ
GqKxwFLtSEG6xkqAFQiFVUXFHnJgVGgoJfjr+kCUDu6V+QeMVd64YQrr4vWsGjEr8nvaYMiEC42g
GaVHV3ii8aPc0OhCvudgoS99witFMFZwW6We4meGfhWtHqzm2VqzuEke9xfjinOAxtb1JDnwW1TM
gVoGOfB9ShPc0GscUclVezCq/UI6VG2LtXlpdktXCYLap3V3IhTAaoXwoH5CNU6w6B3aUq5xfDJc
R8YB4ukyAfNFHHfuqeEppqpuY2BcMK9rSpfCRQy2jPnWlaNCNtxU4e37V7QSD7Ii/vvX9ajS22IQ
RQC+yomsgYYSsqGiaKZx7/TIdraIVT8E9VZqPSICfASxgRaWxTyF/LJ0qkAO3l+jwF5zt74apJ8x
JJ+zY9VOHC8H4QwHadLeMntYa9mPCjrxZrV0zLGidl1906joEcyUj4Cw+d19p1nhlBH71qtRT4qK
mmba1jwDOBOdzrnnfZuoh5Mynqqo3YFVMbIYLiB2wR1wM6bEV9pKIxPi+HTsOYFRF9zN5W7yVDpL
9BbrzwkR1M0LPjSRltB2mmeoWTuelLXcLaXPwlXMhVV+baAzRaItE1qZ0b3djw2sAB7Z+QksA39p
UVJMr21xTklCz3WrtG2FgrIP8FkqCP7UEtWHcZhtdzsNlzEdxHA+eFEcdU+SDZgg35xiusJ4lqSu
4L9sAtY4F+xanHuHCQ7m4KD7zUBh3MW49fxtw2/zSBIZ6qsnQDoVnkX+4KE+3+xJAgUlYlQIF+XG
wBYYT+cK2IMHDmeoEPW+H3+aTXdOqApW4fFTc9+oQMtJktMKup03IkCbQ0KUDXRNLpPYbGgV7V29
nldX8kG46+grGMPmfGX51KAWCTfSbm9pWEatd6i8EH70ISw7pPtsQV0MNSF7OjnXyqLExo1R32+z
r/vgyzOv665A6ZT9FfOqNg4zghcwlKpKVkdDzwsmEitikL3K4tgd1vO2OdJs/KkhWJ7Ls8bfacEd
JglAYr02lwr0q0gTN8RWHNZGDgmzRC6tFnL0+pMFPwkLRoduenAJS2EZkoTB7TAyTbeDu8B+yRh7
oGiWh7JtQaCQr9vI+4KntHAa48lOIdKThO1T3cB7ZqYhy0DjopMx4hPEskCxCfroVaG/79Sl/MVr
ZBeNHVpsL5n05ScaZFZErev/ka6DM0NkR3jfs9h8rZAlw52kg7wPicHoBXbGvH2lqmqR9FeYFN2H
/4DpQs3GbwXgsoMKXASCQe0g1g+dVqa/cJEgx+FCfgjrgnAnbFYKfFJ97tkzipqXzKD5YWgrOqao
BwmtiSlnBg46qrrrwc3soDGrANPb3qXRVVXgPmoZCQwSr2bKLpo90MKo12RFZdcJzB3c2rIZqjTk
YFlci8R28ROQZADswqEFTek7U2N07FBWrTlChuUymHbzREW0jWpHAzdNZpPXfc+pQkLVx598BcCJ
QMBElwAaPb3hdOnP/NptxquldpN/Gk6gsnMhsV0WsbmZr93ywdNA9yuXajC6e7jQKiimxJGGBpFb
wVJGqenNl2riic9GSSNiV3My6Lttk/ROa3mIfn9vQRuMhcH9jTRXP+++fGs7aiJmPRnLtD8w4i/1
8twDBZyeffmucc8GnayDCEhFSmJkYoOr0c2R9lWuruBM3AuQKR2Nw7H8O+DhfutH2hIoLWuRjzZv
KYN6F/8GjFC7tPPNRebnBAY+YKattuBUqaZYMtILCFJ7W7VqezUjrqZs7GAA8Ic3v62f0uzKoqHO
uDkWyyKGXHfz+w5yk3+gpbVzKtPdZT1pWg1ardk/ca3T10V0mJl2nfroRVsJ93i8KyhWPd7Tqv70
/9sY+JJIuhuWOICYOsQIOGBUnPhcR24hRVlMd9GlQN37rw+Ef+ycMu/0w8QkyeZEWkDeHyZ/MzUa
BnPclVdxVGJpoUqFOzamt/F4UP+ANZJ2t9UGaxiG7mmdrode+hAmT7nXttga8ZsVCHfowzfA65Ll
336bfG0jYGbQzGOexHDIu7uYTGXRArGX6l93RRWbNllVN75Jpj9ITKypyIVpAtJ3UpyKawUr/hKG
ZuoSxUHBYp57nxFhrGQQ2XRXPD6CZ0ru1Layf0vYQAwDx6YlnznXWpAfF13Jlhow5gOYtmDzah/8
CWktzt7rOOj3FxUuC8uZPOjR9D2Owl9eL+mokdZdsUz4BDpKzmcA1ZVAS6aVHyy6hE9UEfSx/504
54ytfOVBc08YaUQil5XgKx5Ls4bESYrlJuRg9GPEaNmCSUZIDgjHnH0M+Sz73yuTDOscPhf1z2ms
jlwSjH2K9abgbsPd4V/3bnopjcG/tTFzhSBgdE9Qt2RVteC4ZiP9Mwqu48axn3AHdRr6RigSDk7+
gxMp4kD9A/wXucoERVzyX2W0r9kubNXqp1P7DfXugVXDOErKQwFtiIQgVJcwmiVoODpY7FqApDpl
b+NEe/n8z+ANhfo4JYQj42ioYpA4iMbYOIUqSwwFoEoY+pmr/D8swx+5RN7Z6bktltQ0MRAqjTIU
JjwH7Mn3TQhDIBUYxS1AguwTMWeXllJ4b9HU3SXh+T9xkxEYUg4lWuslDFent0NPkwwSMl/hvDkV
NHdsAwHDLibH5hQGJrdjlMvi9Jw2xlnxKEcLPvcuGh/bPBtt6ThbhoHHATapj+i/0XyPyo81hAXb
TGlmEwhwYR3te0Auk3ayEB9AggJ8DOu0dFYoJcT1Uu/JnlRS727TDNU6Ir/g8hWWGo9CBS3Wz5Hw
iRmkEpKipi8c5pvRrmUzkTvnaHeocSkJfHY14dLloNyWWq+qvORJdOBS+mrQ91PY6WDTEmZ6u6WX
aO+T25GpcsDggMjZnoK8isCNCGuolB6CzDNSLE1YVgLtuZuInU2I7AtWiRbmYXmCwOkR2wEne99g
uvTp73RUVI1YQmGbbIiDlx9/uVVLmzDLd8v7CpiQWtrdcfooFX9VVE+0X/F6SAVPUjIBXKLM/OIA
Y8ZeS1VCSxBiTWm/dGZRTzRyQ2a6JuT8gkhjIqkEki6TYWPC0pDK9Vusznl62nJoJAwTvWyzpmd3
cmErS3q8Rfd9D9TF8rALYjpkKrb53/ktC15gVCM1py6sri20raaUeDDWGGPOM6rqV7Z0Hhh7YGl6
O1a/ZboN/goumLPpN+y4Td4ARbiXm2FMQvd+W69Er0tMMyfn+aCueiLNTvJvZlCtVESd3lql5dNl
CXOm6Gf21SNiF3qk/i4JlR+r50G4WFMgZTPsa5GTss8bMRAnn5zq6oUR7Hu4mguuJ1SDKBIBBfc4
f1lZsyLW2f+GVT1dAbQxtO659uayFPkdYLhe1a4ZBUVolhmjlWEDiIVKQAkOMsDCnlcolVB1ZEdp
LBmYOWSpmFoRzR0N9ADeGTl1CYVKehtCqS0P+NKlnorhI9SGanaIKgvkMYi8id36PxkD/A2T6C8k
R+/WfdWBVhYXPoH/BEjY+G5ZAhCRJ1Ruy3jo0PYHWG40KCGjfQKB0OtRInOdmtEFxH+XFVBEFh6V
f22wyQDBHUCUzKmWGydJ7NqJ9AyZiwx6q6L8Sb1fPlv7NDS4a2/SgLA6HRjTONCuR9lsJHa9jFtc
wj/aOIktzgU3b6QiEWdYGC4vwa2cPasdMzlLXwhqph85A/FmpyPI3YjFldmEEIqjTi6EgIW0D3/T
dmBUdqRTnI96WWLbowhlr2bHiX+TUL6uYL55L5k1tmtokdaoCsjquFcPo7S3WN3g6kENvjXpuVf0
GJyPciMgdvHL9Ury0j5W/a/YUnUG2rX9cP+d+gPUx+B9/Fk3QaUM89sdmsJW6knL9LYIBWCei9i7
dKXL9JasFnK4LYxpC2lVzbAjjUUPmOwXdtjc/XxWc8iWnfDzIDrh89ZCGaiF2eWmlRgp3skhDhMU
iRdzQIF1Qm10K43b11eTjGrWP5SUNto6JroWw7CuWSX/9P2u+OsOs4utut3Zt91Ea6MtbeJQ74g2
hQYjm9pD1+26urNYjWe1d17wOQChPwSuM/K76NLcH13NHizEigH4UJurydMroO7vgIy3SvczgA6N
EeDCnM7XeM7YBmDXPIzitetZ6gFkDXeJvaPqH0A7iVB86x0ZjAt7Tu3RPrJLx7ezA2Z2m8sz+Wzh
cr1yg8/NJuKxCHEniopLGG/S8pdF4yNc35MPEv1pZh6h0GpAGJHLpmRkwqnmF6PWgyeROGFz+vCn
aSGQxOGY0aj6/2lcXDTDVLIfauABzAiigV175btkpzQyyH8z1QB0Ja6zq2IgHkOhdCl+V0ygimVE
1lWsRKHntkFUF3MJ1PjPYjuvocvOY0Mw0B45IpmFb0rBaTct/KBtY7dSXBeu/F+rBMlCRV5rnBRM
oA/wnKcYeki/pUHZfyGAjQ9/5PEL73D4ebU95qRokHo+mXtHm7VFGjVmiQr6ka57vpp+IGSIAovT
XoliSuhb1DL+JDsf0OCTdgiMy0S5XgorXI+5YF3l0e906eHXZC6GNVtLr+bY4FgThOQEqtA+679l
xdVnVNF2X5F38RmrN2Yz4eczcvMz8zteKSYiIQA0Rna2Xhyz31DzA5J2RDRJBZC9docFD3Zl8Qbv
s5SfeiBpnbr7D3dL6nbIDvBwwGjRB998v05U+YgvVmm9GGyZv3d3khbdTlUggbizDzpAbZihbFxE
gTMkps+RcAFZLJdC+SGNvWDdKZ972idPqIa6Fi3EJY2tVn5wzhMr4xRUjTTqMZqE2xbbRjQT8tnV
DUrzVokbSD2AHjG08J3iso3/0wlwSxjXP/hrZxmp7xiWW6U3DCk9jZd/cfWJhgYifp53FPNXpI4U
fsbxOe2W0up38CuBlCQoMJDYY92IrlmD2N7gxlymHZNDT9DwM1skfooSTqOpNQsR8EZpU9FJvumk
OWnSptI+PF2esvXz9lMKOxkuh5BN6icueplTkcCfog4FJd5LAu7v7vQzq7erjgHcH9tkuoWeuXN9
RauOqCxJt0oSue17efOrDa33k+7IdM6/bxo9WvIQrtRUUodw7GiPSvnh74K7KBtXj4DXigh6sht3
hYXVZ2HCK9JuQOOuR/Ga6o87HV3y0qVEFSmTNEci8IasGmHGNVGDICX04N0DMQtP+qMJ82VjPOTJ
dJMYpnOJtcOIAM7zZ3PLh3Oa3cfERdkrmYSEd/QHeSvffV6skTTIb3CD+vLUnnX/5QR40qavLgHU
k4baLez1+3MIRQI9FL+9QGwxKNZp9qIdTS577PQAFYgNjmtLMuvIBt9FCSnIxGIYPTv4CwEFhAne
gWMDPVkDMcEzCyg30wkMEoJZYk012pXcywg/6OC/vxs3anhdKxUyUsxMS2fQh2GaUqRFNnUtDwOS
zeAdo9E/0/i6xr9e8Y5m/+IpkCctfn8ca+1qLWVn87JKdiRs1TpHxROa/6/7WZK+vCWXZMqmff4F
jCVW4sE8kgFA2OePEMos5JlVnVvtIwU18TWdZzxmkFmxQWP0dFt1/0Gwvb/Bs25a26Y1/ouwro54
PhFajg+GGWxm1AnSsaFdDNGzQp9g4mTaxj5e9vZHOlbEZm42kn0C5eTCWXPbOfCyy9c77oG86X7L
SWlppX/60qF57cAmmKjuEGyzEhjHYCLDyeKcXM/NtGfWB+pVuJWIwIuFOM3q2gNvYOgWWuec+dFI
vOqcfGqgtDllz2PCBsOmY3xb7HAOJ+AArOeSheaz9HrtFdpnd2pF1Dv9Xw/V5MM9Dmx3QW9kXE+m
L/KYK5vmEK0J1YcNXnyYS/vfIwPcxNZXnLZrKes97Kw0L/NmL4m4e0wTGkHF+SZKrzGzxWufg0yO
Jj7F3f33oSd4nTlpn1Cn/SMzzrei1HxaLIgB3MDgdQyMzA/PgT8YNLvFG57UIcGzZnUufCAbBtbI
nn878PDsjrn9d/mghnIhURGNnxELykLftRJzeL46vukZAkVZv32DpF6hFQhRAQF7al6uFCuhnujD
LLx/5ZQxrRXQsoZJ4Or5qLyMy7FHiD0O0aw8ruxDdHpbwn8n1YJvk+c17OxVj4LN0JGmQEVm7Z0U
W5wQmRZF1U21aY/uTQ/pJ2YsRHe16ncXx56YpgMvAPgcVgkxSIPZYmm9FMl3fy4iE6QNaRLD5AX5
97ARWliAt/4FU+SfK2DavdxeOsJnaDEmRH4pxt5bsCwaNV5lWCNdaogIs1BdzhZ5F+SVeY2diqvl
byrFY8Vc79fTT7sG5wA+k6eh2Ws3LYbsunosrBlzFx85PT0qYaA/xuKB0HhPkr21YEs+EkZe0o/w
ln2nCS85te5Ad4RSO6EQ5p5kEn4YXZRsQF4WsKvKH3+QVLpaxnnOBcHYkKmJY/WInjBTgjKlmwSP
sHlZl1mNna5IF/jv3L4fjYDXuSv24ju0TNsRmvjjgfc4MC8OUMWjStRhmgo81mvc2NqSYf0DeOT8
KvZmywTcxxexkOMzG5bpxsvukh8+5OgKPL9qX4qwcJVjhMReshM0Ypvsd+uDHKXa8m0v/Ne1fUPw
cWBLiF2Tx2iJAyRUxS1Wo8VgkOnW4F/upjYC7hiWr8NRZSaItnxQwaZM9FjMwFo2J3SpDznbOFXi
HBCPErPMGZ9h4Zr7YVnAxdRmiFzVNotZmWeWMwUStlw8p9fm7/a63USUOMAKUCiB6Zi2vJ33lJa3
/vsxVgNvqq4ly/RxULEsW6MvlMSBySHr5+0eIg5YsVW1jrBQNnVDihX6SB46VkyKvZuRiGanTAFJ
myFu4t7g6lLDA2M9CoPzHSIkIxknsSv5L8SVDkZexaJkjoC65Cl60uoP/YaYmvRGcGKpio0/sVZo
QhgMRvR/rSL/seOYlNCGuCjOGNwKXcg+t+Lv/3B5kDlveKA8N199uvvsOYo+ykUcMcYyXb3e+Q7b
RSgXN9u+8t52snI9LHWLvyV6laPwKkGPYXABFt7I1m5V4ToNLFOAs+Lw54v4IjGHMp2OkUcrivx9
y3FMsI5FggBvl/xVrIQ/hDAxBpYWt/iN85AEtHnkosXkuI/kfkydM8XyR5+QTuM6VEF5qvx/zt82
AeG9w2+8FRngkggwTUE5stUamQcLRSjlhvvmdj5+Y59l54gL+LoOMUcGaLo4Vufmu9UqQOJB2o8/
YpXlplHWW/WX80OOV+PNZ/sn7u2ClfH2QgYU/I1OHerHApKM0GWF7nVeygOB1Wp/+gWbJ1XjXbea
kek4UjUV1iSmAHH+sVfzaXS4p5F6ndg/6VQ1wj623qyYEEXLlRYxo2WQH1cTlCiKIh/svS+wpkPU
fCYPN/CR279EyvUUfuRXD0cGzDp3gD2uNepOBr6Zt4xihaZNnZhsF811W5OTlNI2fBR5QUQLWMeB
4IZgX+guxKfDKr73JjSpR0GOvfc3fBV1awM+glz1kEOQ1irvyIqG26pHCRou9M5IUlCKtXMVj1d7
b8FW6e9RD+jcXjwj/LvPFVSg5VpINyUj2QGSLigI6sXFwGrp8e4zxBYO0ZDiEurRlhOSJsus194d
jpL4lxsXmrCycah1xGNSq7JD1Ha2NXEf6O2IGHT5c/0gcgqUeOYrVHSz3ZKL8vJVp675Rm3je7cb
2HIg1rS77kAo62+ePnpgdSq1pJK8jp7LI7SefF4H6ht9bFzJgSZjuiDh6tJdL42iF3f7VisFDum9
vAf9YLcvixQl208wAvfhNUJXzdiVfObxeaIYvKAUdVIpm2LFvyKiTttlt8DWBRZdsGttMPelO/s3
mQ2RqdzqT7KYJwWRubsvcn6Cu3/8xaMKWJS+f3+KNVAjNAHp6M1ln6IUdUHFJR8CqheTwVXOuiuq
N4s+8gU08vZY9Sa1DdKPigYmhrF/sya6Cp7Gu7Ev9IqUYShCUGhmWdoBLwS6jFXhDUChm/zkc3sj
Ztiiga8PW025YRH6mxRKBP1RxywOVBAXmApxPiKKZ5l3NIFUFu86FXY36wEWSxdrMaJeQeQ+p7bn
q4mebdLr3Cq+440ywNva51qgFtsghONj8az+JTSA8YuC0LL03ehv3Vopp8CHdawzp3W5F9tB0sme
Xh9HwtviyaHtDapYhTAzpwhWxeom0JgsrG7iF8Q5wtmytfrXfewvbWTs/l4IaRzK052S4VDzad1C
aBKT+7s+99fa1NTgsbL/jFvLkVvSIEZddi7J2L+P48VO+kVxjVQwRbC/mQ9EwPHawNAmypxb3zwx
poNr/sQWjY44k5FhnBZTnzsOMUM8TKlwk6xW8fsJ0WdCOZ3uyh54xjJT6FUFZC1rUBgNto+fO/G4
CxOLYp8GCiG4YWpY0abWo6v2FVo7qRq2zrIFwN8gz1V9eLHbV0Upmv47i1uY+T7cKGV+sm4Mf5Xv
Uh3PHgxHCKPzTCfeEOR/yuU12d4pLZjn2Bc5CYnNWVEKzN9W+TUUlHsPmZTSU9Gs+pEVUUIDK7Ud
rIBSkA0IUpy7Gm44xTFhgNvmaokjKShwL1ZSoV+Dvx6I85r1xnylO0qWz8EaGVAp9AbEV4gkgzAe
PowafWz92aJ7kdJscvyFZhK5lxvefQp6i7UPAWEc86M46rr/F8dFTjVphgfww9ckh5Ae+49ue6Z4
QtEyNH5S+IgogOiLkdUPylwSJL17/NA5F75eOPBvElstAn+GZF9QcgG8RMIldCtzHxRXS9O7y/vd
D45wWzsJfYM0HbkS2Cdq/JFP5G5vEkd5dMFABTzMlq2OvH8SYIgq0k+ZW6/w9h/+x6x01zH93ldL
GfE9h6Z/BmcR7jA0FaxRSXc2cpblC/WVDwxAYFcYyLk/8SmSuQu2GiZlOEC6jwcOk7eqFb1RZDSW
6mjtsCL9Ees+ixxq6cR8sbLCVFxjCdeV7dld+XDVZva4L0X6Jr7R5ctODwpyqI+aRMq1DNAbqTdK
0x15aFEOKZrM9+/KDzJkR94V1bdNxHAPesinKJJ+8+myeJMzOFH0uFoZTg1znTiGDXbr2WfImQV3
IGpBph8r1YbvXza6/An0hn2U6InfyewIN00SjFRkfY2tU1cF3WOwwzxLdfXM/rnZru6UVUwMbI/V
eAB1oZNSroLsfr/E/ZhkoNGjjZjeMWQj+gt2a61nHc0Q6J91SaQz1jgbgEmJgwcf72Ivc29JDJ7L
F73FrxRZ6zwrKEGB4UtlQrmsMyC/rvoLwdK25Zp/laaLmbV+0VXt2Mx9bQTdpsJYVjDdg9IDuekh
qJDfszVVuW6cDObPLRLszkgr5rD/o1YCfdOVSFZXuY4+EWGbq1KnDIULLb1oZzheMOWScV9uWSOr
AVaFusH2iKXwJzUMfB5+goOL3hqQkFiFpUHfSTI53O8UxC2SN0zt/QFCmBM+iR3dQg+lGWwvWtzg
4qlXKjsE63ltWutDFI8FQkyx/PC9Xq4Xq0SKYxAd1iozzP1/69zblF7swXtcL7f2LSug5fArQTku
zuSsx+9nf0Q6YGhZNC5yIKGSFWNl/RNeOONdsQQTWMYpjsinE13bbPHsvwUZRzWWYYEEKP595Ws2
ildVQ4g2drvq+FMgNvzBlCAhjCx1lbNw5m9UzxIR2oZJUMXjElX9fxbDVPo426dvjKeCdtLtTmUF
lI9qKk8bXahieLrWAtI6HxgRsew7wti/NRAdiL1s/EyUrsu1Ld/e4uNrbrSrwo0Sbv7QGhh/rHMA
9RgSJbtHKtj06afLGlo0CB8no5uAtb7dBZC00pYkV15oLTxgJ+0AijjcGZWDECK0b+4MGOd2vt9Q
Y1eVRsRAN0OHECzDT5hs/vkxCmIHE6uCcigH23gkM/KXy1ErI4octtWIb3a+oPuULVKXmksqwvT/
hiN/g9kTDcqEI++qgdg4L6Wy452FePaE+1zCR6BijE/Il4vF7DlvYHfg3JTgIsNVQ9wSPcx+dwvb
6f25STbwNeDwkWhR/MmAb7qSVj8LH1BNBNQSvSljjlQUgup2nNvh8y0CPS+VzUj2BxiFeq7nS6N6
JzFfOFHhjlnih1QMz4z4qLCcWqTpHwDRPKChO3ebEbSyHDi+ecugTfsO4SBUQ6Kg6qK8sbidmC5P
X+eGLs8D5iamlNvZEfi48s5rEGTzd8EdvJ71gBM9JcAPhvaYdeZONpYcx6kCVYlNVKsTURdGReF6
tUNe4wx/pBarWfWbgEQdnpLLwjwqESr6/rxjYlYCjk4TqzhvqcPSRSU8Qo6jxrpRpuaTfXl0a0FA
O6XtybdfBLQJ85s3WGbdFZNgaSY58RARCpI+yOd+eGEgMuCQwW98lG55W6G7XxbyRoKnSu+1HNL0
StBu+mv5xrTPfrphdpkb9zVMLvCUCsgGftC3HmUzC341nc0NBBlaaz1zRb9OyDR2uZYPp6tZb03t
vE2cN5LVw1HIvHzS1vhNgpqLqxASfQG3LeKRX3cyDYJp+0ZJ6OwGe2gDKw40MWGBmgtpz8f22w38
UbqVa4peYfqdJ+RxmORmOYS43ji9O9tZCx8YuK0iw48AWD3Dtabvr2TX2OLOVAYz+4gucOuMjsa6
SMerowKky1RQ/pcXxM82QpLIkiK3Rw/BTiHiPuVYH8GOzsxETne3mFqVOrCUiryf+j9M2g7QVxhR
5sAoliyPDsTXq0ZU0Oj+wtQceESqVWsAwxmTdcf/Lypb8WLez5vVqJoeDeXo8xK+wk6zbzO6GIX6
ladeKbXul6iYa25cR/vWibQ9sNUs0KiUNbBoN4BVVeu0r9cEyAVWHtBuonUJ9npZRWPuLA35sp+r
UMXcV0OYV9n07drbSQYi+TZRp8cGOVTVOWC9V+UkesL/bMq40uWGR63s9kqyfgcdSYCAV/H5Yeo5
ichGtkk3CIYul/a8RC/IxaN5iVLueOvSfqZDXJzlh/vRJ/xV2RHIHeL36lE5Ix3S0dQeELDpxsHq
vh7c72xnhKRMvO1HyCtO3iJDZzCIGXO6pwz7V1DDiMoJLUc6gL7QZRppCxNloDLHNm7MQMjBsGT9
15BSTF6jCpS1ZQmeCI7RY88xv18+Mx3j7e41avY4Y0yhy2A5nP1WaLLFZU7LW3BBd4W5e+crPR5+
gm+yt3QBeqZnYOz+L0yMPfX/XaAmtRvrJG++yRPJEryVk37itFam2rI7n4T0FVS529fxCsfy8n5h
J3UA382JCm9IgiMbsum564fepJ8xdwziSaahYbKex4LdZ2XR8vQ+9E44Adnv0s1IyItKqNJWdx7I
SeuUXuR+1E2oE2G1LoUyo61UvshUglslxu+fTt/XFu8Le5w24Q4EXm8FTONoqCw/nDpeBiwne+S3
VSVtBnwW3JBaPLQ+lUc8YcOwtM2D0scP4RwpUB17PxYOcwnFSt82SsNM0kpTpWoYX/dARX1GrRsy
EjTWYgH8Nkg+h49xoOBlvw6j1xD12SQ+Kno/gGcq/mJbB1ayy/hIbempNrBi2Tn5+90keY3uCmqC
eR9d2GF9OwH1iJddUj8Ogq2uSbudu3bDI7Wf/o9IQHEUivVRM1zRN0xhlixRd55zHPeVLRwrmnJP
69+9R3WGzgSIGCDhOLEzoF9o/RXQdsfQ+XRtOAJGtEBfhPwCV7FETOwllKoMcfnOfbWB3sXai7aV
kvnZf6iVRmSkr9dWW14QNVjc+klrAOWqfPqEaDZqsnvhilypxkmCwHFadWh1bXK7aq2in826JaXT
KrB400uAZHz/mKgrUBLlJFS1fmz8AVzActIwQUulKnCikZXoVjf9P7TYI+d2uz1vwHiFvmaztcIN
LRztoQG2oZXmdI1m7TtfPdsO79spss2li0mtwSRD7hPsgUgJdgidDF8/me4YkHEYPqejiVXUpgGU
n3SBUE0LA0d1IBMrA0ksGP/vKetoPvX1v5sp4M160dRyHKxGLWyLlASTgT86P7NeSufMTASbGJs+
wO05TLEVKbRSgIEBuiRqXJ6d18sCghwUyPA8BjVsi0E4ffzd0WTN1qoHTDN9cnbuiVEQPAgCjOWO
oySMBdaclOvEr8w2M1tNV5N/HTCkHZsY0l78Kb/MtwWIQfCSVg11J/kRwc2NoSEuh81laTnRE41a
uh3VpX+8mhFyvnQvHEkDqjSWToFz2ieUyq47312QyRxXBaib84TJak87VroPdy3UeFu5CD0Zbxkt
Qy9teZxC9hS0GE2zkOtuIDLe5Yf7pefaOeJ8mEk2EhT3AsdaqoNrmssc1E6Rj8ecyc8qhfeOVKox
gylt1I7zatFkou5ZMECRJcj8vwDtL7lGhRnj1lqXrrXJySpEd4/vTRppcRa1tRh1WRdX4ChD4rHO
S2eNHCEOyY9t/eSIHMHyzwHV7fVBnUGp6swfTk/gBbW1CwgBdyFWuYQK+1hbYkOWkBX9ZNOfw/55
CCMBZqe4M5Q2BU8ORkz2c7bTPROvfOYSj83x4TLn/rxP194u0LxEZXoLeNaM63fQkKwXOg5GmBLd
zx4V5Sldj7xbTDIuRmfacvNfmmLhjvTQkBnEZYh5EtZi6nf4m/GAISBBNJe9SFB5iz+z+DSO7g3v
kAO3snuxhbn4qfeIYcNCSLsLARHlT9of0uMcqPbp9r4WjUq2wWaDr7pasCd5hAcAWwPf8lbSbRv3
m/Pteurh8FSCGM/03YEb1Unoh+fZKdfr6E2mk2zAdTN6TJbhgqkqi/I3OkReIB1fgv0Og4GkrGSM
yEKUSSkpx065qEFnkMmzJTT968qZLtryI1grvuTQxCmkk/aGCrrXAsL/1UfZlIVH3T0CtJE8N6b2
lpWH/UyFfq1v5/YIfch+8CHpCEWcuW97d3fRNS9xAJf0P/qtRoUnm5UYq3LBIr/JFQAXlDclq2Uh
FGVv2eMXYOzWS9EFADuToIWc1+c0/ZD5SQyq94el2B6S51UqP9634maPUyYlctcWTpGet7eXdPZw
AAiwUsQZDaIC8IC8RHNuOvq1TM6SJCBfPrrFqaNnIUA4OW+hZzlFipzEslz6+uK6C+IW5vXCv43D
4BpYDLA7hVvZzdus7h7wTTSdir7ZJ2vzTW2cOzLCKTcPmLkqZ0mqGKpmYjk/juwctk+ydYeyGqZG
B9AZYvpdS1/aSOvm3pSfUC+ovRUPuQrs4sopc4kgVDyLJanHIdiGUQfg0efA32hVNuY4FfueW576
9lJvLIdzduF9p8pBoQdMmkYdRYY1PfIzTl+LAz3Pu4wULURDM2TjiulbGJdvY6Xm4ptGQTQEXGOp
44UHdGxvH9ptTJbA7gtxJvvnGTDBfucPhtjQevTxEbo8LZQOVjvJS66++qG7ybCpq8KE7uzBruy/
HoT9opCE0beWz0V5SJelgZlcg1Q4otNZwTU9Lg3jxope7iSjkacL/hUWEcLOsMszTTMvx8galxjJ
Yz9jU3gEN6swibSA/NoP1M1jqPPs41to/yih4J7Zq2jh/JK29/oFkGiWvRVGDf+n3QCF5qW3DYMx
0aGGmmAV95U7IJPSeZEgkV7g+EioXjfphGjfdXjvWn4gyo074be1XTI1Vdf5CkF3Q6igBlGi9v5B
xXaawNydk4IZ3QOpiw1OwyO6PzIc+fIkIczirIlY7017WZhYMpgYy68I2llnUhgY15/0w+4ObbbK
rjbg2HlOgqMwJQlcG5idzm652cztQJQM0LmDFIgVnfDYnLdTMySGHK9HT8nnrL5uO87Pog3Dr+Xe
w34TWHu79Spu0LWLXwIF0Q1dwLARoMzhPGZojovC+tSxtx6/fOSYjDVsSPUvI+5VULXjjiz89cal
bHsUBZQHHI/v5z/uYBJvVgTksyjx4cra82rkQxTgyVsSBo2O38w68SNkjuytyvHQykLnq7yzJpD2
8GdUyF+klINHqCzct7AM8CDqC5qDJNYWX7GcOi7sdngeIs7AjtndmL1deYJX6rdx/UCkw+HaLVk6
LRU8npq4gMksfHMErnk/K2HIyEy9+iYTro4FN0R7J8r6HW3DniEgzcVCF9avBEWgRZjSLM6gxrXW
oJAbSIUEUbI/8eQ23ufglgc9OTewU9GeY+i/thvGH27JG67H9RfXEYqh27Cmk1QHSpHzk8RRdbQG
mUu6KzqvM+SDyhDlb+HOL2YiS7v46c0tSkl1k78oH4WXoHqhP1GrjRmsQdBHw0x9AQmYTBtq9sqL
T1z2y+YLYWGEWze4C9kwDDbnbJ8llSwuvkedXpz5o7sDUjSwQwD/Doeo5qZcNlMVEczu5z0d5XvR
rkPw/vQ4wNGk10/yopYeSI/R016RwFWQS9r6wrW3EWb0sKqP7TGlMefUTK1r5ltlRq9FYQA1XUwY
tO5soQhBon9tASDQxM1kV62IO+c0iXUv+AnfRuAFsYc8ucUFz8ZZjFl9lbUHmBIvOTHjQ7tDag34
i8A6ybzGHM4E4TX5dXfkYwO/JQ5QDdXQ6Q3hwKhC5ZvDLIbSI8WcURES9xa8VPmko8M4UA/bKMdP
Pr4nPa/TcgqQVMCU7pDfV2GY67s/nI1XOJ0DtOZ4E8o9g/6Kjj+ZDh3gf2xC5UE1NMrkPD+afJW1
F+pp2h9Xbtw+2reggAzmTvgvHUOV7xqunt3onzJpuLEC2cFiWE2J0Il6E23YrAbSXM4yqaHDNhrH
JXgaOAX8aemReTJHLqwlXvQjvkgM/HaAu84kGbSa7XSJ+N0/pF2UNQi3eroC0uRkRFVuFh6KQq9v
lqAz8zZdl781+77uzmiP4h+eG4xejyTrsOAWjV2XGlq1lWrgS4QQm3HCR57BnesOO1xWsTrYH0eu
Q6G/n40wKd7yDwud9K2iZ86nVYg9IPA9QLQAGy9x8uiSDaRKX9TJGUIHfHQT1gqxMW8IcdGK63fr
ttQXvThGgVEAcBP3l7a1nqI3L7Vf/Vn8afkruucoCt8u4PY3CsAAfJnMXuHvxh+ecBkcOfQv1ooy
Ul93Dm1PpYp5PUNrPgGkfm+0/U7YkoCIS7i0w4Siu5qOOnOJDpIq2+TSf6aZ12xcjrn108WeqXid
j0f2SKMUBX7Mpq0mapvbDDyvnMW9+nb+xRHGBS0t+jhs2Zfa83joo3QdpDhpnTIu/ecdRhOaseRF
iW88XN2d6BIOt/9L5GTtU5j9UCgBD2LJRv4gpFuAimeK0UGOPZhlJsFNK72RQafcmFFm8eF+/pXi
2pEp9pVrR8HWkoX6ohgSVaSVo5Dy3q/Jx656QdljKXlBFfCXWYRUWMQzXIWGTD1KMRN2+qL2WfPR
jMdDi8+4c41ze6xuDiPsPSYzalJ6Vf4zirXMYwcP127ZTfopE9PGBsD0YqS1vi5PeQHOYMBgtIOs
SQcfp3AKfXLmSRaKo+npckziSCZyw3TDYpJFCQ6vfTpyNFaxQgozJnsSW0BuVL9TitaHK3OH8xqV
heHgnVavAepJn/cYQ6q/xnJFob73fnblEK+IH3cC7rULVn8Mr1SKpQYN2VDdOp5gGs5BVB5v6Si1
n9zrdQPR+D/yC4arA1SW52bIhFuiTURZ030ESb44zx8C05/WGT/Tre+otryx3VOyN3TcqiGpJqlA
DtOjjBmDbPODvj4leGJ9/b6uebfVheueNcv1ghvGRGcK3CwioZph5BlxCt7iIwHUdqxRFR1CSwX3
m5AyFIrxgCeJDBbNiQXQGvCtuddH833YHIoTb+BmBeB0vMbMBexbSeY0XbolF0eBbkC1LbT6eM3M
yb/T3l8nITnHuMjPzxPCcIERJPg0Jo4EoxRUo9wiarzdGoUu78f7OGyPEO5j3YI36jlsvkGAZC+t
9aQfjz9nDrBp7TRj3E+xMIFDeoQeiUF/F/AGiZ2MCN9hI33q3q8zyold058xBdEJrelM924ytN+h
C3MWv8DB8gIUOpDIeFWAsbGjC25PZGiXnardSOwDlotd3cEOvr+0QDW5M2R+QCvd9O55DvsJkGZ8
s6oX7J69XeDhh4yJZMUsFSD0TRa9J0ZdCkvgzpK0hyZSkTML94Q16YAVJ1kz+xtnmZxsu/bc3tdD
+WNlTo2AKO6djThLzUoOGh3MCcI2ogL7Zv+PEEV5BjPCXxFRcfrPdFved978WIbu/mI3RIPK86XH
734oNyHwBa3Uoo/liZzdMTIjJKKobunibk4Jfuc7TmiCEHdu02pReiEGZhRtwRe731BiNtobIefo
5tXkxDznIY3i3QQeZMQnnQEkcp4Hvh34S0KGroIjvCe7Qpn4iiJZ7uhGV9TiRUAouKtUg0PoF2w3
Ev2w9aPRb5R0zX7yUC0l/DhiOlRGBIYXPfG8zMJTt6Oca4gZLwxF5WAXi7B0fb5TcofaQ5AP5LOs
hYg4nTeg+wCRlBJ8SaIxtXOFL+Y6sNI8MqDfgq8m1C6ATrjJt58870bTsMelkn1S/vYFRTbNKhy6
3aP5fvlFXykxwFTNnmRJVWacU/HjL/YPw+DJ3mrwoSKEIbmUu6/Zp/mvA1mpocqk7Mj5cBU/xM47
AOE07OJTlq7ANWo5cj4rhdxbH5L9zd2KlTyVZ9LVSxakdfNgb/N1sOc1eKrSAJmsrJntGjg9yw96
6K5SsiYBEtwJ2H8oMmBQ0aTynTrR5VfDHTaFNPIdTsyhfFc5rjKnUMlBh7iIdCyRzeaV21R/kBFL
Wc7vcsbMSxq1BeckW2np6yEbraa0JYu2NkEg294Is3xPp/U0rbH7yK/OtjZc6beemEbWv7QaZUwS
IXeBcwqZG+U+VzcGuRCMXD+4j1i8DOof5JMDkutzt4SbHz96ulbZyuU+fnDZeOmou7/PeGmLZ5kY
6CuENvJnZpnn9fTFvOWTq/dJTspu2uZMA4ea7aK7ythf9XGiSn84IrDpKQwjH5JyMPSR+qhLvvEY
j2sybL+y0FPM/3+u3tlqXR4OKammCdOUd9jBLXUJurlbTPDWfHmaQrQKlNyc4dFB9ilkPLoOhMmv
jyBiKgG305oq2t7y1XhPecSij2oC0weHatooTyLXgDmuslEUqP0xk5cRjmCTSyvuS6OUYqKUVGst
peT5hL4Rs8Z71VnsybhpOFjoHqOv2TAa3kJdC2tDhc1qFTmx5hIAi8yjQ9YCVjIm0MR3Yx4y8ZeI
vwvVRyi2Jq6CcZiElonImMmSNQdFf7GYZq0n/1HML1r8iRD0homgTP2fTup/UOJfAOOB7eRkwkd8
BDjSkHTM+tXlGMXLvZ0lL4em5IUucNO1MmeYYG1NeVkrNKppq/HJu5v7PDi4xZPjiGlYwnZ0Uzp6
cB2vJK+WaOmZu2h+MvLK/ThTektgMm5599JrSuvBKCw6lfoLbouqIyq1kugwbdWKDInclomstGil
4Q/5mY0TtQkPR/QhPD01iB6HY2ocS4wv7W/1SqgK8+sZPJcy6sFX/4eATiWCm9T7TFjGlFRMON7x
KiBVdLnnY+Xo2vI5rehkvzizmXV55vLo9eqN5dUJ+vShwfGPXVj8ODvz97HPY3QSn/t98mE4bh8s
XGHmr3S0uXh/RyYafMd2W5uvOw1lt9CZD773FDeQAjYBZcB6AnxRgPde7s3pe6MTqBcbtizbwWaw
Iyk5bkWXtDYitpa3S+2cR4khTgERO61JyQ0v/NGDo6M7Pf/AvFWYxmRdSY2jHpZLkCR8qGcIs38V
6t2wPGrLiN6RtbbCUJzMPbzovicubG0uuqdLe7Eb8RMfakKjZb3cSAWpIB4MAk+ZXWnmRmt6Ogxi
0vH5vUb5uGKeuijsbzIwvMa4ouUKn2XJjapZ6HG3u/hqPJGUy4WMShw8cJmcv3VY2mIjuGuKzX3l
e8HqOe0ueVoI4b11+XvAgWWUsZ9kKm/GopYM1A1VbVDptmN16fdamHtNJNDr7YlHppolw0tdix26
TzphLnlWb6ohirkKwcFsZVElvzO2Rzpi4yT4rolHsTy4fH/PmUTGUAEq15FZlET/tUZy1BxF9q84
d/LeBaJhPo1XlTzqk4eedGOsLG0URCyefb/KQmjmPTrtJ4MnEceETym9tjgz6AcOkpt8+3XV8OtM
yRB3JNlsYzMGE5AjBtqPtY5JTpBL1qUGnJGssoDYHbPfxhB+18vJjWofLCMpwLLRHOAt/i95RTwI
s3KcKrB0Ci0RTK1ADZzV9GAGAc2Ps1tg3Srp8JLudXURb3TUcNG0ND6z+GGE0Qjlm4zP/DO6RUNS
P/ohv/XU5EYsn+NY9amdtcFmD9WIVB9eheZUtOR8OeLtb38VR/ZmqtfkM345XdzbIjgYmi/ZzVeK
NtD874DZ5Z5zvvX0HYnyKSgiU6F9gEriSZUk+8+UgzPokY+/+0JOdJvizbfRk5hwWPb7DiRzcQKn
vKvYb1vUYQ0+w2I9FF9QkqTLvpnYsTBCprBGMijIAwm1Oa+Tl+8RELAvq+Rglgsh77Z0IrcfpMs+
Zqltpzphi7rWnX0gaysIOIk96+T/1bEP4cLHejeypuiLFhUy4+ZGj4uKSNUJflLIO1SlW8lmkWfM
xDHHB6P47md9Wz6fFn3esgXKChpo5bon4g3z9Rdwnv2w9A+5sCZ6Dg5CqC0ERc3UjJRziMRr8Td0
ZnuNGFNgR3WYMkHXm36AV6aMJsZb7iTQ8fcLor8EQ7pvyXFb0R/OBswHGwDiJYNvV/WizZ3YoIXR
gjKnAW5s8a6wQkNWiSF4p8bFP4+Lzduv6jRYnWUBNTsmO2NkO0QEyWzCMO7jgjzM7HFBk0Sb8wxc
8nIsebXZU0oxDTudTbHdj1sSp3S9oVMa6yg29Qc/vfSbdlMwAWR69nkP+AKr7WOwUrWvbKS97TMC
9r3BbtvjFTxXJrunM9ZujZYbH0yWw7cONBW/k7mzfTx4jp+CHlXXU/zIPHtC2z+PFe+y3uguNLF7
jKXRw5+IoUZt02uqfWKq7e5u8aCeGko8uzMK01RQh6jJE3iiuKlHuBnzLGQBaEIZM5lvzP87mj14
Hmcpw/dv4JKfdgdW2JdT9R7ML2DzoD7j5ViPZOMXb060Ow4GmMzpg97EwhE8QLRNGItVTnoHWbCh
0s41L2d9XG1SMnQXW8kwYymt35uYBvFmxr/4yHLmMufEM0xaxHEhBGbsTTvc/K8jsrncom1/YZ0G
5rhUL0qHD4OIOJxhh1StfMHM5LrEwMhgKmAUztdVu31N4JPI264XFfEzeuNBJpx1QdnEFqn7wVQh
gmsfNuogz5fJ0j5ujco66sVAUuD7lY8rNrBIUMLnk1O74KBBtPV1YtrGSvUPphtaXVut5SBvfFwj
pOTK4pXNT3XhB9ayixCLFA0prezoog0aeij1re7V1z9QdAifSSSvYlaXoYWM9Ve747TxtpaL7785
fHqN7vo++5EcgBivI9eRA6lc4lywnydFh/rIw8/uXFyzuorZPhMuD+gBtw0bq+NeZAmc0FDti4kI
PDgP3xoK35bBHKJD7nnrD98DA4iDZzO4CridEMaH2nB8VjbeWs4+d67bp776UBjkq5DLgNLNd58B
iM460nyFDEEjIv+yNAIsqERijyRMzNamuIA7MlcTJ133RshbDHMx10n9YNDyo4Gz9Rj3Ytr18PV6
XM7zdNl60bsWuB+4A/DG93JYpudFWAeP8bT6zqFKcGsGRgEBf3WPkFaaYyXfRJ5qj7q3Y3LXiPD5
J4tGsPpvF/CCorIQyGO3/BKueSs0HWqZXvQAghcG0wyq5Qg6o5D3zd4ObyXOrexLUX535gZR33AT
8K5ysEHIVbHmDjmPQIvPpsJEcHTV5YoM+Tv2bDxKqyff6IX3sIvXONomld4FR7J+kp5GQeRpp+SA
GEqJpKdQyV8x1oDnCV7c+Nw059Pvs+XhBdFsI97rO2ABRHpZjOZkdJgPecLcF2lnuKJssH1mLlMp
ChzFpKm7BnRLsou6/A+P4HHwwF9stBpphpj2iMC3vArINnB47gPbAYJvTdiIcn5Is6ltFa1/bXUN
F+Cn0VxcXSqERWJokbx7tgNR25ZDy3QObTH5aeQAqDllIWXLula4tPIO4kjHZcQjRef+tHqgbDwr
Or1gxmm0+1PSRCdz2EG0oB8gDnjrpGacX4ouXrtPUeAJgke7gryCdefoNXFuL1Sk/kTOdKeX4yyW
4rosoDYbc5MirZD1/5KjLN9SEpogFhQDd8BLAdIUlwCFjZRUS7wR4dxDUBlrTxZtzpZiJ+m63t92
lfPfmvJsbz7dbkjpnD9yhOf70HP+t45lgEldYGe49vZp1MbEJx8WfHb9NNmUyl6uRrSxtnQsVl4x
1AI5+2/hPt2cAAAmRi8eInHu1oiX7jISp1sDyXH6j8ZcjvZUAi1L00XoYWaMZwSPOmiVuNZeBmXY
dL2TEU8tf/eTkZFfNMXLM7IUlF46uS6iio4pINSti8NQn2pNACUSnGUfTqLNNI/i347M73jvyQqK
F14GLM0Vh/6GYnqDDCcx9+mjakC/MjnFHjsA3Lw25x2oiOfa/KoMgh8LYr0839bPLT9mVJgnwqgi
PxxxUM6tSVV8LOu8huMHifb6N9vJRptgvsmPw9g4oSnhlYsIq3N1bsOGs2HbN4p2htgvyhwyjC0H
AyEtBDLCJwcOkIZj4fjhOToLgfjy5R/uoVMxQwmPivW/AFeloUk0+Gkv7WMAjqHIGb88o2PXeySS
nVgX7xcmPGdWeUx7gxUjc1lYQ1vrtu4pEK1HQj9i808VP5GLPhivSJxi3ZkGOCFl/qOpI1YMVE4o
xrfMmbUR4o0YYXgzBwIX/Ua7sarYFyaeLfMXiMdU2XndlVS68ODa1UO6Omq6Huymv9KEyFsA1FPu
9RxrHi2j0vXrQZ113jaZNox346XoumSFDDeHhlmuOdUqTUWUC6GFRMKw1l+WKWNIi9YJjWERLMU0
uNFyNPs1u8rDJXNE8rH8HZ6S0wiIoicFVZCnJs3VCOGujUYePLK0N68k8IxdjEgskcKJMs6XEQPx
aN+4wMWZiQDQAO3FnZr41LminOkLNvYj3+ySoBrby/hjvQiG7+hIcBTC/dLAoz+jRKOQoA5g4DKY
pSWD/E9QU696u1e5D38L1IWdinA/d/Fhr3+SJl/rneJft//yn4WnQmo7K8XZGudPII2CWj5u17wb
BdM3GEC4wFWJlCC4n9elDOYSTU1KdS71VQukyEB75kT55GuIEKYZ2TQSc9ap723Uwg6TVjMaRp+T
YNQO23wX3lOEaBSmGuqEniYO/yJkrL8q/AXHcFCmFXde7gyiAUYAYEzGtGXBdOh9XpTq8iCDltqM
hnVEjbpjEM9GqhizqJDsrCn/xx8k48GJDt+QLJhtHonCw2OHsrTbc7YRbOc4B4XSEXHHFArh49qF
+LX0uPhjAF26D52jKQJj/a0PKcbB/PK69UQ22To9F9PYja922IplpxswPsTotsb8g4TDaagvB+tQ
JzzZISteiBAj6isplEP3MHQJcQmsL1L7LzxGPb8lk75gr05UZ5Dzb3R8U754tJhndRNEvFaWdKdx
Kqcn/cU/A6/6OAJBYer1UGYjE+wVONUcPPQjEiYydTlF3C6CIMaHzR3Rdm/TXImSW/CFDU3olQHX
+59XM366bHbAFGZF12DwkG6fpzqz13K6BmioKQCSR/ydmrFNDAYlAQq8jYuWryDC7fUGAmJ1OHXr
N8P3CQ9sOWk/83S/+Y25jhhnruA/II5yX9DjJQ/VugMhrdTtTpJVGk0pRD8vEBUt0wcUvSeimNTy
Oj11itAuswwxYNHGnHRnoh86qYHyx9zv6WpHoc78iSBSkm3LQD6XsOoKq3lfjz8OO5zVvvDbcKWz
R9yfAemHEiN1DaaeeX6Y9EoyhmUbnRYGvdRaIdtJKXTT38l1CA1sRtrYCDpbaJeVFs/tTODnMFZT
s/9qs/if+Jdb8Y1GST0li50y2IHb5oiHvV9urFcLqw46n7mc83G4Uz54Gqt9QuKXeN/qQrfGCJsr
0F/nGlj511lGOnCHbdUEF7XIdOcjBb5+TxP8uZu+YN7SklcFd3jCV6LnUipr9M2jqAwYcKHiiAmg
/f3pAEcn7qyMsfrXAW8TAaJJeXu1I6OQr9jBqjKtEZcLa8iMIOKfSn5cekKdTY75nu1uCnosNrvj
2nn5E6N7dI3x2AzIwCgPl8NYdrnvREMJ9RQfjLtihbmO/4KDT/wSPK4HsIYvQetMlpVj51TL1+uy
GyGvhrRzO1BG/Egi6osggAld+Y3tRAEf5x2KsHNKMoR7KcyrOeqMf/HLNe6hIc7qziT7rlwJaB0b
MaIQu7vHB33cYhJcCbH2KgBxozEdZBCkuXxOJePRDchtCy6joEzEcMWRxy+Z8H6d/VsYulRHtfQs
rMUaoZZq9ZvGKcbXn8lkcTvVw4m7vITKOufJW4dBmNwX4SgUUNbMLCV9uvh15EJmaZDcdQPKauNf
Wl5rnRfgtBvtOgjJpeiOHvjB7hziXlcz/hEsdJV/Hti4WNt+C8q9nwMTzOEqUHa2ndAq7v64RzrT
F4fi3T91UU/WJD9GA9NLoMt6ve80Mxn0QkNAQ5m8qEx7b6aaRkuVfEcQq1FGx4uwkAKnLcQFH3oJ
anATO8YstWDuP6/mdVwyyGymb+mMLVPHOjskxfU5tqLK1XfHhiG7nete8aEZ9xl4i8fAL4FJ3ygg
Bl3WO/EoTTUqZ8IAm/FIt79DVh6FsITX+Ai6Wne/G29HZfpWgNnk0zA5fMCsa0OFnrKV5B0os4vr
WIE6thgru9ORUfMQGbuTPvhCy7bMSkXVktvuqCdohUwI9lUhf08mFKXm4fRooZYaGhG6Yl+psUe+
hNv+VmHdnjWUqtNxQW2lvV5UXrsGb/j7LtQUG94gAaVo1Pjz60TfewAIb8DmSn0wjpjjZAaAGpi3
d0XaP/sIIfoCYDKbbRrA2s0rM3La/YNfnjQOd9SnvhYijTDGlcsD5NXM9qdrVhfiN600JVrsL8Po
Meqy8qKLlo73K8gj0Ww3mVsnwpCQbW4nUUWOBxo+eRsuzvtra345brKrSfd1a0YQP+3pec4/QcJw
wOGGIGYDehRFSW6OI7YhkCpbYaKfg1nzczzWYpIua7H+QUtifPxrKlM8uTSU7rGiI84OBQV6gZ3h
hQCHaih62+Fbt33EHyeTfY8jNApmQSWL9YDjrjXQF5hdVRYuTd+FZDZTtn7/DSGj/OcQ9nIzXZnE
UxwTr+y/YnTEpQlB7nMe306or5hd5HEzj0hR3z+liavz4mE0N6d7sTrEWFnA8LBg7H4pGm6f3CRO
+Lcmb8Gf1ZXulRkxbWc7fWdYDb/TknBYzybbm36gBtGN0dpUocd2N/5yeO9mFLWEgB8qh/H7g8uM
mT0lf19xk6pGhsQPfFOeElO0ZEsL7tCTFintGrUNB7K1FmwATRXU1vSMZrqflXSC/cL2bULYfScn
ZmQ2YikiJbyBSNufQvA+FlXZLOflpvh72kUg7LhJLkfFnBYUN9FiaqUclkOWr3Yuos77Lzyg4M52
wxscyUn9Wklc2k7yXM9TwAauFDFCeTlbFEsImRmZQFvobNwbYoiLqF/7ZZe7WZzrBuuPwD8SdVrQ
WgJ8KpSJMxAU9M3dsyXZH341eaJgts47OfmPSvabKBtUcjnaQZ6eNdo7VAwAwWy7Qxu6RLsU3frV
LTc6xw0BViWPl9Vk56ixqLAlQFMqj25HzYHTmzVWpVjJm29MSjRbdN2Yln0ekzjUDz5pOEvBwXhU
EIixnvU+VlT1m4/I6ijhaPqPGVnlnLVwv/h9MrCPxB2QDWxUfr8RxieOTop5e/Fx+lPd8LHf5wd5
3Oc6qq1AL7uJMUBOu/HmYfp4zXggB/UkGTo2CgIrjF0N1Ck/er0MXv+BhZsy0QEQcMbz5aNdhj1O
UoeMtxYs+4Z0xxfp5sd10lGy253IPLV8+Qc7JTazEbOEUMwWlSzbXRACdJnrGM7Ayy6N/cWwEGvO
TFaJXQva8OmbVq4kzk70QkliGLFH0nqoWyhHpEeTjPov+IZzs3puMX8Wc07qTSzmF46XGZ89mJ/n
ohWNozY2rvIijwvHpa8WoSZOOb6EyiNEEuTc4P7/mTSu4CYomIfFgzcB45FA+Fl9lSRrRHQXI2q+
ABeYGRGqryBNz2DqAQGkb7QIzivpcxA0aQXj3DpYUk17G6nMKD6Abk2SmqlDpOjXVPvIDiGTABWu
LOMMCdMoFb+eCrYso54bP8l2qkq63hDAx7Y/peZh4IYQOEwtXHnbTiOUkMvSYSi1p2tmn3GcWCjQ
rup/BLUwxWWLGF2fqVAC4vbli3JFIu6uz1ZR8TiSYcUk0Nt6S2Rt1WFRo6e/KXjfupo6wJfeWMBx
66Q08C0PJyXRroP2fZyXCIZ9eUZrl7/uTC3tGWoW+rI/8ePuVh7haS5pCaHejgwJeoCEiJLNlusL
qeHLyx3lGJjxg3PrszrQhXApdCXvsrvX+Tx0tB2U5as165zA3zhAURNfW3f8J82eg5mniEzGHi6x
pdlKFqA+E47uJEP7VmQKFn1IUHfUbrbawkJunlhBRnyyg2BV0sxC6QqXRfvEZcdyCDQvNAbSrLQw
Lz5CSi6j5T85Wg4mGijuNeUkpZIx0DLJMbNCEcnYfSBYhY/6p0RYg3oJPWnotJ/z7IZo4tbi+BSu
cbngWs0jVbO3Lgsz+1j8T+mvI5q4wJyp2Ajub/snhMFThhsKiLzwXnkzMAs4W2psYYaD0HAVvO7q
8DhdbOe1KTbWscfgf2Dc2raDPqbROChBtFA9eF4RVoaMlim8uMLDPyFux18xIC78mBZ9CWi3pygU
kN5T23A6ACMEpu2dhyO+F7zZm8kOkbx3V28RjXVQgU5+IflET64ULBXUhqcvUd+8Q2yk4OWUkLeY
fKUoZWQNNpZZ9nIijYf8iFYOiXpaVSz0di2/6SW06zpDKvfb6+DTn8vML/ua3vIhtzDwROH+KURK
88PTLp87a0upf7DY/5xxbkCPMxYtw4hPc5PlnqYhjafl91BuhBT+fL7U4Y31BS7nU5skrmxcFqif
N+l/1NbybFrN0NESvGxUL1zvXqEdaQ2CsGWnAurGkDNY2HYQ69YcK3sgz8E8ezuGK7s2wUPitMFc
KNWNFSSVUGluvldUL0xlNeDDYDPB5RfMFd35xSEtaGOQIiM37jNqZaPufsht+oM30IyU6UYKKf4c
vr3nVisCtcEQz57go3QF6hrkLxjfjNjBd2AIzJX/IqQUFIjmr2Lr+y2V6vBGOt0nWAaeCtFTP+2s
OmA0moHS2TedQlFIp8DQ/TiJOYWP6NecZm5oFid4E+UIJpD48QQrlgR5UOxzLHArCUGkQVJLLJgb
iyrXHRXdnMnj0AmKeQbhhn7dtwP1FsSKkMuUiWoOmC3xtkHRtf9Ns7xOGvOtTnkshee/Fuvm2Alv
+Nmhke0twJCr9CWRJghRDKNR4nomctC27xwHzSMFIkKBj1i4s9WU0Y0seTQoYU0z8EBFNRcENl5p
KNSB6hYtozTQZ8FpSZFg3C3erv1wGTLWq/Jexhi1UEUKaBaKC0uvwU8rUBHKzxIt1OrBsYVU/gv9
iJYy/NX8qVydpFI9E8ac/iS5A4Ug95wDqVhsUymYwV6xgnBOlZR0y0SoBO7kfVmt2q1Zpmfhk62p
UaZZQGR3Js8GzBNjlnBVL+UDiurzh+B/TxKYQQ94u06zUEwoiU3pHWlf/Bye0vfMJhOaTO/E2VlP
5b0iRwp4DhtErOdXBWpJH5Nci9j6FodQAMNBeQaLiJyUZShWE0k0G+n8+1zAmcfO64O2W3uwWHFO
121qcElbJfO2V/J/cTwxWmFbfpe1bIaBczXVnv5i1degnASOzsftqBhH+iLlRnOk6s43YHxGLZwg
DBRig6HGiBr3DnoKuW7HPX9AYfP4bB4yX+GVIU6JhWeadj2r5nlKvIAgTuBHfsdtlybd6qvYfIDi
qGpX/C8byyExXGkV+oAgp9rUksQuXVTFjhHNijDI4u1g5rc7aWUQNwVUQPZ9VCBwooWLBsj0hOcU
uSS33aaLfztH+R5jB8RtSloo5HOugrmuATHqE+zXqyPe9jj/Pwzu0rqiNMBo45fEJu++i8LZ2ZPO
5Lhv8FjIzjWhbrFworKyY29MJY/oHxTKibq9r3J9zEaUQFEUp31CgPAer46qnYHzvG+eUncrWKo7
x0PPm709uiCVabPeLJIqDs/VAHugXtF49tCaM4ZqCMLeCZwPagu0pXpYMvhOiED1k/M7D/NY5yM+
zLZsmzU7cAQdg5JFfpXbfXL5QM5690MS7aw4Gb3hjeUMYFgxTYmrHSU5WfJxBKT9iZKR//ThlK4v
iHK+8LjIin/l3QZQDS7DBkE1948E89SmrCt5rT/s7PRGsljdntWfH87/n4U0IPIw/Bsh3Rm/WeOj
FW0esCYoSBDmOwGKZTF+uZ58+H3cKNx+J/s37O0p/2rzTOn8RaYH4jb6aAtT8XqhwqFlSSMR332a
rXn9Q8+sJCBRchY84vNQLRRgVidw0SHWgpoMrZVd7dMFTH5deF2gEEee7mmHnA/06LJpRsc1SvO9
H0u6Y/7L/WW4QpmMCwOWoY1l244DYgniC8ZzYZssYqJ4bJdq4LO38qC4HxX/TDB6Agn9KMjQ0dQW
RfLfX24UbaI0cWDYaGiKzemykO61UdDuypVhqK9bQWe2h3CKZlM4gLAI73jG68tgmJa6lGlEQy5o
5uNNoHBXebAXkXztmNseMLv7zz+k/HxDAf5eo+6DDwQzVEd3yuvoBJgvFmBG8Df+V0FVZ69Yker/
qq+GUD2nkHLFSNxGP5awRerKwehmpn0AOBdT/fhPs4ZvRy+iVqFsrFWGMIXOJZo5FrWdXxG8Gbkj
JmX6vcFGSjGaU986uvsmiG1cSlpNPj2eLbL6yRmQWa/vJzwNcEge/pZfAByM4kXV4tNm/s9gRkow
ZJwco2yLsvIZKzUAh36194rXtUkPA7XQlJixswjAxfX46GUqUzLEvuH2+nk/IxKTqC++xeTMlceR
IxFOY8j/HD4qXXPVKbgLSO8WHNB2ML2QclNW9d57mzGpNd/PwjTGQK8ZlS82/dkxzJAlPTA/McJb
6S2/aE3fnbQowio9JCMhU7GdbthOvsc8A0ScsO2j5CCeQaEtzIKGzOPsfGxfdql2XBBFbSSDYdlT
snufqYfV0c/a+vgCAoOaE63Ds7E7WnaunbnrJaMFNH79syS40hzcQhv+YIRRqmOLB3aypj8low7x
+5Lc95OK4mSIM7/WPuB6kbIad7RmhoXCy5nvDiqoHk+4Mt6gcbpnKzkVGzENxjQ3kVv2FkXNKlg5
RxMnv6fHRvSZxSnBDsj7vTssCahDuw1vdvZpg2tnxrSXBR5nSmcehgRRNERtZQauDfWST4ANVhnu
yj579L24Ork2BoV/+Db0F37IkIZ77RCXaGWgJRBZIvnHuTIgIbDV5V8GCLi3oiwcuHGJRM/Biadq
LhmgeO4Sb6er068RqBtdo7psHXgaR6wRE+YW15LhCIlOJnn21/IQgFzN4s+kJ99qV7/fxEmKjXIH
8YgbX+wOmyqbOip7n4wPtPAmgreyr09pRg7s0V/8NGUU7F0JojAz/l76TWDxVjhWtZvue6AGLyo8
7bV1qnBlNr3aQQM9z6KpSfot6+jm62USKb0kiz+XfIGBoNrE6WaRLG4ZeyAKu2Pql2NXa7GWI3rr
7lzJF+F03AQFT8ptjN60dbTK04LTK403hZjb6GJa9uhftSVPsrqgxePEJlhFcL3CVKwpgFjO6F1V
2AoXtRTKdF6euKYg95T1k8wpW21s5dj6Df+9cQcEVgk9NWjfJypNoOGUk15A3RSdCEMv0fiiDc13
bP5d/Ox33RP1gcKQjljgTcP7LSuNYX5paxYp0cSp3sNXrA/a3w7smKoSeoRnOjlQPPDzUmhSv1qz
73uimlGEkShJqcRluNBWd0s8U/qZG4YaNiS2cDr2G6Vsfhi6P5YHZBe9dZkZawYS1AgGEvRYQs4M
5UrJG1ONeOJ6fTjJd4kwF9Hu2AbH2F3x4SuhN83YFyHJjANwaFBbg++E0PTmuun7P+MQkpYPt9gg
pnqnDruP09daZRgFYszPa8B4Sq71lIkZZVjugB+kc86bbOa9rTCku06SiDtcfj9PxaSREC3w3Uk2
NYb4zISK+W/rek2rFb3AbY0eOKz22e2HRx6cBf5jZ+0Z9s3r7KgoYOCR5JA9JABGLszOJbb7JeVU
iSnOLR+bwIEcDeRNeD4Lf80babUyH+L3wQ7oKSvI7LFK7gq0Hm4OaGunNyak+PCbNptiHGaocphq
YC9rBJV3aFYDDOYRrqT+k0SPFKOBjVRVT4+InxIZUQT5C8YIZHCZRtprd/WsuQeZM3QMykDyRKRk
xieUJRdTTuz2modSYV3GlTm3FbN7AKjwtfYlpFWi65xSPfPHymOtEc0ENRXpTwZn5KFu2zyH3Yf1
tvTAZF59P8FJegmgj5UT0/0cKzAzfVgyvW8o5oYuRvlTsgRm2Zf+c+vq9kiyMuBXMvP+/WfsewzA
Dfef0LPkQXiAKfgI6+DMbUGDUfJ+pnQ94nFZFIXLdESBcER8V6W1gna8B0s25esYqMT7E36eiNn3
E6xFoYNklIeEFeW0xTy0cEvZuH9eBC9u9VfnbrgF+B/RW800r6SYpos815NLRRlWKMy+JSN0874R
SqDYhZTq84/v9pi3r5tcxJ9kCfw1P+cC76W6MRSTZ/keFHMGaItZ7M++Ws9zM8Qjh0Wdf4Le5bWA
ih8xBJZF9IwOEDnAnFSKxstQjegXOmmuRTiLgRpfwUM/eQOHEyNGpW+n4aIkWYOLtXsiG3iSeDoc
BsMWlhoC5HQX7pJBjW7XRtMi4EVnMDm+153B3pErarFT3EmZhV+XdMROgU2bDUdX4E8LbC/wN4Mz
DyVwOvKBZPsakHrD5kk3/4nFkRXZHAdEH9mtF0EealCO+rc4QZpe3dNTTVLI2udtk3TTCt8mopl7
Ewtv05DE4zHWskjsVQ/ZjX6ecU8io7uImxKM7agfl6fjdzudyjdCKCizJl86fLZRmilVyMxAGAu7
H0FhFETQD46CFX0PJjFSXI5QApYQAmw7JqSJkk1a/qF/QsOsObJeko3W6wp6acoDcY2ruSwrDE9w
cixaJ6BYVD5sNKMU/J27shImjcQHpMXZ6SEsnlhQnazwDYJ6Sv5xU6Sye3j/xwmLa+hRUo9T0y/G
LbDhLO9nBlInotvVl3G7IOkA+N80AzJr8KQAHhyyYKK3G40tnuVVXFd+LtEzCz+unwgyjnqFnTw9
xKWYA9ifbcBrkOmAOiTfbiunssL5Z/KKb21Euof3I1oWmaDA+w9wXkWuZGTR3abZPIzS6rx7fG6F
0OnF88xc/tdX+PsvLzR99urWWbLqgRZedmgQ6xrS1Ek6SZpo2cJRbLyZuBCzXYwtFBWA/6aYeFsb
fpVwQQJAO9SlRyT0pzdDppjEnWoTdX0ne4Q4IKJRQuGBL5vz+yiTay4kWRMOs9Ves1o7AdQ6Ph+w
eNhbhgl1JYpm5W9+Uf8KKFh+f8klUgN9UDluZNI2Uz61AZlng0gu6ptUnQZ0LPSjcREp1oK7Epgw
f6+oSC+iHDesFi7LKzo1Gn90hJKhBEVrDeRnG88W1vVoxuRPI0b1aRh4H5zrdelZOwKUKwKkww/l
Ok7ztRyGBMAmP94WP3KzwjE7mGTi0tECQaRZmMpGlcc3Gtotme7GIKPLfBpt+yHRthKp+e2xkA+0
Ui+uCTNIa6Ctaw4nHzsNqTCjgAbSJqDocd3XAM32QdHNqFPP06x0DUp1iBJ7UDQUsjXK1WebCnD7
kw/L3DuRdcTcapV6gT7bA4W0p7FO0xlTsZZbAe2iEcGLoGlwwg0wj3n5mSyJj80w7w7gw3Fn3zQh
CS5viHfsofj8RCdwrybDYUJj2b/wXdW0CiY/sN+8hSJHOKV29m62oI8gW+MsnSQp9muix6Ov8u/u
Tkz7B2LIynoqz+BLiWhxgCYPkI+xB3tBVDVBFXdOB9+zTuMKgZanSOuFuXKNOQIRNjDfceDjKkWx
H/MVa3RvklY3qiiuwp2Q1Z2vZFfn2iE2APOKfTeqknTv/HQwkLkp9+M4sDVbVv5aUj8sVOU74o5D
2Uo0dziH6kTfQt6tLKyNj7yhjHK0qzZ/xJ63ROtiOPth1Hb4kQ3ABgekvRsEiUt6XnK3d/cIkCPp
CZeUv6XFBDNJZ7HVoYaJFiE7U0oWyXtNtywzVZ4YUby5S6YmzBRSUC9VElXIJoxWbFARkUuKCs/b
ElwBkrKK8b6dIKBhYInr1Z56bfCX6pazBtUgQAsx6yV4dk0SmH93PsH0Vtx9955YfU7p3y5E5mYr
jLftNpD0hSgiXdbIX08m8f/Mt/zPaV/AslHGRYpzftbTHGQrIBjeUeKDHLnjOhXfb8uIhuKL4ycN
OfdpQ9NMXhm1iDlli6R/FMVsog/i7lHB5sJ9eTw9F/AchhQiznX/IBvc2puBsOPDbRBLykxG/qXY
vIEHYgbZ5HkIGOtnZ6csRYPutLfhsh8B2ClttYw0FAUIxRTpckIhxS77USpKp1jdqYVx6gVgkQY3
P4N23JyYpEz8eNjqtG5nA+fosSCzLiGMqdIeDt+48AWWMQpw0ISaaSxsBZjrSjsgelz3tYVnqZzG
CneBfcZI5v46WhgK+zzpjx8Q9dONliVz3Y8eMRGR6QfmSRjxsw8gV1aMMyFvqpBuH2BON0vD9NiQ
GRZfvukanwHwzDAjEpvav+nsrpBRPzIyvUhL67PxPIosvtAwJ9wqb0znCgJsPooVZpqlXoWn9lnf
8UJL+hlJEgkAnv2CTCUBt07yDVRUvZbc3S78sJoKHnxm1xdIXV7XGNmQ0CQLgDQcFUJ4gpFBoODq
BsjV4qnH/gg2yyxVDljTrIyPw9LzfmoWoNTNrFxWEGc6lDsvoLyDMYh7Qfmjl4qnIdsTWKE1BNGZ
SZX+y+cEYqLBs3JPi088NL2SGyM0Dpuzb1I3DGrvMXtjpvXJTTVkBs8zA0OL5OLODWtz0A8Q3KUL
nmvUGYvOwYevq7p+O3YEGc7mj/0opk4Qk1UnkSOZfu1KwV7kyXzFEFSQJz4Yd3E62z4UwSm6sy3f
oCzIAeOCeD3NAYNzd5lOU2Ym3cn+Gj5+7avO3H8ulhOYTDM2lRR5f3tO4k6J16akVm6wm2FIoXDz
AjJYrJEG2AIym+jh01jAh/LH4ZFbjidnfd9WJ8b7qCZgBXl4yTsDNT0E051eJwbUhsL2t569fHh5
UwJdmIOa56vqf1+9NsBBU7JoK5HfGLabSdAIufbydME8pjPRQjNcO27yVEDe9ru3bVsmwN0Jh2X+
tX2fF/SdgSsR2LIZHC7Z+m2mqqi2OtoOEB/xzWtgOoyQQ2xOfK8Z/axrIT5G/9VS/Zg3qSczp2x0
0lfISCBoqJY5HWSEiCoWnmeFZmSTMFAR//LM8q4tNrnGYUKtpV0FmZxKAhP6dN3du3NcZksnC4k3
uZHA9dwFwzufPs+O4ZbJsqxLoshuHyDDakANIjzSs6dYPqEG9EaHBrJHWy7LZ/Y7ntdv8+9MwF//
+rd5H/yNNDX44AC62kvSXNqhAfmIb/ik45GSbZtj6ZZ7md2Dba3jB3D9XuM+swojM6IxGQLVoqOx
zJj9mswyk8BkqXPI7OYjb34ErEsBEKVD9jpvXBNzHMUhvh6fajm4DUN6BgeFNHVK7GxzoH/yKV2r
z/CC1SsN0rIA8IAz2gXnllL6MAitPHG8rTlGq2DBARHgcx4YtppaqZYL3PHNOPUx83gr0ymeMTkw
f3tlfdtLTkoxBQfSey8izOQRSl2IU8u8FijfpHeeglBSqFJ7cTVwUr/kXrGLGLer0AVaD9VrrRtf
W3KedKD+Hx3zeE1wAwTZcNfEoXyWGSpf/n4qpAtEqk2/Ec9j8c1NFaqAj8Dijv/o26ufPY3BtiGP
lP7u/ackbP7H5yNdLxzn91tJrTQaSDI+sNfEP9K0qqstUexIIt2JGzOS5FbG2n0LTqWtigw3++0b
/kOw7FAymwd0uTbe2SlYInGcttvCPj7WkwEYfAhCe/EvCXwSAxZ45uqB9YhTRFDzTbJqLNimt8T6
EK484J7WTvYO7RmN/MJ0IzEQ3T168E6oX9GEtV3VFNZkjJxdNBW4eJxjoyOLcIV1lI77Y3GEv8x6
oMOUuMsUEDwRjU+gesTGo6bMO6BUHG1WVWXIkB1mRpudBVLpFdin4Sr9st/xedH+CUzVsixedKFO
nSFpO1uXpk7dqGYiAsc/J11F4Ap1sLsyVGNfye/nm9tBfwZ8Nxr+Opgh+ubCSEN6jIbrSgbJVhVv
TGPj7QV/+nH6brMGu6ACtNRQ/24VM8pfHNhmCPmNPO/iQXLjCNAA40MWvRA9IGrZOOX/QOAYAWTx
LVo9LCgFFWPz9J1Ww6OjKLHLQ+9hLKMm0NWkmmusGF3zZUF8U8w+o3fVZ+7G5mqXUmaoD2txwRPo
WwPQtPAJEg6OFsm3Xi2pwkVPyFPj1qUJMwGOyRrXiy1S33vGLvBdi+jUTBcwicYhLRUnNi/vQvEX
y4XWrOsRA4jMctdBmnAsfHeuD3x45hR+plsPF1gnzKv0EVYVS/UNK6sJdkNWdclJX2iNH739E8mw
fOmq8epQKo+dziupJiFl+AAIYisTBhMLHWM0ldSVz8KC9dZPoUutCcOUZZJcx5MZHhAuVDbIt3Vx
M7OqLj+267MaAIk4zPUBfrb/HXlorADd6uz2QM2z5FkZNkhEX7BRZXctGMckz36+5PLgvO4pKkpZ
IhBuVxlwyiRbSgX4SuOI6CzJEa0R11WTc/e6OW7/RdSx4V+/xACFzJ6XVYFtdBflskT86SDRKYoT
pYP2UR2SfgQYM1yKnfSxrI2wAgrX5iluPRCuhWQD8683nqkp+xiNLMPYfX3p/PhoTWLD90MOC6S2
1ZkB3ZtcLKFKszYzmeut//VuTc9SECEVdvcKvsXhrEEdNpO+nMVe+Piu8LAF9ykEpKJVAcCT0k1V
JZGtDHNedYzA8andelD/zhgM6zoAKQ00M1pAtnXyESvBfdkGIAIjDAvRQ5n6MMvdv4Ido6McgvRr
H/PEP1Y3Xj6JcNJgcF3GsGUkv1Q9belSUaEyhrlqFgqZu6DbDp6HD4G8h1/ZZVsx9Ub7Chcre/GY
DvUi0JfjbOrYZUpTj5T+aJvMBm8YV30z9MRu6lZ0fkuc4XcIcsblZIFwhcIHNZ4BasKwxvT4sWsD
KOcN4s0dBVdHQ8TPmXL8EmppdOmAf7cKEbIfmJnDVencbt07YKqQJqZsAVypBKMhaXfFVvPJK+YQ
Y2kar02fRGeb/73wZsnmhYX/QqOrHfrbj23+HjP/mcnPmHEx1B0A41Jm+UuvhASWklk43p1mv2qz
BUk3O04ov2zlxWN1CWu0WC/IGxYP8nYQx3H2EMhIyuGnHZM+FTKbOx2fOdAYneMoDgXCTnpIG4Md
4EHajDHfBUE8/ZYkNZrCQ2rUUqUOjX6GeFmBNnHyLfHyzLP4PgnGX3rt/bNmY0HQisgKv3swUZE0
P69/0ueTKZArXJjdzJVdqsEimP79PPCLsKDHAOPJHIQzl+zoY8+mUoNmr0BO5aqvCVR/xkTzZ1Bp
oYtDIEHJAqKGLnRjAvlQMhbID79OLv9dJQwoEae7cpor7chJxlk1qElmuz8ZXR1XH+60M5wfiHOs
5zJtK1iiUKknVbW3sKeXMS33Dcer8V4fEur6LppM6+Z9zFmmOOKPY9ADPbJCZP68GLW5a5/FtJgl
eNOzgc1UJ8Kqgx0XSNcto0wM4/dsPolWLYQjWMQXqzaSkf9ow16mhN0uLtv9A5OoiX+wzqgk6khk
YfpdgHElGeUhIf25FkMdI2B9Nw92QU9SVsi1AoNHn/ejpk5BPXopHWcbafU1OcSpsm8HHdau+39j
s5xHGLs1r/imZjZFrL4/CNA+P7nfmP5ZamM0i1+3CcTOBNNaO1p33FyTzWO3F7AT2sZLKO6CdXm9
Xbta3QPE1EdCaO+wEBXxYRJbNb/wuKCeG3OyNnxqM8xFJkjLeiToSLUniMgN8VIoOcUbBj2a41/3
RRRkX7bItRkTl79nqkAIhPuFWz2IQRJuTNQ0gyuQk5fvI8QxnvUyxQj4SthXA32e7S7iqduoVvrQ
k25ujRgPAXAHEm1nn+30FStgqwHDe+EuZ3vPqpLoOaouNiEkywIzTevQk0UeNaaAB8NZJBvxrCcp
eTFexUrGoCx1AsCHaX1mp0Vx+BL96l6an/Kqo8T/0XLc9in13eGulLZ7Q5sHZE+0l2tArasXgZM2
tsdApCRm7YIQccC5y9BKY1sJPvCF2AcJIb68XlceR3kKLp20XfJgigdGFvWPOf0/W1FBr4SV8pJx
OZ29kaz45JhcJWwtf68iDuAqQ42h/rTSZYfmY42zdQ0UF9iQfTczgKGuC2J5EhrYqS8xr1t7djsC
EEwxWN+THdVHh7/EJ/+ecAMI3l9MPAVqvoKSqE40oqszXWQkZ851u3ZCt/IWv8Bj32/Pq9CVRI6U
aaKPvTWKo9sS50+/Qxf5V+jZxfo3RAEBWalyeWB1RQgjJOghvG69ufbRi9US6PxvAq/bmPtPywkN
EpZwhnOi9IAWCgk7ZEkl2PiAvJlnEbQBTZRhjerQiZ0RHN2kT6n2ZVzojwecxdrv1wVTnODUs4aL
tatq2IFbq0myS97zyjIt2TPzFBL6BqHqQbNBw1rZbanUQAEtuOfMUkST5MRXcw/Pp/T+dMZETqdh
Nl2CrKQLyXM5RO3rehjJCiwwTM0iRh5W0j2Dha9tE2+3Tl1VHKu9HJoozY2OYVTiHxVOLxtjqFbL
pgSVMGuPWQyC4x5JKR/PwBUIt7v1LyIcFtUecUb2pIwiYU1yIw74pf9z/BPFfsMIkt0yH1tdSB8o
Dia01QfPlDZGsV5mkC2pn65wjAPA0MaRDsOfG8mfDIBp3SjB9cb5QplazqmZ3LiIui1kwCDbqPwy
AFhEPOFxwb3de/ZZSy1gbpQ40+BUV0CzGVGgOuo64kl5qOL7Z8D1ZyXdsWlqKXpvfNetj+tSK8UV
LrhSMJVsNJWOrPgvEdjH3IBMT4eR2rbno3wNFNjWKdNDT2+hy/3zzmiW2DEzo8ouTT8DoJ9JzowK
sHs8QI6NfLR2h+mcV8MyD/cpCt/L0XUiIuxnsVqB9JPho/BqW36HqmcZzdHIPLHRFiHk9iJqN+yb
KSYy8Xsgp0R9lxhJyozOHoA+pE1hAqPfibroYkFpVF93hdt8nGdvhkjqGImW0o9FYM4xxizD1Pvc
1sQW0r1cXZI5m6+QUiBiKNlKZ/AhK+HYvwXFH2tBbAoRBLatPxs48W/XKM0cT1OzmR54TXQ4GjMU
S73Ky1qE6HynpJQxyQdR4RUbryv+s0g4k+tLA7ykImROQlynEQsEEob5Wr9CZ0pCBipVQYw15xDw
58T6T445PZGupIMFkyfVedv52gYgusdCvJv5onUbtgMzvEn2y++Ep1LUEx7I05Iivo8YZPIV2fWg
65V2DSvsRl4Urj6+jcTUyB0IXKFvvmFq4OmVjdohV/Jjq8ivhxv8i00wc+PqYTu9ZfRsSm/OQQd5
xH6ZTgrGRCYF+pbw4dylrl9+5BUEo24VDn5sbxDS8xk0OHqUndNfYabwL9GNVOtn0+O6iHnAxQqV
TMiVPf0DC0jcVS6lQ0G4Ct8MjKSC/1IqG5qLE3Q4Fqnuo3NtNeJlTvEKIShTJj1sOlgIQL9ri14v
4OuqHk4exD4gizxyBUrIdAzAO8sdgzkRYxejeuiZ8j1hZwzHDYmBTY0fSK7IjfdEVSZZHMqZfSRT
k/gP7qQq0aJjyjHdYD5t0fFHll8F+zQCP4K1DFDCF0eT5yTG8kHmTdLnLi9PjWSYMDoBjq8vQTJm
fA7KzH/CIRt/Zb/EpQYyNqAYIN1vV+ETwrhc3aIZCogpl73oSIENPZFhHAxF833rLTnlIo5P/dcs
Jz0iIg81mdjC7xV5gdSX/emOV8Ibj0RQ30sNOi4cTbR3Gv4BMA+OjcjdwUpoImxvkSIkxnK6FG9m
WDBa9+LGZzzB/MJH3AqoajHtkMRtWmoagcBX4fYYYD+RuJNmnyQCyPpI1z5Vp6RGTWh6+by/FBl8
tssz9JMEV5gooJS8TMYaf2OKvjCnkWR36INWRS3hcOpdNwerH3tDcYFetOCJSLWl7eB6nnj0AbcU
PrrnYyYNkGSEzlvb2ONFHlvf41bvwbNup3XDIukMO3ioOiw7ymUVKEgghRgG+Zl1uL7Avu8JJ1Vq
H3hmQL6hF3sP326Y7f5NSd1ojiNCcwryFTS6lXCFjgVB0yb0AhJ121FlnyapHipy2EnLw0BuAQ1j
NpMmzJ21ERqJls90HZvGfJpW75+uuWqwZHLtWYUss1G99AgI8LmA7cUsdM0EpNIZt2cDsSuiWu1H
Xtr3ieQuLvHfDhriKHIcqFzzkFV4T8QI+LCr3NgIlHRZG2idtuAHL3Fyavm1CJlXjetzTipQwPIG
9Djo84eXkuIoM0yPiT5ne8HoSNbv3agiDXYnXE7EiyOAgv44fqSxSWIhQf0ATSz+eIBVBjf5aCqs
aYWODUstwXIbqobVjDC5UsdrkayyB6AqYbCtC++D3rv9+ZpmzDGiJDd6xZdeJwocLNdXkCyMASzU
rbcqfcgiuoM7y601i08JCt9sbNT22vitLpJm1Ol03ucejxoQtdUJ39SJ38mMOaZO8+E/TyZPrYBu
KDJ7flkAXGw7feZcRgOc4ztQ4Mnpe9HQAret62xEfpr1S16EoenFGkeYiVl24VRbNjpybUGketoe
JtnrOhSepgKeY1FSGI9OX/aJ7n/wk2cYPmO4x+YNpwZNeVo0/o8A6/x/7SSjf/W7pNBtEwRsvH6l
8jpQAJdcTTeYhNHcq0HLGRESEuFSKfP1e1tP48NJkiAwHN+srp7lDNi5foNmRw6ZdbLZqyTNWG33
cY40AqJMe/+X6qe1RhdQxoQ/0mjg9VVoA+TWb/lkteOSkIpFNxAM8iogqr6M54GzKuBfDXHYX5sE
Nsp2SB1qZMQ66D+lesFMYV1NZeysa9/TPe3VcRjfEr0ncbT9hPfDxzOB0lHP/oXsNiRyqeor2Rrx
RqaGYk/3Fy2MbOf+ng5GQhxcaLzM5BXPf8G/yAqn+4m0Za9eKdx2UkTiwxKiM6bOP2T15vO9q0xX
7nmyNcKSsaM2sD+C+XmzgPuXwtHYrGt4VKf4afooIn016NYUfIMTP44kZrzn2Drr69/ZMwYueQCh
YWO7IVl5vVzIhOQxV3ZWb7KuSiCMqPa5O/MfBLr0bOaQOzGfHJEmE6OxK6HvdJufqg1aqSOi19GQ
Jo82sH7c2sQDIX4Cpm/J3XCjctBOyCcA3wd10AsQj1xCs8N82tgViHqI/4E4XECOlc9qjW/YIE56
/pbwcfqJ+5Cwc2eWqVK+JuG5VkIl2xyVodGsgcnFKTQjpHKsP5xax3M25lozC+9Khz6hl1OBZnJu
LsauOr11bAG1iQgx0AL8jm6xvIZKNZ0g6vTqTqbGT0nmpK8dAixwHNDjHDKOHiWwSezMZR4H1YJI
8HDmWfZhBREVEnFdVtDpQW0D23tjQFDBTt++LtlYNwwUqajUWzzvtduORK54l1K1QH9iqAt8UgN7
Ku1ixpogcHZqEPwAfDEGiHqYU2V1Xoy23nrRxVrzVyNsWcux2+wsL+HG94RxZEh9GxpzG0JnX4UJ
zn++SNUfgBUtrzkhM7eRwl1Y70deepgpi2fuyKrxCiHIZrrzEC+Dv/w/63Z8Wle3yYcRB2gZxZ15
Z3ANxVt1HY2qbVcxcz53WmtjoLL4JqWO7qqJjd26X7lpE77Qmv+5FhtQj/pn84XWhTHcl1pK5DPC
vkn3FnBaQtnDPe7bcYiphqodI9uPaManpDNU/Ww3JNJ6x7OEFaBxqdO5d2cD5rtOEP4lUZVknY+M
av78ewjDVcgd5bv4OHbbIhu22NU2wndiKCW2ZjZ6K8R3WAzHFjHTJwnBNuPxgq9grPReWuOZFkym
838RRK575+MKy1jOkTdJpxClkSviTlqntDDjG4AZfh1eyxe3wTgoKOJQ0lQC30BaD4my8D+XDgGB
oHcaxuPQI6uuqQYu+TF+YRBLyB+BpKVKbcx14x6qHE15OJBanz9QXGHT70SYSGoGPVM2Zy79e7E6
D+JYZzLsDqwXFvTo+DHXm+FfRjVoJBhYA1y8Caabs49EuhP8eku2DE/cqUKg4RhppYRrUAkhv0Y/
I2ap7mXr3tZLUs2xjeb1IGyhFny/DLWk+8tSEEYwlFKmpD7Nq+qjSHPyg0lj4jf/UAI9IS8Hhben
w+aUl1DFNcmixwwlSbNKJRvtubR8oF3Hlgy7lfCeSGP7fHrpg68SNvnSHW8ITgjVHsPh7r2OKT7s
184XIGNswL4J0QejEEYsb8Qlpsy7Vhbx77ZsGuTu27VYwcDQ5o/iG/u3+iF6lgYQg3H0ss9EC9ID
z4HYRZY2dgYU+eLJ3ipNPY7Y/X0RYG6u5QWH8iHEoHx2K9ylOWb/XXLpO6PJ41YtMeoKp4/8D0sr
kDSp9qb0zZpvsuB6oDZyuI5+xblaLmfYuj1Pm6oxNL+3YblQHHmo71plAEP5+woPexW5lXlhRQKY
lmDslqrr3sieayvUTbhzF+e1vFmI53ZAZV3vMbAHxv94Hw88+wdO7ZarZyoqbR/LRB72z144ksQw
Rc17paOgVdyKAHePqRZ/ZARL/odvn4X6tTmfKRvYt9fQJ3h0siBLZvtQsgyUCqPZ0Eklw/BF0plH
cHJ3VmsyXw9dSopsdOAkdvT74NtKX2tt7V/biiaLlCQTI5BfHaw0pWyqyxI8SuXBm3cUNu8eWRHD
IctGQi6D75s41dZZXyMfT3QPAGaEz4QaNh/WiW/DTYq/KDlnCwm6Gy7Cd7g1l9gyIta0nG+ayYpb
r1d2FI98FMTfF8STwGXmwDCUOVSXM8Q1lvi88ALJAHiLEfK6Tw01+hVUJDuQ9mpQeYlpKOqJ5fFN
q6/giWxP0DaS9yGjBUrCfO685r4I9xnbgYlXoHKvlDnNHwWD/CisfnJbffrSDQZyfG2Q03rhh4Fn
+k/Jdk7IrEYoIK2ZkeVV4rGI4/2ZH/3mu/6qQD0ellyq6+YdF8u8kCalmssJx9RUoWX59snU/i09
JDIgQwEEDBk41F+Q46oQRXZcL1edV0n3hpRaWerYekb3P0EPp3nQsMAowVKxKP4IlvUnZhky5QSo
Xm0R8qTKCkUUB6dKoZ7Hln4W8RF+a4pjpZt09g+DXOBdQr9JLWf2jlb6JuZ6kutbV5I00pu868i9
5cY5LoPzWaUAnFe+50AfW/70dITGB17tCbY2yQNGe/hN3RHeCRkgVGANNY7yysbHPMOHUpkIdQkW
9ApJELx5dr2phr47e29tcGkoOsN4I9mGFE3S5Hik/EG5UR1+gjjJSlto5MUEsIHTTE+onqHi8zJW
DujBjXVSu/4poqy+dDr0a0x1WFMGUYf9CG1DgBIZdQqFcpchD+4Ys9J81pZzrO1xh8yCHd9c9cS3
8YoCKRo1TkFKj3mnKwBrFKDBFTONZvlfmCHYBkGhhxBjJnsL6cgThsEpaQxAOJ0tF2CnDLqFcHSw
ctIsI81vo/1aW70sbZMR/LIn1anO1zMwZcSDD8GOlPRINJmbb3RQ0MvgWloYIUUHuV1AMwXwjNQ2
evm4B67q+9kZXzyUD3Ku+DWOoBSS0sJKlyBpAbdRAGSAquqyMKz0n6Pd1iKVVh2YsRyZUkKOXscP
GKuokRHZuWYg8DzyPmTi0kj9IprBnRSg8PqibsQEkBAJpiywtzX0kDQFQm6Hf9n+D/gWvHJn3qCD
771QISSmheBXdwV/x0RAeUaOh+oV+rMugZkSVhkvt7+hwne4s0K2Zxt2EXJ6zZqnrxWXFjbaXQmC
2T/pmOql5/aCGdb8uT4JXSZF7/WQ2z3L2wZw1eG0U7BxjzQG66mugI5iAVMoWBsOI2SJBzBTS+Y/
G0d7rGKQ0sJXko9QeJbnIAuVS6QEJmMDk0RNCKj8JRwoni4hpbG7APTi6eLfX3YK4S0/a0Fee9Ch
WbUXjLig3BBiq275q1U0onWCRQ80+bGxmCjZvsMlOZJqe/8ie1SidyU1A2pXiH/7YjZb6gU1QTOi
DzRGLjgzKoCZ2uQIvVIR0faa4A1+YCEKB6StJ7Vm1hRYjP8ZcyR8JREDduzYgvci+Kar11i5AtHo
8PGYI8zNLIuIeGniw9Ica7A3nWO01AW/DpgC483XrRPsaVy5uGfhnjfJBXxIb9H6BTV8pNLi+xSJ
weXDrAscaR0K2taXok8guGVQ6xrv3kuXxrJhR7iZqMYeAeR9d1ton+23f1qX4l/PBrDoyekJrkoO
DRtxk5S3v3Bz5/IrZk4SYWTsblUUYj+Rx06yyZVw4HR0u7wpXsKeSIss4eTQ9khfuytv/q0/jPId
UE32cGS7n6xUarhwtiU+pEmPoMc8b6gfhh19YjLbafVqBp4J7EocDxqLkIU9cyPG9scaFgsvryv7
v+/qDUEnv6VicreFBK7sw4sz3TyUWWWY8twRllcv3r/Imp/uqpI/WzxU6j1gL32O4mBEfQ2kuuJT
L7NCyxzDB2bkj1biszYvCqdhQf3yNwSoGB/ISqFodNHv4l0gRs+q1mdtBm093HxWRbBp1yNnz75m
Tfvtk4/MG4LdscSkGsodfjBZZVGrPV5E0H3fb8OGwPqsuDxZh3fPWsFC2yU+0PArzXS7cdiDKBAh
hmgMj80wfFrHnBaZNgLdJXoo0s+oQzD3LAcIQpqJLzFfW2dUe48793PIsdSll1818jUjcTKbEmfB
1Gns2Mb1X8m1zKzeWMwCGe+Hmwzh4FPg7PmMgmuij/NH1yU2fTASz6gEcLaSNLOlJpyE+LTvbjya
kwQuFCxJSANxKi99PwPri0iE59bN6S1N2SQi6+Jc3CwSLRZIR1ikBCpS+WUcVqXKma7/IgTgHD9g
RS3mrqleCymsQDtrfUESHtboXMrkOwF7Pj7bXBjAaNjYa74rs2fDghxZropTrDXmqLDJywK7FGKP
k4lrOJfSUBJrJvU4vUX+bYZ+b4rcauXZcP/HBEwjnywttHKzEWmXU6jKN4laUaRpd4VLkrRWCygY
HQzg8fMvYThGwk0SaCz1GLQhzRyPF08k34LK+0mNh8Lqn0MMcLfqjbUr0dZPniuJSd/TeSbgW/yO
TE+1raneCElyf7iJKjyxJHwMqIYNlc0xVOHCHxb0kinFXtIzhKrxekOpqi37uCljM7hmnIIxLVjz
55VgwJIUlxdLthdD1zY4IQ5V4x5gbeCALiAIC2UPc+RudnbwIkCo5Yyz7CY9ENIbgmUzB0l0N7I4
NOyfPsGukDWJbZGmPn+3DcFGMQ84a9z9TfRUeT34fMSxoS33wanWghkN0/x+54rKEZn9d9+WeY/F
Q2+H4tt4H0VJWx3ENOMLJ1D/C87O4QZi+POI6gB+aQYFHBGnL9ZMpPU3346OtMRmp03TAaXAVxm0
3laHEwQmFJFWRKbjNKFlD8E9m66aA44obmqpUuAc3pq2XHZgb09ykgCrpE47G7mzFAwO/vF9gg8t
ppQmKziL+Ia8b+74aMrEABXcs0imhbJgCKxXhQJkk5rPRh8eecjmAHmer8gxIyo2zNhiPq6TDiHW
PbAAbZ6c/CUCMatwhOhWruiBYwsnEwvpGstCs2E+pFcKh2FROzsHYE1H2N+U632alfx1o1+dwuZr
YfLnlFnZGp9zrzpcLpSvuZOT2tMcABwfZeFRVXvuQdglmGVJ3pxlnpF0UfCUKKjqdjjdHg7hNvtQ
r5RkTy3+rnx4tR4RfyI5FaVc5s43yggh/hnxWNRSnBa6oqoEwk2KhRU9ygXngvfXXnZ+y9wn4vVy
JD9QkB/DuF3nWbf7eEeljfFLtX1OlIvBD3VQWgqMCYk2UKALTAVH6Iiji30x6SYJj6vTmGlnmBbo
HHruAWvPvarXR7a2ODw4yE6Avsr+IkieLhE0CCOsN+HzpKuoiAPpEIfW44RZxudjQH59Q9NlbmaK
Z+IbFd91Ch/D6P/Hiqf3rVfxyYE1ed1ANj/zEzA+vzcvyHqhaONTu7WnMARly8MbPKZgkhVNToOp
ZdFYldKdRnsO9ARYPrVTJopMGY46ts+EhXfMSTbDXBOrKRdd/YjHo15wcKTsGYuMMneRosgsK+e4
6I/JsWri1VDH0FcKtVBLoKxPvG6AzFmsgrO1XusqHnHBafHG3dfrLaOC6FBryhgDyl36VBsY24JU
In82e3aoC6sFCF2/NotkXHuZ4dbuCXkKnyhaOIxGkhysJ8cmcH7TltzpPwu2CrkXt1RVwZkkc8d0
9GfqBzPnd4lSfyB8W9hKgW8iCsFqH11NySyD9hdbI92GeQ3cDeOLAvmhUUqu1XdSw/cmtZ+I2oXo
J7uHM4FHZhB6B360WW1gCUS/bD0KZE4B0UjrtRCv5xh0Lr1gVi5rEkHg3nC53SO7rlEWu0P7EXQe
Sza8qaOeBgGRu5vwVEWzdV3mrQoIqaWfjeRoKmSkBMe98V7y3SoCkabt5aqwDWW5vUs9lWvaG/jW
I1TuuBABZCy8vxsGJ0VdFRSUiFZXibAC9IsXldGyaDtV5xPfojcWkdi7poPFgzYAZrNkGo/paypQ
d3a0HvjOpNMpdRLilTcRflbZv42Swm7tBqsi1vcuvsWpIz2cjm9SNvhWUosarCZtoG2+DPP4mPxs
RvF5k3WOGGdK8uxFrhTXUorxIGJUd2C9F5q9njShXq+BTKLxAcuMGUaedzdxwJO2Dnv77AzDdouE
Z1E1/Ixxnf3IeEDMWV5mse+MY6d8J/VXat8KteAmYpPZ4WDjJdnnr/fPn48BO20tq8/UvxVz6YUw
lJ5m81Gn+Azw4+MfKpvRBR7dxdcQPFM4aoYNrUhc8pIDpZyaVbcv7ngdS4g1CZmd3vjRofu2yGA1
p5TMi5jhCij8zKDR/golQroJR77O96G8NTUp8dr5byL8lvJBhsIHQNCpVnFYLsaIm61upyEbn0IG
jqeFdnV3ZCiPBQlKMSJ2fs2PbLE5VMDbpDbyapOj3PA+uJhMOjDBWf0heFDftgJQ0QeNb7yOaR5O
0tDmweSf9ptV+iCqB/7sCfF3Up8joQ9r4GnkJDwT15ENpi2DCyqkjf06siJzCZLxC0gHSOkkX0gM
AD3OpgxNm2gOCAG7GMEREynN1NT2uucTKwjiCwRQmnkt1+TLsnoLbxArGlDqy9iIQDwxlVmhN5Cj
I/hE/hT0/E41/TFh8ZD3X625XsP+O4nGr5qqhK9ET2vO6QB0YleyFEpjbAlnw+Gce3u8pQwFr7lY
JGfpNgg3eSfa53XF8Q16VwUeZ9meeRDodmRgj2FlfH0tOX57uIX+FGuM1FthdPDopKMrBvU1DJe0
dvbR3FQTbKj5ZtandVsrJ43roGFhEXzfUziWajYN+PlMcvBoHd2ibQ+jeRJNF60rkCOYZvwZSPUy
UzZgHPILlMUJoGtcheo8LQDqtbLXgDmjJOHeaRffGC5IcaqUYOPBAAd9kB+X2yxaRnma1EVqATO1
M5B9FEsIWaS/2JndjSw5bSVwsMQa8JEtqPFQ8K9McPGmcm3TTFRKuuJ1DYP1w/kw1m5wSeoZRfV2
cB21O9rovlEvgb/svukbzwoyAuvMsPKaAvZ5E7gWKb8CKoy3L5OafbBZ1eWmAHr4iCd/zk7jQbgY
KVIaO2qdjqXm9Klj4RsUcOATel8mGAbXIy8KWyYJ/6IfN6TX4LitJPcIt0kwIFMqx4fJTHzdlte0
fZTVXWQ72OLyiM6W/qCuDvJJvoclFgJqahgvnUGIS/P6Rqqn7pOwGRlyYCivEDYbgmVQnP6wdTEL
2qVeTFgPfSDzpzOmx7J+2baUUNWZPfbsVsLgFKul+3m+CMZF3a6MdL2j0N7Z7vCYyCy0t/YKW6tt
htTDJ7CWktwqFivP2UyRv4CtERIH94kHzsYiOk7wdEuvBM5uOxREK6iVN4qL8n4g5zEbkoesKPZz
OesXe66Pah8AYrjvqvhAm4tFJaNaXdUqkivRjW4Odo0En4fyEQdzU6RVe2KL3SABoK+uu53U68qy
8RVSeFMs0oTa4KareOiHd4jQZeYNGqWHxE60FIlfVzehjNiBEOUpm/qHurEjwOUk+yqjubSMYJBJ
bKrfnRe9uuLxa36SqIqx3TlPcjcwxfdaqlzBqbWrObM6XRv6JX8nwrBnbDdempAOtl5xUUUxqxMP
c/rPw5Sm8PyuMoJ2Poy84yC2K6l2Z3g8bL72yM1UIz8hb2LKQ33gXxbPAoaaImzkCKD2c2bZKGwN
Lb0I3LqzMsR+h3qbGSl6nmygdrhlzbFOAESLCPuCBI5NKZlbUcejAak8iHI7KwqrD8r867HWtqDl
jwzX14cdg8hQ0cMk1rjd4t1nPLLO+5m59kVKHiM5v2/8xer1Hj4sLDlgDNvt/p8U/oBAy4Mgtzc1
aY+KBhEaXnt4TwQqJqE8ooYb5nk02a6lArZWwNYcyeqQWIWpdwniAK55gHExiCnbCirLiEvQvZj6
5hpNeaZTEZDWlduajgMk66Auih0vAn4qDIjDzv1nr+obpCQXRsnk2WULGaZmI7UeS7j5oMwVPh9i
iWKScwBDoaf+XzxaShTrP72PlaYW49bGYO9RJ7HANevTnjYmVWqr9fTpDreAW8uqV4eprVCy4YdP
575O0Sb68cDTLvOoi6yDvC2RCEkQs7+CxTVW5k+ga+FUd7TaOFfU24E0SH5SEW2wewAQhpdcI4yR
Pxve/XH9fof5Oa36wxXcTAzR5N37AFa9ZTW+LdXCudoXVKTJiZ8r+7Yz048Qv0ITK1SrJhroc3IU
S3/8bGpLG/DvPMBcftfc0Oorp1NBF2PwWHIkDu65ejVtbbf0SWUI4nITMx2yYqyiP24tEspQd3OZ
11y6s9zLMHlbLgx1ywhtQ6F4yQRpleK8lvEU3SmMPmKksbdooL78PwkmDGwJXKBrEzr6BL7hd8mE
hRXfaW5s5UkdMKNciMtcTZvTZeRK+cBt12KE7yNCLfKnZdfg5j721AhBp4fcfzkc3s/PW4vFGNAC
2dco7udZu85buzb3LEmY6uCRrqDjyJ9+sAkNFVJN42imuGN82kQsF5d7Z6h7YIbYm6mQ3DxFZ/QL
+IiMIFxUqOOyku6JMffm/RSMJ1iUTrqaEH/GmLyoVOcTzbLYN1gLlWnetTms5q1GpUhFwaXJY8Jq
20l2y65wn1PjjdHhGRkNAD9dNWZTOzqFo+onP8gBZirgqQ2PNyvuvmmtDYYlr6cLQZSLhmjauI8f
aoaE8E3m9ArJbEShvELUPPRwvztWj0C20RQaVXS45fb1qFR7W2oKezAWfIfDdbB9Q92rxvKmjI5h
+dsrK8TZ8sZiu75wpebUeDF4/2fXdhluZy8PI/uY66DXGRbRcLcdPnD866RKTteOzhw0/7O6nBdA
ks3Zo84Ic/VuoZXMPRkJb56K5pDrjn+AetQks/Bq2qRBeuWPLiCOQSzFebzcDh7IT1A1feRnGLIk
GiKIKB5amIB3NTKXFy2+YkXwCthTuFscMy8JAGTIt4QWDTRnpm5YWC5DEBqC2uvdz91T0+PqDbUK
0LOD2AkbxNc+qZ+hLEEyED6L36Zy67vXk8cAP/Q6C7UGibRMUeoSg7MNvAgNmT4fQnnDPfjfyYu9
nX0HWyUdNowhZyhN5u5oNr1BkgI7nutQaL6upKV+UxHQjZ+tKuaX83FNL1Cp1vp6avEK9et9ZxR5
N5cC42hgwFebpYAtNLXmOeWkNDqO7uF2Qs/1gzceRZIBdh513AkNea00dcuLIbz9ZQUIQlJ5oYAQ
3GkbbmJB+ciQA+VmFlIxK7MepGSIXem7srUUSQ+sUKvcSB5SeaFgr6fczkzDVrXd0HvzcJlc50xH
toXRl183a6XiJ+tZbaho8ab/6u1jJaiT+KW8h2Vlc4rHFMHvztxrzzsZ/c8StkVmU/KxSbcoIrog
bdsB5GhypqBXu68o89AC/DjAur0ndseB4efBxlQGKG+x/iulGxf475CvPTg0lvmcVJT5tzfMqFKn
7UphuRUlFAMj2/5PoMynzaWymw2mnSDI6NlPUDI8RTfoV/Plm9QhNKXAc6QWjfFU0aG3KT05Vt7C
dks8r0ZpQKtRwVImTdQF6e3W5I8qNo5EG1S3DqHKIVtwUxt//iAvJGINrzpQwlcTXvrCGVqmEBLA
bPTQQP4/g+SKSmDJLZp6TArHGkx3OMsT6yYKAm61oDM+ZkhmRBDjiY2Q7216gDOdd5DW9DHbeiuf
4/Nw1u7cST9LRsI+9ZUtFNRb4j+np1mhsaTm8GtoYH8gBCR1FuHJVh/ay1wQ1q7bhbCVnclX0sM6
vYjd5yx/0snZQzSEE0Ux1ckeuxm6KjrHokbTSDL1Gioc/Ou3M/zW20GvIKqrzQ0R7AUAapjSK5T1
O5ZPnAbtineRyvnxbx6CUdccezA5J2kURspQQfW+XPQZSwYkjU3WTC9VUkzCJH7Q+J/Tc+oUD/Ix
NUj74eDJ+TlGPwi5zpF67XQpnXe+cMB04+6ESTpW5b5bPgvhihKnv/qJi8/ap2VHpDBoLSIL4uKH
3hafeWX/jOky3ZNRirMTBgoy6uRTlN1fiPv80UmIrgKX68SZ52mxHxP1A2q5xdeyD29k3P1bX4f2
p6Xc8xQkzULXVthq0HcQ9iXm14mHflbubxhzenbBmHNy7FIHCW/JWH6lpxbnQTR1gpBaqQKqRWiq
4KQUC5gzVE3PrUC3DzeWz2VLyrZfPn7lR432iDzM7TK8QPNiOl8Z3HJ/+YjPk64VqfKLT4sBoH6/
ARdyTAAeGlYYynLkXYdFzodUzpD9dHjl653aftwVh3FR7SfWkYoBnrg4b6s7z4YCp1dcYLwqMZOl
dGLLghTTg2VgvAiFUmD//P1/xmyf/5nnLcUjHLsSV/v2Tb7qZEIT+a9z5VhpsVNH9Gr/KIIV7K+k
/hFfP/LnrpwaeKmS5n7WgoidBu3L9AROnAJ/If0QlW1GIlCDMJyioO/amBs6OSnwI2uVm3Mgz3uo
25jk40gy2r6gv05PWWP5bctwjQAbyunykEV9xVCaiYvNXcv05IICeiJHjP4bPWdMEn0wzpeVQQih
KZXHTERn9YQFv7cWZ8iPHf2v6nF0eefRiwZAIIzWtw0NFyxV5aDfOnUo+X9jPkhqS4ivfCcR+lWd
0fR3hc5Lj19zyidn1PDzqvvfwTOuDujId6GusXAJWnwAlCOsboEqf7uYqaqHuiE0s/zgg3372ViV
6cGzsTMNPXmMlf0HzUQ+wm7/s8r/+doxuLFZz2/Lj6UjNt5EpbG9UkcTorS2wknyBXwdr4Bze4MQ
sSHLWssONUUaw2XX4x9vLNhxpoVorNE3yjQ0/9vjRRGTXlWh87JOVTYj/e8GqZPzksD4EE34i7+B
WoHNE0eigJYcbAF8bBS83WubLziLyLqtmULKgRWb83LsAFo19Cp/h39jGaCOG7h0vxaAJbNN60SK
MDCd3H0BgBlB5Ms0UdYml306yGQjChPUquSER3sexWT6IuehUfoeLy3dirO26OZICyBVo2uRfH9X
GHN3xU+4OUjmmGABAH0epBtThoyaJhSuiQ3o8LYPM/b5SS525OloArCTk7WB+9//82i1juTBozeR
jc6jecaHmhpR+lFgHqCHWSFxEgs3O5EY8mT/JWv/4LYQ7GmQ1dSfo5kniUE4UsMeYJ7nuWWH5fIE
5uAhhc+ilyhf29qVJEmEZkKoxzUDMAZrV4S1R6/AjRgoQxJ2X98UWc/W0MQTC3DRfsum/C80I2AM
MsTO79tSRNqyv2vCn5BLQ9eghAPQrvi5CzZvtktfyrbjorssbxELLjJ9AuxobTo1dP45gLJk1YZb
umgC0ITRP/ZyRADqbtZzS1HsTeCwyIFJuYDPXmYvxQegUpZdeDLMaEqduTwZ3NP7KFQ5gAQw75fh
X3zNNkIVLHOqSPHR0AeB9aJRbav+K4cuBfpATA7/hEurXekouoihi75GWgHJEumQdOMZyc9sBmah
yeLwiQS2MUFvF5Qfe4f+TxGZxdeBd2OibjcSiwUz+ku7pIwQBW4Epa5F6HGM6YARWrsaTEBKDUdR
LkG/I7TkPVd8qwbJSzo+0tY+HaCpJ/L8rpyB1eiHc5m6XwJ7VLMjZWhN2gUqhqAny6sj5JR0OWST
0mOTusAH9ZUWt5Tnh7eTgWALFSDPj61MRuDiqnqShMAw2YZXP+qvBB4h+57uydFhfrktkRIJ8HbV
H9lrehfdlSWypAdeFqWCO3e5MQ5LHDDz3utbEXiIqk//2oy/VS1w1W/6/j9o9BJjLQ7THIAYEW+n
jlGpu2EF1QS0FwODQyxQVBz3J9GkNjrFFh9kQaQeppUenVBYRQtZp8KwjKHKPhGqANLPITl1tv46
EJuHCJehhDR5jGre50/F6s6rpptSLa/GIS9S2jZfteqEAmd3huP2rwIdkmny3UYrz0AhkwED14eN
YZECbx+m1c0Th7WW9diFPyIeWJcWX/w53tZjb4HxpCh0WQPd9RQTFb40L3SvpI/jy6C9/HvSvlim
aPcPHzGxXw6suDCEJ347vjuJagG8MUnOUAes91NbDAfL7fJcnQ48sD91vP2429fkbwOTmdKsjvQ7
nvcdFOV4f0W+djkES77VDRjb88+vTkyiBgNjia2fAS6HX/lmGmKPJyjgwxaxS2wOByMDS/SS3KI9
sEDXtBBzSHi+G3XRKGOqHiZ7dRs8b8qPJe8SSod6fHcrEIeTHizry2mH5aFEobWcM45xs5/nAMUe
GoW7gxXOKqyT9/LfA7xiV0OXKdfZ+M8tj3GM+q9ppLyfwI4o80qMLkjaMiW6BWl4ZICg0HjWePFi
DJG1ZpNe4UTxzrXMsZ6M6hlDUW/t2VEo4bdj7z3NcVGk/6c5dr726quTr4TWoNkDP2Xdygf+KCMZ
vHZzw/EmeK48Bz+6+QE1LN69QSJgdFZBZK+Jw84bIqXRGG2Hu44EDSeUvhl5p2/Cq4Sf5gJd3DKw
LWlcxBCIkwGCbL8EiP5HIgt0umV13XUpKEgq/xO3z2qiO5aYNY6UH1/5doVl29KuZ/Ut5faEbU8w
vlMkwNBj9s12irt1hPm4ajwMtvJdPT3SshvFOMv7dfC4vfLAi8jU8a6EEA4DCiAe/3/ZjOjsu//h
mlHpytEfpWEqVBXNeWXLPSpYlfCpnlzzmTEsYJkKwe/qDvqdkEZoEst9IUkVFsoG8764d73+73bm
QmTRGAy0C4nRlO7vaLApN5CiuXf/tkbf6PAPiCQYq0eyr7op4lvhuu0QkJ8gxzisWYQuE81dN1EG
Inz+znKCvOGOi6KgolRwtXpi7T/JmAwUy7XVhxfMV4G3QhAXzBgvjP9Se2nrSU5OKduLbZyOrxKq
Jmg7OUD8aXD26trd8N0vgFB7DXU7ijdYhHEIpa2PiBdn87V4P5wuwWU0haa+NYlgxfB7xy6xY1Qb
+ATeoS8S/sZ76q6Wt9pAI6vZ9x02mDzEue+3BgzbdLHOJiZO2TSCE/aKH3GDegU5An5fvNkNGi4q
mQLpWan8em2VH6xhn3965UxtiZIZp1HXM+pzHbzDZdcmzXGqfzR8CeaJkCKBfga4JPoI4ModrbaG
KVsI1bbAp35Cy3LAM5z+zUCbKv4xqgjI5kK33zTgqqSL1nX2oyI+cuCuyTyufvvmL0Z3HbYiWhju
87/H6beS3aVT2mioixn2zAlUfhdgsab/Z4fgA89ZSdPdLIp/SPvrAkkvRH3qP08Y7VebUNrvHDky
PVRLZBdg4J5jolh2gcEWLlAWPJh5GUxzOQ2r/uSYKcDjrw+unPbVq+R4qTNmkzAB2nttYjsqxysJ
oDWOxUOr4Db7Vtb8HnZ3HmzgSS59PJ8XdirDg592aiCBn0bkPzThYFcqNocivrkPlCwC+8y1d37e
ST+fName7Afp8Pg1y5H1Zh/uXD0c+d6Zo1cSe5V37rYEWwb88eJJMHvlXKt+fxeyvko5L0hzJ7ks
LtyEQJbeee0NOxeSe9vA/UTd2QQrPZSK0CzREo/mEnbvhI+XTESxkWRopapHTIsxb8t8lTKaXphU
v+mbdo9J6L2IgRAuneFXtjMQgkywnby3oj+rW8Qkivc42ejQ1ZAcFlWXq9v89+33wS4cow8OpSmR
RI7HlfImGDHI4oM/p24HVDPqfS2p3XBwiTaP594QifrDFGCs/pYK2Ub9oK51cghnWe3wrP6Qh3CN
TZdT8jhA+JV6ibgdyaQ88Yy2spYSVtmDw6HxkyUDI0Oq44ZuhG+Bn6yhn6loiA2bU1Cs0ion/7pc
QGwOmDbeiHhShoq1QYYTxCmwxRMXRrn9ZdAhXl5vCUcEpUZGroy6ENUs7RelTj0q+Q8Kl1BzegNI
DQDZpzEhC1nf2QUl7OL1QamuLdy7ej4n0JkwhNvaN5ezRdg5A8q2DgK/MDJgQm+qeeGgM9nmvjz/
IjPbLckdmQEOA71Z7w9mozKp+3LsH02rEasbROzmRje92i7h4EZcZQ2MZ4xEnzhshMnAzbGBkAV0
ozA5w4zrgkikoTRo0W6mt1MuhKC7mfH+dEzkQeJCyprqF1Qb1Ies0ejlvzEknx+5mjL0EQpR5X9p
meeK+7JoI/PP00et5cvASqIFFP1ghqKQcfMeeDJ6nB6KPbIstew4OlYK+zZaefPMyQW5oTBGZxpS
cvf8BlNZkrFmwQPjqmEAIdiqdCjqLco9GaY/emfEQGvFMyyhaZVEEXjI+xrBd2DsACNKZpmbvGrm
/2IXXsg7GxQSJIUv2Vzksc/up3Q6DrKD7YJttis15VFZH7GL1puYYdTfDLadfa5FlaakT1lTF5Pl
t7ZQG9izkm9ztANihaGRKgWHGGyG6UGYNLWt/ORTg/L7GsAwnjMPmRIpx0Y0GgNT1ZLDFP0v5PPc
Uh5hbuOFXdA23ueEOyX1Cu2eZs9QcJOZSH7tJsi1fCNWtlIr0HafHNJ5orHtxJSENavuTscfQVbQ
iZOtRqASklRnpII0NUz6/xasIo4E+EcIy5FY4jfjp4MmYsTq0Wb7D1jAN2zCgAJNbO4EUHfs9I0v
GhgrsXpvTuVsiy0LqyViuGOupVZGje4SNpml80PowQiTm37ilDNDsa19xMq4QoPPiKdl7l0pcRA0
kfsKEn0FPMcDgaaH10LnnRfKbB/6utrNpCBxwFzBEhNHDlxGry2aNEUT1qQLPjhGOWzqC7rMpsPO
cut48J8Q8jeHo5GMY2D4NpXOsuNHp6gES1Z2CO25KP0tfT+uq1OqqKPuObdY4H2ZvmtiFCOU1ffZ
de8u0xDV87AYNdj6R+4wIBnh0jWG96ME5aYboLlVwmlSf6mv95S3pAExrogKovgrTl/Zwu37SYGW
k5vmG/X/VU4OuFgI0ggTEhbGAWsBwSjQtWPO///Ko3fY4AtqPchjp6sQmHl4ykR/S9i6sYudhJ7Z
iNQpYCeuGm86A3zfcjud9vuQ87ZJacTXObywTd6fPxi4hDY1DeDcYfupw2pzvxvX1vxPfUkps1LQ
1snqDAscRcoOCpJEK4cn/Z7o82Cene62vp9fWtQYbM8lY9edAMBboKUZbFyFUj++ur5JMGZZbiyk
lu/1i+oUlwMRG6VqMoREOYQ+ru/GI1XME/c8BEyO1dNwv1JfnfiL39hxNSDdGd7s2Dmwr6Oabgo8
CoSJlDOjA6v0V29ON1DEKlgbTctfmgNqkOEH1GXORfGANJ2luRSzHnJyTNxLSAPfrCxE0mxJk9w6
ClL+bWOQVV/xu1eO2zbIVfYUxwr4Uw/t7lzuFqn3pZKBXhRCg+qmv0pkndh0wvX1X0+iA5Cq7MTU
o42OPHjK39sJHdkysCl1XXGKXny2AKFfFjU1/W1BTlTRml6LzB810qTNOR+TNaWTdZbtddnTdSK1
QRp2i9oQ7QTfKK2cA8Hkqv0bs43Hj5QiKNNa4PBN0uUTb52KUOcAg6oRef0Zmf67TffIt7cRlGAJ
oRtGA+uIdRqNYM9wjHvZ6774CNzXBSSnkjtPvFJVFke1UrhWvOQ7LZLcSn5djjv5qEJx/mO4SzIV
iysukK6uzI8comKDVnfuFL1qvJNQFAWCHikLlP2uc9UMdxiBZbVyVRxIgJK9odxc7sQxCK/keAcO
omqLUm3TfpsXlEI6PjAkxQVQfRaDrOHkYS+u8QFJO/rB9gggwBdmnpIay7Tq14pcZZrpKQjXtR3H
ySqAQOXxzYfXP4fPaY0CjVL5bgfu97BqyVCHqaWMJqoK8M9INRh1JDkdTIhj/DrwJoOsbLmkcnWL
OrRXs28XHO17h1otGo/YuqtC8ORYkEKKQ9z1arkH4jBoRSGNCwRRcspBf+JoL3vj1KflMtGrgny7
typ+ow526JboiwZeTkxFOZ1vtjsOfBLiIk5OC2oV/pldKWhNN8TKE3A36j6ST4uRcbui2s4Eg3i9
lehaQer5cr5erYmaiGDGyEnEi3H/gw8pYJzdWQ2654upHBxnpa5ZWLfwcoU76SmPGJw8j5M2qsMn
cmYIbuvhgsO1RtHi8vYpa3b0/nUy92L1kIj70ajL0Wf2KXd+oxLGAMieWXldB3x6jGoaFUYiPpoD
Q2c5xeHZQwWV5xO1hqLQfEnlHv2o+UW+TRZDKK+GAVLmifJyzpOd1bHnY4kuYtZowZjZafGhU0UW
3lyVrXZu+idG2emurlKD+4U5GyAHZyyqG+tUzQ0Jk2L/YntKGroKD5KyC/X9MnOTC42WObLey1H8
grfJ53Kba74ebH/k1pmC4O8eZwJNh/MXLXrrd/UNHoqATJltpCQfXZRMnoTkpdY8IaV66yjnYjM9
3DQopdWcpluaYFGzt8pQqvscaGjPrnI5oAxaZHQKneBKdnk8Wl9bNT0W5FkOwzPlnZJVyaK3KJel
Ew+bns0jssZ4k9buLEyRGSQRo9RfqpXPzW8bQbpVkCOHV6At4vKM0Cw10RfjnErwQoVZRU/o6sux
sm354XiK2c8LZfDCcDupWPUACtXjNWgNUpCxBJnWDa0LOuOlsOx6fpC3cbpvZwTRqYcAfBgFkpNe
ViLtewaTW0UavaqAd9V1Fas1IfnKLhBhSdv7VnUUJtrhmzitcEvxjdiWiFj+w59dp6DkByve0Foc
6e/FmdiE0Vhpr2CjiCYs3r3w+rj0Lufwfow0+3EC3q+TXyVAdL4ePDm9aNVzqGr1wgnNH2ugXmI4
HHhHeoI9vERReGffN2i3HDqlB+LX/9+nf6iwOqrw6dtWtMSRPKp4vXPa7XKsCCqyS97cqp5fOK46
ezW16hEzDQSAzw3QqrTcMfsY8YJM6buubFuErtTVhDNaVnUFtu5psyUgEGQlj6XyCZpurgWbXFwD
Bgxh7EvG3RF0EpyOSpCbVePPgFo2TeIAz6AbqV8mlsWrbZZR/ZJHK+CSaK6QW94On8I3282wJfrV
QgNcyRiKcOOLSM/B4pUT1xl7H4lCO3HXzD7HO6lmFjsJE+M86jPh8zwr9BEH6Jbs72DuYG56369u
uMxIceBktBNdOR95kS0EZUpAsy5w7HX81jjIVZXBSPUam0dE3gCOr+7vnQT8/Te6w3zet6ISPOqK
BF6Arq8ksLkVZHLhKCFFO+JWm7gfzCeMe/HXJFmB3KiFNw12x11ahO6PG49UJr4cYvVgJoO61AsD
EHsEajobITgbAZt7SG6NmqHK4qO4nfnIaIZajSmc0fgw76OrThZA6HRq5RvTkMjKX3zHzb3VUSIY
onPLmGSq77nYgiGBEbitO19d+Ah6QSqtrsn1eU6tTqw8JlTSbSflIREIqi8/GhPbqfJiS/HooqVo
sjf/bKYuRmZT5imFVhCEvioCmFfwVOHaTGfnaHKz8/KF72I06XFomL6EGIq4nID9kfZo1K4w7GZN
nBaRjqDHpU5EIRh/0DBiozZzSrQE8nmKkSkt2c2LKRHw2ucpB2UAYf5w3L9iLxu+rviBsgAOfXRN
ElAr6CNwUOe4p2KTci2B656Dk0PMSGIzRFGXBvxXzp/6Rjh1x2fDzBtTJCbuHAVsW5AgdovZutUB
veapblqgjoY7zvyFWeRftsH6JifAXWTXgoWJspk9p9edK7XTef5pbmj6x67IfIPVKPUwU7wnSXBQ
XlFZt77eXb+nLGt3jbo0luyU5UEuyK12FkDHTM2r8WyFY38Dv1NX/kUQSwBTaHD+aBZ7zqq5HFAX
CYx3wCX7Tsztt27jxLje5NDPTfWE3ohVGD+Hd9FPGNxnJ2YuiPVXNZf03FrnPmZO4RhyxRzVp6lz
IMHLdUSncgkDqRyx/zKZCoxDIRjVvp5niV9KJcxtGpsIpoNAjFwKXk+z2wZ+Z/nNfole8vL+9OkC
z+897LwWcsuiDdfCftRO+UqwViSeykseaNKGG4ygFSJdjRoC7oZAgmFvn1U+asnh2viHiVOFxp5s
L93RMLVN0mvmixE6ncPrGSSDhEkpqzsBVdESEAs6XqQGzMCkcW0FliqIxNeUTNCp0kY21Jj2wCbh
aAvWeklNu8c4UwyrNIGt3KWNXesFRbOQs6RAUB5MfTPokbBV4ZkAEfkE4J/693RE8Bg7pQcnJNV3
hMXpcOwNZ2P7sqcB6Yq2uhbwwda/rittNPDlMx6wMLwPbw3yfUMVaqwC26HOGV6NDGmmtgw8LLb8
cRFnDzerM4CFzNwzt/DNaztCiu83/5NDESmEnwMRsPSSJOo18oT7AE+VKpGJJrnrQaH2F546vu/t
ME/0ct7MNrKgZ+CwE0auPuWp+Lkn7ljkuk12NOOmXMPBjyaCWQsmDtEN7vdLbIw2tjtD5+QwnAVs
9VdHdztQQ9o6SNxnc/SDaDXEUQA7JxIw4E6vRBzf5Y45Ux6akJDZ7y54zA/GLeDoFnmtE9x5RVSR
MTrBhqExNnno96NaMCAsaqqAt0XNmYVVqyyofrpeFOH3oSHJSxrpOlfI2BaCVOLcUuIJToFD5Yf5
ajgR8JNADPLRSuje3ZOL54mDwR6fLjvJU8+9CvL9ays2KgLYyJ/P/MmM55UXaPK9AkqzMGxF4yGH
aARaGIjOMUpYF/Q2dK4VdQpNIxDuS9aAPU3Pq3MuL0Wn2be/mS5qDYG/6yGjBqTm/ujt3kc5ZKDi
K52PzziHA5348t70Uf4vNoY5VGf2xRkTk/MltesBi8Kj+hl5/ynrXw7GscmFAz/i/CUU69rwCVP9
N/hMqY0xCKQ7kT8RdNqdkOHwTrA1CpWGRoh6eSxzpF3Uv8wF7jn7xkGnK7UM6KtN+y2cEvp5wMdK
jGn+B9LlKJdiicPUlHV20pwzjcuumfnovxdaXDhjzG3fLgFeeTv3l/s4sMvOS2UGYn6jZhw22L1j
KRh/MiETRVgq7k6zaHsmdCOOm2ivzvXInYjWluYWcVEh93VfxUzlHLDqpENhR/+LywYDef9B2MYT
svg/3kMEQBFUU3WSFJi76iwTRoblQF68BvpHEL0ZlOl6yuX21mws7YgcGq+8KdUeIMwuruocwDI+
B+C3Srhl9vWacOpkWL/KT+gYMups41lNwHZ8Mel+kYaGgw7NPGCLcHzVsxQ17sxttDgYyDeKyfhe
cXTxri1FWTN97WLbWAMRiNu/hfs4paJy1fIeIshoPRs+qmtkKyAFKVFGbj3e5/QpOBQtDlBWD87+
PAMuKsXxDY3hNS5M62yFV7uaLmSDVMS+h5uF9xchSpsl8bZ0h3qW+TDbz4YyumhQEdxqmq+y3SxF
QkSMsXfe/NnHxWeZ0Fc3WlLDPN+dl6xfD3zwabWqlZrWMNXZJF1QdEvqImieI+NXEYFTLPp68wtc
dNu3VNrRpN30rQcX7gADRT3KABgs959Ni04pWoY4nNmCfz8NC9TjgmMbw+/Paij/BYHwDPAkiejb
gurfuSeGYOATUfmNaCi37JB8JpByubUjlkYJ7RazcyYZ5W3E9d252wlw4zfjYXAkDniIG9P5nEeW
kxmZumZVyM7mkiVUhddOAlahv8NrLT0lclBgZh44fn7f6QQElTOz9JUWM4UkLc0Wx7cQFHaFXwJO
OW5/GQANwfTxm7/zXpoY0oFx28nC4nFDXJ1KQWJQKGaLI4ReZmJmDr155W5YCFIEz9B3HeDXpWex
kapj3+XOglFSEdfY8Ggv9lv2EPKC6T9cbBTbcEzw0k2ICq/P17Nybm3snEDqI/l8ZXunai3jLPwW
WEXAm1HGUu0HDIrIIvbHL9tkEVyce6iiY5eDibGx5xMW56LbLJLweKR8xjB9Zi6Z57bvPUf9RKj7
2lu0h/IYxGDlGP6Tcfo2i6zR+uw9Db3giU6ZLqqy68MqoFs8HGOl6G5eLaPyGph1AIgssJDsr3U2
jH/D5uspeTlEYxoVoNJMG0VArmsN0ywihoY5/AclOat2SWI3cqNToO2U9N7tYS9eAK6GNL055yFJ
E5E3lOnfJN8+Zq/iojZLo/yaEc1ed1f2zhPLn1Pmr+OM4CknWqgPMmRO1vFAn7/X78ZAX9mocF/C
OXEflSqfxB9amNlMN7EKXrBA4uYaR6FcwVBBVlbkOgqTTVBEpVzi8hqyKfHPzeaqFvNctRibvycz
QYegH8/Rvyj6wqqHQGftUEKXe7E9H4UDTEnZEzQ3Eznkr6utv/N4vBgpnxZnX5Jbvi5QRkSTvWfr
AjG7MtQdMgLcbeU21xtiFWOS0MgI6TDsYAN7ujzUJfq33s6BzoxIQpS4+ePW7VRvty8QcdluEwfM
OxR4AGluJ3fva+FrP6kxHl/HZ0x7ZtvPJOhLwq8vByuZ7K6bli10mty1Tvf1tD0w6lFtV05CCt1e
L1cItuxCoBcUSo5AaxX4DcHWhvcpbcirDvXuQ1gq9WMVJaDmrL2L1HPMjl3HYbgcifOEPzD4aaEQ
YbV9YgASCAgHrF1ErAjXW9UyIp4197hVNGmZ6B0S0mge3s35noiD8aYrVlGuulQZEyK2ESrX5FCn
85uLgu9VyHKnnlw716zEjCSykPmhr8cy7hHeiPTY/JNk3lXqZD5ItWHd5sZOuE3vGA/DJQtsoEfv
+gz0JBMMKYNnqCmtlBe0op5kfYSq/i7MTUGT+2lytABjqKCOZ7J446snomIUFjayRg5zzjuksluy
Rhqn7nDeqseNIvyeijiEi/Acp4cpeBI5n5bJfghVhyOBKpGRcHMGfetTdPHhUI+wYfvtVi2voyv4
KgDJrJJ6MTQaTUK3ulJC/EuZ5rZzyY9KuFK+LnNVdkiHFZpFRrCQCnVsqvDYVHcdMwCrGl7YgR8u
+48IGt3aCSoaASvSdAwsrax+l1YaYBJHOVd7gzJFlBtySXsaCB3H8phHrTd6ND+uzEqHK5qvtiPG
PQGvx6mn6LAhkBq6nsQalR+61axcxZpO3s/EhLpQYanRFPvwhxyT54U2LIOOiLlbIiSTrnvof4o7
sOzCD9uoA3TdpDqaychcvTAVSGC3g+mqABNrMWFZXnT5Etmu5y3x+xDKsk4fiZEwR19fTCnu6ZEb
eOxxSwpwQ0nlg/z20ZSyskpIOF95o5kk0fIA6M6DsDUw+2cNO/hwU5OjmdLAM4ofzobRlyHLsUwA
jJ3xm+MkuT0hOzIgri9S4UyrihEI11s6TkOYkPDUzO9ZrDYDXo6sFNfcacSZnHrv2BmsNVIpRIJW
l+wXZKAbidNbmaE4YyRzwFhuJwdrbZSXyxYM0w6jnL2b7J6ln0lN8wl6NgdHkRwvPUjkpSCLt/F1
GVR0T9vHN1D+7CkP4pLD2ylIpQSxrryY1PZ4IB17aKfhl7cY/SNy2BzdMzdIkPY26i3i1/UqU1EI
uWdNEkgXbNLPl0POC1y2fjf7ngWPdwnHpKsouyaXDfFCy+jzs5961ugl9SIJjh2kqjJxtaaNTj+I
BCgnTYChcNZnw/jZixTsRw5NrvYyvehBvL3D4mKkttnTRjRp9bbOmudKrtaeFSu36N4FSYLfuGA7
cFHpOLclIrVGUMeZDRd3BXB7VoRjEcg5GNhjUR8hj3Uoj4WJ8mumbtAiqJZ50QxBKX1V8FX1Tvu8
NfCINfm8t5XPKkOa8kdsnL7Kt5zqNmjWcha4RnITWGIPqytyGm5lHCBv327HkHmjctDkDGnXDcZJ
flBI5KZcZCC4x6gyh3APhPFrkelkNKzzRoDlhrNE22FVBcwFDnQECoUkAY6NEqGfIrcHAZVg6Aa/
fqW1m0hxsIsOiHsebtla9ObQ8CJSq9NhX0EGHSfa2nRB9LSR1Uyf553EjvOtaAmY0+A0Igvu3hhb
eg5u8moqkqwiPaannfBjnLMgHb+r/r0CljkWWWe0inapWrhC908Hre+WagaujeO4r6f/qgj6k1A3
VET7dzW8BYFS6sB71DFUpyCPhXf97kBTEZh4tHivdNa8TR+fQzQ/qjVoHAxMsNhLf9Kw5eJU/J0L
LhkTPK9SKrUBa4F1wiACAd99O+pyDkwpYNZwJc/WnIZ3WAs58KJIwlZWY2VP7azlnAr6xdMSPZvG
SP1LxySgEeoZn5tKDdFZt0Am/VbK0hnyoe6mI+jiqtoZUob4EsqWWuqnDKtR4f4ZUoZCW+6jfg1v
9Ft7MjG4Gd4RRDB1fJZknliOpFJQYjYKhzvyMOq/h190xdrOgZPS1Eu56qi+Oq9vRfo/GT6QA4Qr
yDwVGdRih3nNr+8THd0TTrv0UBjxNE/ehxaEUCWrHWYr9qIljbADVYipekptLmeZK2d8GblIIpc1
upbLMln7VbJFksB41qPguBr+osmmO9fbiLqGiD61k64oPfvb9yzJGrxu1PEINLPXOGWsHPA3jW9p
Xfu4L/F69BPPjHuhDp2cRMsy4Xz8Gzm/b5/AaOfUmLre7FgKrQ2VLeb8AVqj5HJgcTdjLK/W/GAn
nKWQIg20yDHPAn1frj+VnWpK/2ShuurZxHd/NrjGBEFIvn132oNbrvndywbxtIOCohykwl9amuQm
6cPJZWgpx0dhjiFotNThz03P+wVpuKcfcflpBRXAAjf2hbZ9eGWMaN3AdyD73zeDPmkTqOIkpxOt
C3Sc84KXQEIJ1CHyKK0IC1m/JCZ/IANjGpMj1aPOH9nRcPNlrqpB5t+YJocnqNTHjMWHdpuXiKyt
KvISG/D6mOM2QK3h+3jBgLQQavNuOrN3vhq3XizrCc44/ZJ5PH4XYZ6NQ17Wx5BqfaJcVRWGA9Dw
jUr7cMAve1rifJKlz6C729Xv8e1/Fa70D0+AG1/7/OJw7Rv7zh0hseYC5OnGbm7Uduylj/KMw67F
yYMahFWl1Vl0FEzQ91tauajXzlrHa4EQNBX5joIyEuuKEl743A50qrNJeKjKb0OOC9lDXih+XCmN
JYHFaLmXosgvXjPPqIrnsPPNZFNPB0cd+6HVTONsNkD2ibEpo/eV54m3Wy2ELT+za+4J04e/wKy1
rYI57MWxugMuEMBMtsJKRM/NsRYX0Vct96JcVZssLvJvJqPkNDmL37rShMem3qgP8+ee4vhUuEoI
cwBwzQIb7J9snalo+Nf/tSIfjcdEUhg5NNFAG7QhO7UYtn9m1k3bEsp7tNcf5GW1hgCntzh94xZI
fNn51fRmQ9giPkp+3CcS2ZMgL9xvuGXnkQzlqdPmGIzu2axVwJZDfMEZ6lKbCiQ1Kf3Owq+Z258U
/geOaOZ8k6xeH2Q1/X8z5LBG618rEKpgPtN0c4CGsZmt1WQMi4XzzyQtixsLsgLXXOTCqO4fPDd+
QU53QxzpULo8+wCUGWOgTkyKXzIzcc8AcH45QusE6G42M5oSawEWJ8yVm3mgG0Hs715Qn/cNB1tL
PAgih2H5zM6SYaf2ghW5LXyjtJB5HyBpCYDaU5JXuZObRHWBqAS8DRskHv4RKqvmaq1XKwzWITvG
D9Wc0gD729oXGGFpOL+AFBXRjhEP7KcEn63ZqklK+9jTvfnK6vn6PF7HUN9sRjxEa+gFV09DEyNp
DKhqtLaehjkYzirdOI9aqXUjt3F5PMqcJnoZ4eg3vUChuHRiv8ft9XPqixJ1Ymx/FqoKZIkRWMBP
by7Jl5R2QNRu/MLzqgWPa1/sIDZGZ6VKXRZUsKxFkLaWElFS/sB1U//aqSYZbAaYnLIJG8Vn58SK
KU0xWvLPH85lK+8SORpEEa/kwxgeuco/LIYPkeNjv0Mi128Qm9d9EE29nyngi/pKlH5WoYGQVlSg
6piH3MS75A1xl33Bz6ywYMZPLU36ENn0bzh8GyJqPsqlRs5rkS+aHh7PzxlLdpEGaTqOEBasiidu
NTjI2elRkJ49lWLOcPl2sIksUV5mQOhMb5Am6JZNWA1RILJhjwBp5g+3pmHZauo7sGzsfRRheLKn
ziiyo9+n11j99cJAFeERYGwkMuLgVMcVYH5sxb5Sk485+pGvKlIyZ+zhDvRAEucrARr78h2Jp4VJ
p3df1P6DXY7rVGtDuR4jm4UwSqVaioHx2LvBsVpzzT40V3e4Q9G98Yc6OnPNsQcMVxC4FbfSdAeq
XvQMb3UkJ397iWVy1OHV9Ok3lwMRl9tYupxdgH4R3DRdsxlX6Qw9wvgQWyQoW1buhYxcL43UlY68
s7NOvlNRhxBrz8YdfqhjiHd/So2VuWaf1E0evu0XXSFfj2L7cVDdI1YovClJneFfFR8AopfPO+F9
NAVfk4ljOplpsIdhEWWfUdZNmSPO9D4V9IeK/VLxy+mGxwFEc+QfLIA4qtC7fYW2rjV0ziZMrwnl
ykGLSQlZcxXow4oYtRzThrHROp/W64k+foCePLEZAfL0j1Pn7glNWcO19f3e1/zDuaUwiB+bD5mB
lk/mbc0HDyHWrpD2GvJW6GaVvo7ShoWfFDCKQMut7EnK9262LhSuvXEw8C9djT9mEVaX7H9TuKtj
vsZIQOcCnCKQye6tsMDoBd+e4IjBKT/i5FRdV4z0RFviTFnRACO41lffyUVTz+NaVf+t9EJL1f6j
uaT8GlY8pTJUXzV1v+4jIRj+Xl7RmDzvkxNAd3j+uoe6Yx75xBSZQAV1q72wBdNIZ98t+R0YWqEd
RDWNNc1SB7LeitH2L+at8hgsQPdJDh4G7TqzfR2gfKSeVJci4FdeuXg4hEevC9Viy/kM0H9aaGAr
3l4vM2y8uJE2/NVgIu2eebTkpCHzOUGk/InEFgF2I1ctSmiqKnptJkp70c201JoAfuQ+GpoWsCgb
wguinWqVxGCbu9EVQ0YEXRXmzjgIQUoKP9np1K+q8JrWTJYgFyolr1NS/peM0KP/Qj7Ee+ncl/jT
p4PiRs+KgcuDX/DzCk+AWoj/oKa7M0d+uNbYPBHYfrzQsujRZWZ7/oGcvFovAWJ9k3bpFIiVjhYB
mBG0FwTW6OxmvcDg4coXUJYVW4DlUYVnIW8H6ApMoeXmncDDCw0lMldgHCwaSNazJBpnV+1ER3/h
CDtJSztg659yF+yvUmfu7VlJgIhJpSuYHRjSzDBmyQUzR7+Se+qXYYNcJznSZHZg1fW56r1wIWA3
0KYaE/j0YcoWJHgJV7ljgwiHAaWHefo3pcNxbyd8DPqW7r4+Jz+uHV+uidJkW3OKDU1oQs8uY6bc
CGptvRcWJ/eDfzfPMSZnS+2lCJ1TV27N0X9qT0hNScUrjLQS6LItws9vAgde3CxabHsFIyV/0ue0
xOeVWY3cT+bfkxzmoY8EwhodkfA9WPjhXdTYqplxViDa+nvL8Eq2j354zg4OKEYI3z11Ochbw9wW
APEPaF3R744RirU/rrfMJU0e4NDUdQe3yoapXddRk0tAy166p4ik1ExRLkRt5yODr9en2M9iyrpd
gvainxIEjvfalGTsGGlLzjdT39SNDA0vA2uZFOYHmxXmRqh6gi9lX+9dDS7hSCXuTPkVo5WSLc5j
Z7oJZ5Rn98ea/8a+UXfgYtHovjA70cWZWVFal4p/gJaL5sc24uj6vB6GUo+mmV/epFkKnSPI4oFx
GlQO2FFdx9KX2mX+Ya9R2jMgcgvkRZ45QK87LXCjld+sOYmtZbWu+/Q+uXd+my4fFhNXYr35t8Yb
Aounpr3jd93M9bDo9Qw0oYAenq1CHZt6nqtp133isjyJ+YPdIRKqZC2tqxOHsa62OaI7uMJPmrmD
8Wb78nN19MZ+DJsgRS/QV/+VeXjOQxA4IqDU+pC+TzHoDKcruigvbU6D/34GNCRdYs3YOEvnDleV
gMqX4QjXjURKOFp4kCctuTS8OVyiwXntm+MIrDN9+aBXJxd8jGf5yGgyQi1rE9lOR3uZAtXlAHqE
fwTnw0aIpOo0RjtiTDxxf23kD2zQZsr3R9us1WxJ2eOOp6ox6cJmLSEvDsp3qQz+flrVszbYl/j0
9mUwYMD57TKKac/4OQ2nr9wCjCDW2fBGwEj2/3r9KDQobP3qEm8OSb36/TDPGReWYtCYp5cv1iwZ
9/gg472Yqxpq5DKFclnoR0+HiPSxqnPJXCj3OcG59UAQ8F/Whi7APyD8PkkiqqVjgktcxdiaDw13
wIdqn4Zc/FgDnD8OKA7B+ezVsXgoq9fhRIrJQD9lvKlxEFIcnmAtKXSK7UD4uIU4UaTEmvDRpAi/
zZWYkSPpHVQB2U9vhyt/iyY3Bov0WfwTilMZxZyyd+/UBjTg6W0XQaWNEpMBwZF4qpYmkbay8IxR
FeTOMsVQTIrKoagPws9r2wwJgMnbnY3275Q2/i55EMZIFD0OsRZrhy15XbUeSaiTvHVzS4WtxD68
skbbwDDdGazgV9nOiQMk4rox6kLo4/XBqvYtLgauhBnU0daKINDlKZFJRB6nYnR5ktgy43R6Q4FB
tgArbO+qda+9ynKi37lqvFdr9A1WJkuofOxwLE/x3XdJFZeu1CO95foWR0IBQIBIBTY7NsssJd55
zG56vCAsY+hbqH6zCryiEPNCzoSFEfyywccy/wrCSKHailrsuNciaXONCwiry1quB3JaUailmuCb
muA7pxn1ut5AVj5q8XMns/s1cQIt4RObo5eZVRKKWOKS/DDAQyPuCNfzJ++zm4KhqBQdpenR7Pex
VVNCUUsOWLuq5tayt5YZuJKmzTwaA66oHeGuyKUjuoPMpooVgyRce2JDsh6cCZTLP19CEF01a2ml
oO2YZLJg3FoVKioRWN0BJ2jyju8mDCguKtFp8PD4xI6Pfht4GYpzjbFUI/numBP8vpXlmApExQvS
Vm43CMAd5R8UHR/TAdTQHvMn7ghNhNmzCzahsJ/IvtG92rtx4nWNhdYW5fqh1TfwAuhjQ++XDy1+
5cO21bU8JuW/BPr1mjXPLgs9Q5QjT3M2PtvHc5cd4lXTTVXfqlXRu7diHqDT9tfcK9CkwLthGHBD
+W6nawhaAVaVPoscG4GsR8CJZ6lQs0byAHtGQXOvUtb1Uh1x3uxTc0Luh7hJuB59Po2+lngImZEB
j3VjDxynUDMOcn7C40I7CJXMSJEPh6ie9kqQryv2b0o4/vFNImCm4wBYZNk4qFxYr2+S7kgTDlPY
hjGE2XBy9qikoDd43AHJLU9yxC8MsXeIrhCa05xJ5/5SqfxhvrXD1uZ+GV+hqk0HM3poNJc9LxD2
yuzlmzNBL36Lu+XX8EiHnhmu4uoxj3NDFUpKYseqHZBUWryCYx7C7auKJfNMBclTJ2RLj0n2+Ttq
IlnAw8+f1ODR0aKBsLLZA2AepyeKIWFNlKGDOLhDZDubQWVzTjAvlK0p/V3OtwtLjGW/8ZxILB3K
4uJfAdd05JZ77c25f68ARxI4eoOC/Mt8ennqRJSGUGDFZeqYdQPPr5G38XitwRBxV2HwVmQeCNVl
FDAKGhwi4aB2CIXp8LWe2VEy6QHx+1ivDnzTew37r77NvHk+yqzYOXU9pr16wwTPdLq5VYbNWnHW
MqUFY42fju4RPoiwSW9j/eVd2EFiwrr7gXZqo6X3PXgNqCNuTCewyROjyTdL9gWmBk6pWl6UeXTG
gk7wEQlnVjgs+4MYwQbIKvXRzUARL85DWU/8KRN4QPpLdOHL4xHkPr/jU7M9jnekOQZ5ogq3RHW6
GVh4JpT8HCeQoELH0CKV7X6yxjEycDoGPS5a2TNv/KnBLQOxOMe0eSvUId4FDcyA4DbDM++aiZvs
oB9eMaZiWFlO7Eeuw1NffuNVcbZAOY/2P3tjxiIkNMk3wY2Htvuasawq3CrKlSs4wbw9FOFEInCM
uCjhNTE6kQZFT1WybLkyCfp0WZZrh2C7NiL74gAQYxWLJpCLOFvjxVnfJnh3icjYG6rY7ILps1R1
yWV8lTX/U4vpqEj7pPs42BHF7wfCFBqPzV1tO4hYuFVkATUKDa6zPSj+AiYlp0atTDgkWQ4QFxhk
42iU/Lr1yeFGjUP0jnDBPRSMZzxEwHUo0pwlrnmnh48N2qnLe6SxUm5zEVrCfeiZmiS9GKGlBe6O
3olFUfEEZKO+rTnrEA4G9CEuhpib5MA1K6zm75t4dYqpeJBOJtYbWJJVK0r+6/p44E+Tptb9PX1A
AUj0i3f+w6trCsaDOkUo4NbtAlVWwUHqvaxbPyEz1sd3IjzUDKKcRc1T4HdQnb6FvXR/YcFttp2r
puWg+h0Wt7K0AEro7YLVmuzr2dX8JfjvatfCdTY18R62qe0O4WtAM/sycPY++aTf+p37f6plMGjd
3aLZ1EcSAV6wxdVeFuv40hfAgQQ1ureI1Ed5ZcBk4V0HQVdliQ0KsnZCFEj6wHqw6IV8GOqFdE34
7eElzqIEH8H7nOtW9orSWnXNJwDfZYsL+fhnmzF93p6fDiyciOner6G7h2Lmn4utJ5IT4ayKK4Ls
M85BA7BEWEhmDevr9l16SMCkQXEqWvO6JsrTWjgbfyUC7rzTlZhQk1EOJLFNrDKWtUCU+rKS0lMV
E5Max8DYtuTDZa1A4pqVpd6BNhmT4G7DlJ1b09UrD35n7wXNs++g3I6YuuFG3ZrlWYX4QcTFpey+
nza+gkBufWvPpG3RFmpC7qL53GCUtgYjdQEchfczBfEhQ8GYYu9v4mtUWY1DeCyJe/g8j+Ruz4ol
uO2gXh57mtpCdMRpIzmARuz30k6Bf6h51FiEzlEg9B0f7kZItPUE/KhFCkcAcZ3a/1PTA2GMsF/e
sHtf5BCBJF+lzOGsiM2MV/XiwQCKj8tNL+g+e067zevO7COqeXUtOb5P8dBZhccudWdw3/Uzwhzp
1uo+LGFpF/6mj7h2DTRxd5/1F3R4Wx5BWfRsA6HfyToCqzhGMwwuI3c7ay8qnNQi5M4K9Gm3icpd
rA8hfFviXsuiBzr0qqMLnf9LSWlMt2XCdt+240sY8nXXn2+To3n/owfJfBEAzNIsWKXDJ46ZSTJ4
k27hgipGPO2vJY5VBtozZ5svscunv10f9OpzWkm2V3JJ5s7jUbzkhDrO0MJy3iNicEgchQHIeyZm
uYI2vRgfaZDlMDSuFLv1awn6S5Kcx8uCDmx0xhygOZLtnXw7zyEDvGYHDXXE8uQx+Mkwgw8csloh
prazdmeNtt/1z/lBQjm87xzOubuNEyiT4dlmkiunN7yeR3Z7Aap1gQ/OeyUeIZtCVte6IBzqfByQ
ZwKUxUDgMU8UWxKbLYvclJAQ3RKDJxn1Ap5IjbpIyB4bzXmutg6ckzRG01dEyd0dgypqLvMCMbfs
7HT+OJjUv9zLv0iPvzl3qcNAZt9X3O+qndq5W0ozvo9g1Uk07wHu7L0Fm41xJ++VfVVmffgtUS0i
OjKP7+k29AV+3N/JrO1LDAxh2283VFcY/zRbuDYMJ7c/1dT3IYCOhiiLXT5MlbPDDa9mv5vUJMUB
W4m1ad1XB9HjnmQXbfsdOnEmp/WZqDnlKcW4qHdLxvsxw+yjTWdtHoTMEN1CvmbHCCY9Wk45lMg1
7dO1B/WZb8D7UGZBJGbI/7VJvTK1T8/bf0xsvqVVMCld8rFnsFQPwp2jsvNJX4iyPMHVqgZYqGy2
TI+QJBHvq/GFHBrC2/vhpohf9lEe/IoX3G5RR6UcPVTtJQRDqSa8SY7Vrwo6nGN2Fi53LAD0AGyQ
6DzEgurLCQ0Fv0OSXutBarddJKdncL58z328MJQoQtnxxQQQX4/hOvAxubXaPgQ05v0VGp9V8lOL
Nt9080Vm6CF8BABcev1iDzxeSRgoG9W+T3dHSE6bsezvdOzDNeAXHPxlgqcx1XWDoQgdXtCb1MjT
C22sRoaCp6nMV7U/B5g2WK3x2aS0+hrEYGaQQ3KOTtzmyKFA8VqFzxVhuT3ZuL8QY3kLljyVDDCZ
ly1Mui2D4eCSLtbRSqOZkjQC/aZ/1yw3rgWDDKqkOWme1R5vX6nlHjG2U8U8obkNIIiuh6t+Gv9h
EX/JKZG7Dk2u4AV0xp0flHiZ7eaIwSfxt5rQyWL9w4secM9PSQWXVrZj7y1ypJekjYVS8ygN95KP
wkjXFF90io1F8AXAOFeHnTItPkZPNZzagWe0BK3ZvBAzGCcUgG1VArNyV562EJIin2VRQn2EKKoG
lDvBaE56PDk2i1sm8D/xjeD/ri9fk04FFNYgbtgSs8p2FpdEfOiCbTfF938dLsjzA9WPiCdQBv1S
110+neNCL+Mmh2S8wSx8zbN2KICDo8U5wvMcnpaLCZ1LDdg3GodABIdN3V7iRZq8kalzbeNgbprE
DZV+IETVm0Ige3dQohUpH3U/ACOawfk5g1YuMpeFgqI6CNB/3jYDbgh25LTPGI6r3Kg7nJ6bhTe1
/S4lLexpyRVFRWWpQ7K0SOqIX8aIo26uMahJMeHcTYe0gy7d83ut2QGb44+M6WHC749hozQKe4I8
sPXgsBr2G8dsZNq4mN2X7WqB0+gx7Vq9aJP24s4CJNcGdK9T86vZ/7NlB6VCtExEkH2PIo7IHbCu
pGeC6KKkBN5ZBlgMUdRZyPq3yNUmS6bToaq5L5i0R6p4bwIwZq5aUUjQJrdtx2ityHfXIFk4nKMW
tsvnPQO2VgONKt6GPtxpTbCmvF/6SlIzVB+ukW53wMmhJCNAwwHbayMSbN9KdxaJVOndX6KPS0pm
WWRVIjiRAkVNp5Dwf6pJJhI8xQZ8DTDRxrENRWKqseQwhCSRgsRkUZFMn/h2cXSoAZrmRGpoayPu
KGvupkofQS57iET080LP/QPyiq0R9y9l4sLZtapvH02Z1NckpEv8eu3mYhsr/yRKnMsEXXK2cJsQ
H5b7Bcsa20BqGlnfsMkYa7DQdyHU4W6JZz313TG84nkdqGMLN9qdaI0rV7JqbADTWRVZPc8Pu/FV
7QyQNBMs/U8f9N5mXzmMFrCdOAADj/pObLWSfHsGkJx/nX0ACUzICdALl0tCe9dZpchVaOWRHX3k
WI2u+0QhMIng75h1YSh12Q42+slmeMDyqNhxWi9Tr5qzTPIuVh6oIG4u5OqvGFo6wigQ6+mjf9lK
QLs16f6DKp2PRMcIpGORwjh6OM06PoQ/tJyRzIfyDZ8Xj4sghKGF4bcakOKHQHLm6YJEF0D6RBn9
87o0KVno5r4FtarILW+hauZqdxKb6zoJg1e+fIvFJCm8VsF2tCFqLjJ0GYwu3mFRDC3lAAwGaMxj
mwHsTjJjkSe7CRFTcezPHCd5c98AHPahC+t6o+qLtM8Z/Kd6+qbOMG68j+EVKoATHrghWu4TqpsO
C8jhMv8l5X5PvlXobNDM79KMkLZq3phSNH+U4H/1hxiaw5VDBXn/BwSDSJE0u4GAwPSctyk/J3EB
vQX9+6I5xwpR+LB/AZZ9w3qtm8D1K4/njslMCa4BBH2zGYLxiIrajlThDMmiQknnlA8ztCfzsNhQ
aMloVzEVQlXhOwuOt4hKVZulk77OcFYBeI/PqT7B/xyjzJNiaUCyL7I5dCZEbdxKkPGhgvvrPzTk
Zh1svOrhj6ef+ueFu4sJt2QDU7BCV3CT/f0ep4JeoKeRuwmRcBdBndBG6jJkw6eufUi+fk3hooHl
U3I4kyWOXSzMqJ/At0JFEFIYEOLGP8EblhNxQ0z64FtD5fJZEFSe8Pwp2gYPxlkRpoujmi5YIME/
+ye1STsGJ5WT3UdmYFEGqtgxfxleeXm4h5Z+FcXGdobt6wy7bwSX+XUwlpJGB2PhtwIbDAe567ct
DzmMqy62gsNwA47f9cjkpYURHHlfC0nOtokVFivzOWyIVs+47hufYLi0WlWlP7AGp0wAavZLIauO
HlpID5ZU7UHcDBPTxnrtI4bB4Bu9FM8Q4WCf3bikV7J6FpmWfY/0sZsf3Aa86H9Z+yBbz9p59Rka
OKSrT2lIPpf7LSzbv5CRyiTfJeGpyZTeveFzBT1k81LDrrHZiZNFEP5shC/VGkcP/s1YxA8A4l10
Payaik3bMuoMatXC3Kjs3vjC9AMkZZ4H6eUcfk4TYqnCmzROvhQPQuZtHTAXJ7dsnPlbZdrX+IAh
0wKZfgDVS/UIP8xXiUAgZfgo89tiCCc54cC8S3//jzPQn4i0C87xLBIBgEwZvhjLtIAaBlEIq7WN
oAtsD280qstRSkXVTnJMedPpw1UDN92uR5VjNAuOnPy1FXiziDlqv1Wa/0cGGe24pyq0BncoJvSb
CcKFq0Cpa5jYAGIbVGsE08jPz+OkfwXwkYFGd8oVE3DdjxH/34pFvvmd9mtILtwli0Rqy2huf5oF
7HEPJ/yVjUJjcLRlvCTSi0qPdMexCLmydDl4E8N15X/bpmCC3+N7cpHZ+mV46C+Ny0OZyzxmYWd6
lawlODIWPZ+/RMZcpLhPuTaAiufKQKeSJL+3vRgxftSz8L7PFjCONgikALL4MDhpyOjfHG4D0LOC
mpAZZkG0kOcoJhKYYrdfuYqG6InZi+Uv56q8lVeghs+1Vlo3YJ2sGD99p17GHPxoq2EvRXoaG81V
U1ef5w4WNsjs8r+jEr1pU90Um1bIY6CHUtwKuHlV3lUhtsW0q3Y+zAQsZqHg1qO4izWxb/0pvKcz
P9fR86MLbaAk2xQ+kNlcLeKgsOGwIYbPVEZoWb48s7VwHNAjM+rDFFZkPhIrPVLj7XKOuQRmKvlU
G56/xCZvpibVvd7eLl4BJIADLgQdi2al91GlkZHWbiUfRpN4jXbGZAjihxN2jb7oxRz/coWSuysr
yOqlPUg/4uIEzf8fvhoTxVXx7DT4NGw57ck659oWLqHHEZFMsgZ7jtjiOsc2Xw292B2EY4zTPkwk
lR2Y4T3YgtPsmxh7kHEyCwidl9XBbzaFIeeR0MXhDwqSon/uauA6vzo/lLF9Ad19YMxixRtPjBm8
Dg5xMydURgv6EP9RDXnxvbRfmkrA8kiWbl50dm2FeClY85Q92H9M8mlmdQeIrFM5Nlk4vnhZTvk0
W/7n39WgVXU+sWGJvTturCJ2hBYsLDbuVHBPw1cvZaLP5GKxUAhtTkE8a5n0orrLYP8BWKXVX9if
TXO0LGACY60Vvmy/rpAo4wcJugGBUiANrB0Rm8Cw7+wNthqlauMgP0hcAA9OTZB6bz3m6o1Vw7sG
N5h94tIPIbZ73cZPHJ1uA3GGQtMNv3PmHjee8Qh70ARgJKj/vQe2rBq/Dd2o4pkQ+W2O1H3WX/u2
xlTqvEbO4OTXvryuU2ilk/5x88Yh8v+Fe0cqvku/qYJuvMd4jJ7/mqhWPXUsyq0ym8ApV9PIDDyG
l8hfgo/xmbb+47chAg/OHzxsQqwGHquZW+7k13Xgjr1YbYcxJ03rccM9Phe5fBaTAYpI1ojubA6z
L2OEg0G/i3dAlKooZx2V437PuoBt85HC+sp8NrVWEeWIX2u4NTZoLsHwazpJt2Vw6GiTobzwPMeE
e22K8AZhMDNhA9LKW3Mx/Vszb0KsF7q/TQvQP6rHOX6FzLVmzUBazbBByTV7z27KItLf1HcKtbto
SM1w+/NoGEzEcvTj14Wxx2sromIuQwkB/TR2DEQp87b0Cf7tzEQFw93rLEdSeNyth6dBlILFGEAn
w0HNi+hVU9fhJkmhIuEoMW9LuZ46t1C3DliZmWqYBDu1X7nmeaNHSjNym/dT1l93Gv3Sj91kAFNp
iLccNLQY6G0nWWFxi/09bWDZobDjxs8M68o8uW0RJyknpGlbwkrlN2WaiK6SINluaGjspHfjGJis
7dOr6fVqEgUAuRbyaTd8ILkn5koiHi/S3z5e3JH1KOtgFxLNpLGM1scTRpFJ/g03m/G4KDv4jz2J
XcV4fh5W7hQEpg572bU4KzMMGlzsv5mnYe1RwoHET4Ycy+4TZUv1fYRhgfVWXpT1+P5xJjCm7uNF
cS/pQm41lWWgRTBdDrYLJyncqW+bF9yNx/W1XKGaCh3US8HozBQmJ0sPKyXfuKAO8naKOlmhH4mz
9qvC7N36BYcy29OpuBTXP1Zqf+UfOHBdsv6EqYxTVdF/edREW98tOSZofzBJpeAN3coRbqFZWuA8
q09w1IhEPPnAgJ/RFiOnFTHaheufVbOTUNRlQmAAaHtFC93qrYk5RwSQZTFoPAqOYZC3chmapVLS
obvs4o7WcdP24riWOslwTYq6HW/QpcBpJTqRnDj2nyqkHOmc9MkJzNJDmN2n0Dztx1BqkMu9RSVE
noKX1SQZI5nkVhhT+fRXY7ic0gyOhkbhy5OtLUIzzCF+8Cs+drmMRFIGueCCPk17BfKLM2zXAz10
rHksoFbcTbaIzXY1ytAlTd/JoDcNiSYf719j+tOxLK2kiaYsI0iw4xQavX9E/AbsPe8B010PAdXo
QGMK10oZBze5K0R36cEGxM8kXDLMHKfDqBT+okFgd0SbljW+5uzF2hj1YWw9HFRvj64egrBIEW12
Hn5/m7U/rWW0OaVLGybV4GoX462Zzu1j6SCKPy8YV6liEI+/XKtkoirkgi4W+iJ9VUhXtvOcd/Eo
kRvwf6L/SJLYgtcTQIhK0sWv3CpqRyt3BX898enD788k3P2dnBkY8Nnb5hBFs0Fp37hxUWpnWhRf
yzNd9sCI4lm0dy4rNE/DERxKkMPC8thcMe596Pgf/EbtVc45LDFdnqAq+uMeRP49VNnb7VSoT0bI
0Q/nyQP4TYgNPsit1hRJO8gmlnXVys85oAT5mqO6OBS4zkxuoEsEI68MCFVK9uGIeBBJds1a3j0I
63cPdf1x3Etf54vemsU62E9l783abAgN+bATXFQJ2xkToiS/3jJc3uzeDD1YzTk+mWyGD+Tkaobs
1phR6GEkuQL4AHASN6AOsh7zQjELv/XG7zplV+urCqHP2IBYcmkWycOvOXJ6cOWmz1fUH3PH2dUU
MmUBOfnIK+4Yo442oGIkNYtg3TFW848VEt4Esa/+sW6R68GViQxbg+Thncz7h1GmX6QN+PszM/dM
cZwyHxdqsnfMz0WM4pSx2CPTwGIUH+q6caP9R+teEABNlxJZjOwfRvqPur/83f9/GBdWCTJxYi00
hiwonjHaIT+zfCYr4raDmzlrdu0sjkdw4691KzYAxs72v1hKXFJAQtvNfasaR5QUfKNYEXo/itOs
UKKtzmIwSoRbngGDuHcWWtak6avb+i6BIUHYYLZTiGYj6w1iqCRUDxRDXI1zi3WYIzvjXT4Z4M3f
3ERrIkXOeq4vV3okTk0gIek028RIPZ0CJUQPREeJ00RBCRTzNCUbSkaeyIB3RDo9nWDXEqL7S56Z
5mFYKrzs9uRXmGok7DYDJrOGoqHybkCni5lOWB7ZHDKpxTa4KngPVsRJ8ucanSeBEFAsH4RiCyee
VKp3xyFI/mOWv4sFYr6Pwb0+XpPFEl/7kWbul1VUxILQx+GeVNI/tU3gE2yCEyt1q04sd8yyfx89
DaRWoTQBKECqIpDR6RxL+SEXjlRAnOhC8JXsMerO4SIkixB1seS77nnWXcJmyTDCMjFMtASkLxw7
A0NSmBYAjxqp6hoZeAqvsCjQhdeyIVqzkgVwYLLVhidOIzIUHw0x2mpsDZdSeYZ6Y2alnsCKnpSO
p55T/ddY5faK/gGX6IoFxdI+LCuwtz9jD92yx7gttPBR1XfG0LnbvMvMePiGKYAAj7LZNrFi3UVW
TEIxeMwF1Nlf0HIPQgnp7ZaXge4PUqBO+51UkJRy9sboCeU/FpiMTbs3QiA15bAiD4ormE/1ATSJ
63XPlee1lkgMaSoY9XoOdh6r25RwPmCEjBU0neTOiC8WUS2ZGjBVu+4vm2oN8rL4I6wamiAfnB2K
5Jgyf1z5k9fEf2Pi4htiHWqh0ZfOmGorAABmnqX7uPf+c/zBId5HMZVUkPMnDfJvqlj/owqLG2Ke
NSmJWQ2x2daZvGmIcVC4TpI+3xpNyZd4kK7wuhZ3NrHJAhThTo6uWkA0yVjMADgOoTOvuJuOW20i
TEn5TMsARKwMtp5Ci18NhSJA2Xhu/aOYTYKkPPrX2b94g569wLukeBsIUE8op7F0zpte8veRk4mK
UqXr1Zo+QR3Dy0gMbqEG2NxIZgeiUWWvUa5rrjXH4UqQ9AS+4k1bh8Cs6aQyf0C2i3myypbowyVg
g4ue/EvmacStxqEsUVQF3vO74ECbwnEdpPi/Rok/Ld3T5xyuTB58Xb4xysisQwEkcRgtrPW64vAQ
ZtlkSEFyJgxiJZQBwf1R7mNy+Xy2RkU1+OMOIo8AoCUP37RWQszylcNFvSQGVCqNmLT8a7vcejyo
/KJig2zKVEieTs5oNwfFZIfX7RhgrN1YkTDCv8IZDesoTcdU9aBJZxGcc8gNh0gVouaOZY/+B7hU
ASo9P2TVRIaOlEoDMHxSH5UqjpICtANDyi/Luxbf1vyRh1X8GRme6A/7w/vdJSu02lSTiRsy87RC
c0qnm25DS0AG39tS5KGFV9tpq7BGf9GX3hXRK5NtlD/NdT4bUNqZ6jai4iqanf52cTjhzYNFU1lw
i+NPBahEDlygzm0SFJ4XAI2C5o9aD7inFOkygTh3u0F9Ozp2QIuCM3x5xj2PYtEcIVRJlIg4TobP
id738vY5yG4sDkcyaUmgJeUsXOvc9/uTcEv6woCUbsSZeM5k70Obo1wl8tgD/ChebqtrUWidtEhC
QoLGB9yeLSR1NeLeK9HX34vso4l+txvIHsKsB5wlO4J0eBVwRb8+fc9LajgNuAWKyXUp/XH2TWj9
jOrtptV0LpnXKwuD3v04d8b9kDLiKxgB+XbsYTKTjQ+PbFvnWT8hFhU9/cGmjBZSCDotor+a1H+d
y6MJna0+x5b4vs42DjvybZLFg2jpRaJruSqVm89ArvWBUE7+9sxu9pYo2F5t+dkeiqgaWU31mW6Y
kyzsIl51iGaVodRsWmrMuiEfN9U9NhlxhbrhCDki/oiKCl3uyJKmAH5bNgRSDXGfbyMX8kK5fRwD
T+87MbV8ADAOZ11rBBmUmpXLfr26WwwOM7qVAhNQhQJZgdJNKIyqAeH/FywU9KO636Il55zi57qp
NfPHX3Jgy+RBkFa++TG8DPxg7do0QjZNIDU2/QtC1QK2WirSCKxTrwxD+PLkoAkhSt6wCqWbr2ti
mDqMvL5T7jb6wulC7hkAInyqJd6wIzFvshcOHlJ30qR2gsqcaSk476izKkA0Lp+2bNC4q4DK9/PN
6h+oWOESKWp+VatuBeA/ToHg7aRqxAOgOi7zSZRM2SatL8o02h/qQVadtn379GS5LG3cFSlRDIjZ
D/bteCzJgO4nywMuVsjAfbbZ/6bSVAPXn4MCZm2+UrRpTz8lbz0G9p2OetrMFjeQ0ZsOtbpD295J
GC55H+yzZ5l3HxW/gEu0sEXeRff6Jd4hysiWvM9vHfydrduY07LPeMrfNFI/DZUkm/qAMO4RPYFx
IMSeyRFHAzDoBBZSHpjpumHW2P4b4UCnGeIPcsRPOKujsTk5xIFmIaKvjH6GORcXIPZeEYib5WT7
aEtEwD1nb+NGHd4fHX594n6CRJRkwmXysA8hjBgcY68W3js97b4YwfjmJDuH8X/AWGu1jlvRDiAV
1aoTSxLb3Yrg5dgLYq/apgxiajKF3YptPjLvVSSMvBsP1cyJp78NJekKpq4hoefTzMT+/UKb6YgU
wuJx4jfqxRorxSd9eqnMzV5RqRNlxYx4E/ES74brizA5gBpzrDhUtnP3MF3BEurRPwSnmcAFcwwg
iEaLNljffKkQcidrUZWK7bv/2Z4ugaL6VywSmUnochG8smeopQCoEr5+Y6cT419HmxHeZ/DyieOr
olzaZ05cTecBBNJS7IZI3+vQwWv8bi1xwL/NWxhGOQZJMAUJ/T/ET9kKMh3I81dz8xeqYyz+AD/q
6CQqzcQ0w/qHsNSx6JrBTV+29zqrCr7CSOmDnj1Vk9oJpT5sTjmfdeNInxnFiGD1MkyxExw9v5ua
LOjsFmmxpCM8QJVLSPhVY9hGUPSht2DYLa1Idf09EuQ7QN+spCSuGzh5/AloRXa2x5D+2i+OkdBU
MtysvyEcmh3uUMOca3QMbTt3vcS0PVHX5oX916u/2doPlmJ9uqkYpnfFbuR3vX+e3EbzaUzOf+Kf
ODdDccY9vUceqZSaNlsiFG9+b9+woRs/WMQdo0Bpl490l4VdZCMZ0rOkQK7+Xu25+3903nGxlaNR
9PzzdgQ6/GO8IunRZSIGj1U4YcfyINHlw7FN2MobaQH8shX+pgHX1qW0W2/tbjUZfyYugUs2uQom
G3mPjbCgSRDNWEzJlTYEQonqpQvlenKzXab9/GbR/f1ViHdXPnfy2aCRK8kKp7YinB6QDk+k6oyX
YpNeXVmWLP2Xfqay2VmyC+E8NJi7C+T1fRiupJzxzK4L9Ziwyk0F8VVxwxFCxz+6+FaWpNaEWtTY
oj5IfcgNNJbDv5LvjqgMTkVK5LSiHmB/NLTYQyvzwG2NrOB6XTt9HM64ljykbIWG7cfGcJfR3aMj
+gG2jggGt5FIevuQyiBoxNs0jffcxKZocC7my4wGU2VI0Mvi2qmke63uEw5RN1kIGpFlRIKHIaav
9f9fKMuC8EizaRbrDmcNnCvrYiAJrob0TSjryx6DyOJjY5YrMENjoNAjXOCKBzULvnRKJJSByvTA
a7voEAQLvrP0qSOtqYY/LoeJpcGNsN4tfIVXxhOo4tmcVWMw9aHafVNfxPbavfKOK/vntcTOJ9qN
gd2FrigiWlbh46ylSAB4/D2ATTsDvSDialYnIw+zmegnLuoHNHfV1Z5xq1/Ld2u0FnkqaW4HZxn9
Xi/9IdLR3Xko5Kk+xKC/uw2dwvRiUrdx1ZckuuVyoNmfLmzLfzPgG39VGfZAO4fDwFRGbnQST1f2
3/YBrAiZhODHbcBBnGB5bvdXb+6nseqQF4odUYXvMImuxIlgajvWWcWXf5vMZzLuGLVhcnp6ugko
QVs4gcyRpU7Hw6JarUxabM7rB6L+SOMXPh45/yDHsGiutT2W1JCMa5/J8WTBlLyCuxjVURkL8SCk
vVmZr5uPsL7EMdpdzx5xnZzUztBNrrRXSw3j5pIarQU/Os8R5WcLGHFTbVSKpUIxV1UGVyNOljGE
sXIYeJvU1p/7eNnBwOA4DXoH62OSRl9QtJbVBhxOjSOkNKVstFcehavIJsghx0tYjxPxIuw5gTBO
BciBhcslajJG9ciFpON6cy7T2d6js7ttuIZdTycMEJ11RrZd13EHSydfQsxjMZFXDNzfRePyoKpa
DvFLPysOnRkkSbgTUQZ5zNnxlaLiHEuxuECNHRO+1ITFCk4oKrSC6aSSipcQsGOh0FUUfdUV/Ou3
vI5AFGXbc6nV76rxBKo9CbgKAMD3cK0ukoF8OuIQZV4NaaPQNhUVGBIK9P1/qdzVzU+hzCPHFSGI
gViUyuu/HWCuPVJClWhxF+kR0lzhfK42eMsP3Oh3rehSGzcMTD3nfre42SMgAbtHRLhQw4nZlzf8
o1rR0ByKvlRkIOy785+a2xYQiU8+ayJ/jGcEZCBupgt945wcfmKitzBHuXl5Noe2P9CENuzbx9/0
SIo3eO80JJ4dtzqVP4lm6xqFX4zp0FVqoq25N9eSl0OvZgYEeEHla1C531ucjm2Hbx70TJImD1Ik
lGV+kXVVg8vd9bx1ogirkzgSK79Vc0k9+ZCLUNWLKN9deFs1ZFVjDEn1F1HAXRDMJhZLjmfi5NIJ
NYZLSq13Suj8p3OTR0YASVb6WUPl/JG2rOoWd58psbyNcTYk+YponXZSD26BeY7o8TPvDMqtupDS
RkBRZ8ezZi3ZhK8q0vAnYm6/vHfTOxGDb40glJTMN17SjHBpI3i7tpHnIb9bv3RR1a4YlUiEG92y
+hhUE6waoDhYanR+9r4Lx4L7pAbcdAYxAP1gYQvZ8eILsvNkwA8QYL40xBaUx9lY5Gwdn5I47OGK
Xh0s0CxYK4bO93Zv5TehFzijuU+1fSNUWu47gEZgX4gx1MEy8Tb/NuE5P6fPMPc1a2xkf4EGsjt9
Nysdj+Bm/6SSGryQkL4ablX32gWSSJ33c0Mv11F8ppwelM8F1a7bgT5vG0wlkA/EIkvBqgf3kZcH
zhtVMJZyymuo1hSch0GMUZc0ydxbJ5AEiFOno/Dp5wGxcNl1Rc1BjT1c7RAJV6az8UvJDB0+30MT
JC18VxgcEgADdFM71L9tek9m2R+TazeH3WliHesexLkr5XC9wxtxD4VpOeJQeKElQVr+6IwmsIne
CzBwVeQ2k69LNJcTrgjyyZK1RG5yWLSdfPm1MLNMNeu7GYdMQfvhhmW4E+T2QTVEwNM+qFU5zguy
9Xys6neiLTmawaIByYd/3yW447Os1td6gctR/IikW2zjN5sivULGxMqKcGDNGX7CxVJ35BSVp29L
S11vwLCgivrcslcU8qnTqksZkFAKimLEZH6iBtWTbIThVoJVXrJAMrElvvOFzNJq1XXUV9C6aPto
URLWxdxPFB5dARjuA4FcNntDM1SeYqinViDNC52rAszL4cblymOR0L55HXjBN5ixcvxZ9gjx0sN8
2kmdkXhjvmiH4WKh+1S34erIEPttTOcNCruxtV5EUDtEjhFizwaPPD81+yK48J48IG8pB0jjfR8k
Rkw2VlSc7gsrXiaK0hA2uQBoF8jHZMPqJVgtAwFNsFw3FtS1PcQKa185BZ6ITV6zMR8h4sbjDbUA
QvebWEV4ysY96NM69U71rPIsV1PN5/ML+QfMzep8RdFJ/YLXLdXmkBhEl0qJ4oBuIPOKb/ffFXTy
chd2lTjFozUk6A3ZznHANEaxfmYHd4BhJlix5t5hzJsF1G9zreE4nBYctuPUlUySsibE1eKyjFSn
UByVnFHkr6sWfZeGS8uzAtwAAY+vsG5G97f0w4cf2Qx4ILOWCuH0T6Ts2C23hAzsU0RwlzX42hZU
xfYGPgb3PkKQqHF5hxu5S5evMRNidYXZaHZcqGKZnl/VOL3vHHd2zDumYEkuIeV5Aua0ZLqhdG75
fhVZ68pSj18T65XL59KltDDBJUx/lEc/L6jaluLPequ2/PIOxEnooMxx5BmIeQ+OXRIXS91lGFfJ
3cZq7uDiWIxGwpFXKhHNPObbYGWN2WVFOG8/YjArq5fwVC5jfnB6L/qUFfOfEfKm58aUIcYwvong
vfWiNItxY3FMQ8cES4TQSBOJ6nm9NXxCP2mtyM/rW3Znsey+rduPVns6ZQyrhK/k2+5+3DLcysIG
UKLVM9/VMJEQAraUgas9Z5LMxLOobbJ660FMDCHNXbSgnElg0uoNIDGpRPR/0LBKdzVMGTvfJWtP
pU0iOnwrn9QisETBbnC7kt1tRb/3MfMtTVfKlx9hHcH7PWXLHfAIzQUkR6oBqAecB74cW9UMxD2t
GpPNENju/cy3XUraLIQ0+M5wOKFLCQDwFwTKoqQWfJKrktSMsz+q8UxJuEFpJ/mHo1qEbfgzWl2q
+mZmzfj4dO1ruKCphUqTntReTONmCbqU4bVabVIGxmWk9fAJfdQiZCAdJDjRahBXSr8u/BqZeqNF
fFQr5jDU07mKbW3jAP3JfVZKegC/GmENWYNEwRnNcI7EmhMH/fBwFIcYHRuxM+NppDQpi2S+4pDK
iHAfk7awPDJgoC60Z785ki4bd7WsMxTtjATqY/rDJpciYvCa1/OnK/mEoO6VFeYWnv5uAU7dV+Yq
022xlQDdlysnfmXD7xfPFynWzn93PMkPpwmUSD+pvmRUtB1OcCwPoRT0hKidHQ9ZZUY6PejNhTAf
gsPpLyR9r6QTlpz62xzjvPt3B+WUP+vIDT8/jArXbM4384S2f1DzLwKyQ2HAKlWU+U67xS7snz20
BABtVg/BAalKYvEnIHchcjNYQJ+i4eL4OjjH0zKCq/qYIoResAsvIEBaFvxl9A8/LIQ0Osqd+R+q
EkQfLFvSfmIFvl7ihRmy+wn7qJAeb4AJETnWzhePW7tpgZEzPmbjYTDg0FBHk+2sZDMCqEBw/Wvn
VWW1zBYhNpPlGBqXLNnnZJJb1k9AwR0aMEGM4SbjLebyoVk0Uc+6lcupQuK/AyCd4AKDVxlI+MQZ
8OB4MO1YQaHwqgzvHv7EGpNnOIO9GcLRzURPiMqW2ahWbbUIODMIgyhwGwP+rhxPbFVtipq4s79M
mHfGFxZy0qnS9e93DXaDbC5S5jUKiA4kcPTmhgYAb9N2LDrOF9dGghd06IdpzRtOGmLuf+bdOl1I
4iocKAdw+LEgfjaYp4T+jqUZnA+vIJT7uPRT9naFcaZKDeASXwDP5XZcv7vUNCYorfgUtj8pVn6R
ArD/ssBi+p362OnY3xM7e4Fb9RaSKVPXFLbJA3tCf1hkBeQTMmev/ZyrytyTEQNRcRFYEK2zQNTx
Oo2q2Zs0XhoWuVl9EVRQHju6YvyRIHCBfGAcigQHc6w38ATzxRLy5I9jkXmGF+P9d+fypywO2op8
nW+7HQzV/R68uXtOVC1Kv2TYbLcDbVS+zLRkJU5Io5YfSPcgch6qPjPW0eBQXRrO0sFV5w3Kw5P7
oZrZf94q3GmaieC/aQLdj3P69gijWRElpROWKlMfYXhWKUAojgzUCKyeVhSYCZLzlq+IU26j2dlH
HfQKlW5tUIJAErTqLVU3TfI9gVkeZ9bpGG+FEC/yLm9DxHJZtji4OgXV5VwHJHUc622o324oNebS
K1OOxQazIgxWWbuEuEsc2pb5c9U+P4FnMnKtLixZgSAzO5bIa9czVnA3RdZIvEnrkcSBELnkWiGj
1cxAYE4effduZbiSim7q2nbXZd6vbdX23DjJOHpZ3uNAaXZLxrhlWiX9luSHMIMtL/lUJQmKh3rF
nQl1iKBnD+C4yJ+4Vdw6xm+VROtWxU1T7C5Tv0p+nzbT2kgcs2+cxT9TjU0GSePm0+n1B/ZPYgI0
HqYKbetc2DTmuySirG/opto4b1+vrN3J9d+rfpkVmB+4cgncCHcZcQXnR228f+N6iHEF3+yLagE1
FRL6Yua1yg6ejY8qPKHz0gjs74F//P76ZPOsbV83/WR642G3zkaJ/AQVczADMgEhNclt9Em8K9HM
IP20TCtIhUcYEQpo9oktz5pqRhcmAlSTH4A6nzehSSRa1JV2eNfBOCnLHs7TE5+0JVqfnzz3MHl9
KUuq8wUNHAMWtK8UFgzn/MudaFgKzlyD4NtSWmjPZTeyxGyvIb82Uyb/Rsbf1mv8GysoOVHTTWxx
CVXnbUzcnxFPT7zyJCMJ2gkatGO4llM2cNPdeQkAA56AKdK4gc44cPpNtA72KppkhW4OFXabzIs7
VCos/2c1moWhuJVzHz1ZCODdauz4o5N15zgrGUqYWIfnxsEUAcBmddP1j4GoRE89SaOytvhnU1tA
F18OLB1ztKVX/EOWpN3LnkOoRH7eqC1zAarrZgI1Y854dO3JFakfV6EgfaMVBeHFV+EOrMy3DEIC
ogBCk6RLRk7ekqSepkDHYPV1E315LPT5mCOgwby1XYBsqSxa9UYdiM3RWvxdFjOxT1P0DkTieySC
JcXRVKHaNiwzQYedbL7/whvvLfNTHXQ3onjfH/lvFCQ0Cmt3bg7ZZ/FDQ6hZOSvpPdrfcGaVB02m
Mm18bGT4TdhSzgTsgknk41ybjaG5icLU0cqwizOi/+eE0k8uETGJtaLZYdM2P6Bu1VXXyKpikZtE
/ooG7m6JmLD9u0fSodOYAspGQUB1nIZs2VtR5CfZJoBtLQCd9uFvmKAKhYWKLEw23fd+F1Bbc3cv
CUEzzPo6HCbTgZGOUO0cCHE28LMmLWwM72af3jyqb6YAKiDniD5I6cZQzKNcy+R1n6dyHgP1Na3H
H2k3NrpF1epkeCWawb0OXlPuKvcjQMtHxb0bedvB1jvgDPcbSjfMx9ikvDvGpBMJ6bOQACoj5NR3
fhasWxkJ+CQzbskwDQPcgysoYXlGUnmAcfEn5LuKr1sS0IYlqjRJZUlsIhlAzGGCrcyzT0o8Jvfi
EkSYTYlTddV1N2dsEQHh9toEPbTtkbRvcO2NKcJ9JW5gSns4L9H5F9O0AQG4jS8/dxx+JiuatHZY
h6+T0wD8XMgPzeN0IDUZ+1bPhPr6/1jmEB8bKXpHAc9N8sSwqGoTYWUWyuZBbZlHQX/tBxV/3kKb
bt11dBSCOy3a65Jvlpk0l2QZdypWMSaUNcJLBfd1Gof7hWSQGcgcfImHOqYytmh8X6ggDOguZo3p
rzrcidG17m5h3Unc1CmbjppTmbohOFAXIJ2BqPGOeVHu0Le19QT6pvgvCeszFT0nCLvXX8mR9DII
1tJZp4qZFrz0I4NM4TQ6UI5WiC0gMCiNU2QZwjJVLDJkWImNLtnehY5onmkv6kv5sT+9zcgoDPLM
0k2CFwb1WoQeiyhBGeqwX8h9zFqkeLPHrZZSFYKJXlx5E3etqePpzAFqAoP4eE9d438+Rdzioiq3
6m7aySBC+MdSvcXWp3mYrMz40yntpmKKNvOYCC0JyA4Z/6bWIJJLPBh7Jmz+jyA4czNej7uUHEYG
16B8KsGm92WzR6ioCxucOMeJY+nAqwAQ7OkWePud/tHzKWpoCJViBZTBV/sCVs75gqt9u88TXAx/
XTdXqjzfw96CUZ1dImSkiu4L2aVOP9P8ZVB5cGAD5YrT9z0Y5EnxBWicCzoYI9JD8uMMeLCSQEiS
Zl7ZvT0ZNPZhpyFiTU9TrX4yE8A2TPgkPdzVOUicm/bgk3STcew8bc4MRnatfRzT1e2iNiJJtGNQ
PqLK0OmNVy/2gXpZh+RO7RZGblOzbci39j3cF5O1Cnh2YZoRZ5BuK8ZslbhJ1jxJGaRYblJV4keQ
TKJpPWbkiXfVSXiE9DIgUpvZHjlBFIxdbcJ3e/D8S3GgsZyoELZ3Y45bKlhcHYyFQv+28iyho9F0
kv+VVwKKY+TjbHg7dROQfBxf8SieTwZS+u8hSWDMV7GWHVUslpAq431JGDv4X3n4LlHjQdd7kZpX
FSOfsaVaOA9yTpWREgdnKjXK/c6wQEY+1aFG/wu+1TCQ4Jh9rLbg8XpLPXEci0IV4iKPXaZcC9Ju
ltZ4MWxtVRynXk7kORqRctRaaEFh8ZoUR0SooShiVvrRfyCpqFvxVQx2ZrN6TMjufAPqXvc02yhh
gU6EmrN3we+ivSL39ZAvtqjNzXCfsISTM2TFSzsqEdFYASQ9WYEKCAYRsdxw4t19qU4epvIRVgeO
GeA7nFdkTggBXBugO+trkuk2vyekYasxcBbymRUgF8/eZm1aINw9VbgF+nuSZof9ie9p1wGuxLtI
TPs6n4kpO6f3TX2PlSPwVPRqB3ToqxyM7h2KRbAWzLAoqnOmlXM1KoFUBvoHQ7hkAKyzGdK/SR7L
eCnzEyQsQc1psuqLf933Yfe9eF2R9YaLQJiE65/l+8fUqsaDalF2X0BMNZKeDel5ui2iudkt10FG
ajp3AIdGJWyNrP1u6+mnnhX8Fz8wAXO+pJ050PAeAj3BYu9eP7Bl+o8eb5qamxXTpKt7vCm1ctNo
fJOxr6sqZ95MNHJfEKygKGMMzQuNyQMDTjmleT1dFcmKwTglr48S25d7P+FpXsyuTr5oKfjlElCU
MGizaeJfRIaCDALo8+WUiVXoydUU+TnzHOSr9FPVtwDnSO0MZfShpss/M3dIWI/vqc3n55GE06A4
xz8foYK5/nuJ+35TjWhzYwbcbXRcEDlE03AAb7j5kcl4AjiLzuiTQFxFSnn6RQNgRwFzy/ek6FJw
jiF8xP6ulxwm5EFAcoo2Bx9Su1XVtJW3NGpeAfDMxeVNRIl8lym9Cqfa8EFkF3hPtUlo3AeMi+B9
apgzP0WGEYWmXRNGAQg6N3rOEzZ24+lRGdWfi2B7PLhwFbpcmYVqfKQpETXvfhuIc53oK7sZIaLQ
YzAR4P8RzVH5+eYjXHLybh8wuTTZDmUHI6GtzYXmI5U788xBvCW7OkgS7PXOMjy9hxpCijayv1jE
ditEEhEPWBeRP6ARzMLZ19VqrQBwGlmk5Vz8wXJveUVnqMJf5CgzvDgJ3pRBVfgflxY2Q7EvjnJ4
4A+SW+Wepp0U9WM3AwKHc6n58l5T3Snq7+pbHFOs2G4vsIQ61sGofiJrAGFKYm1vXK57hwVW1tAL
27gjjMROk4SIJooV/LFjuAGEdlspRDHnFp8oMz+kDzqURTTVXBOiCsmRdpF4IqbZZjOmrVMVyv0a
yyQiVohAO8QSpy+4yRb2gTKwj2uO8LfeOXmScp48aMsKlghs622WzGLloywAwDLDH8PVI5brKaaj
uioyg5UF3si6bV7cHE+y2kV0inE5PhRZzoBlKIfZvb7lDYnYiBHPFcJOyNGcHoYZ0Fqb5k11yQ7n
hYNXXqcdxH9vnvztVAZAepVCz0/u73+VYVMIiXdGmiNGx4d1nTauD+uJKgKoXvK4eySdEalSxh+/
e9bnT7KY1e/0GU/xj1TdzcK1io67NWJGrTrqtZ5o+/za6MtiqSdcmyPINXZ7Rz6GoLfFOsrXnXRB
S6vV+YVkagyo+reC7wmcgQdrI3LLm0rIfsdFV+u54YJOx4wPkyihtknB/eQO9VvlvC6XCT9V+2X/
xiRTqOa6PCGgaqxr8WbTJw0E5b3XXAUXs9gBhxZJawVDovZzqdbZ6+XsJ0lnEYecYEC0ijG3jlkn
5cv2h/jLO2YXLxyXigW+rItxQX9F1rCPoXqvwFctm6/SXrK6jOBytbTPzhYaYX/UdtfWUfqKoI9Y
fiMRQ9v/Psh5I+hL9TZMVBnkN1OXpZ3iJ8yRpjNmIYiDmRBs4BIK7b+wtoXSMuA2DjZhz4WgrOp4
xSzXd67sLPB87Fv0iRpBvv0ls4aLAr+msaN0GHGLTf+Qws1pd9bk8mUgf2O+ulLXPhk1OyHflmok
2pLk171sY+2HwrPlQDinfRfB+IO0m+KdGUbxLE76yLQfX6i+EwcXyR4xB8SF7F6YCMBdYX55EVuI
VWnveSIHVdCwO2eaQRotlts0yefikpL0r1VCd9+ElW+EF2hH3tMk91P32uz6ieiMpDR0lCCezQz2
FFhubkBzTbPwnlJZ45ipmUoCt0sBMhk022L6ui3m0aBqy5u36lokXqM7Jf57R4GhC9mVu0RNF1ya
EwJU2yC+OaomjPyk3yp0+4Pinqsw5hnR+0LCQAGtvVm2+O4/YjxW6wsx3czEzloODapExVKjwxdW
XfnCHZrVDFdNElmdVbeCHq0kLCaMlVhkvA9+3JkLorcnspg0q9RAZ5ukg9/b9sUNkWEPkGduqatl
0TWh173iXN4WPCLZgExKRbDQx1IeP3o6XXFpyTBrvqHVuIjVtSL33CZjzMXJhzQmT1UiRDFBIPZ0
Xvx3zswdxTuAggqVuuIsE46vz++Kaxx1G1pnguooRHScRV3lFSuj6z665UOxnIyMslQIVXXWZN9a
2e9diH+pq5ZTgJOlp1u+3J4wnqn2XwjCkN/31ICm8duOkaBu8UzmmihTpARw2fmf07vVxwLUTwKp
dD/xlFrGVoYDrtdTMizrgo/Jd2+mHS6XoiZj6OdycKewaiQAA8QXz8PYvsEzp1uU9yi4CnNhOPAV
Xep7KFD53l/waBq6Di5qYUpG1Vi3nvUo3Wd9Izh6pHIoDlXNEdL1og+mJq6uL1Yv5e//nhTGg3wN
O8lxgfl6CcmqFB3E/N/D9/59a/8T44nmk1xB70+/ACi+OBKYlA83BUJMMaGGJd4L183NMVISB5xN
tPwEXOuaii03iz7sKX8bzHEEYMMkoE1/SrAvoR0AMf5056amcYabggWWelQqXrPeupFXIy7xZAtz
52BO9qXqMe/kD9sbsYqgDrsbs/TMjzYFLMavC2WpeAdWnUdqgyAnqWTAwOWvVeStQrTKkm0ndh+V
9HE9tfdPmsi4a+Sa0miEzBLm7sppKsGP1SVZI00BMyhXlNLJvr5Cgxb5MNs2oH9oFwomx97bRY0Y
q5nLU9RdyQC/6uo76ASiLnPxTtVsWLxwX5YBq5lYcbbWh9qYwHrb+I6IUffr9FcJEgkICKGhEydO
ZATJdrGOQ6oLOH5OaYU7IE6tFqMwM38Zshih8e0885XRXSvS4Y68OjniXdhQNPVWmh/ruQn8hOsE
zeE8MNG9rrXpeyTtUM3om30i0h7Put5WY255lXhXkOEs43t9HNIWSVcmkrgi6/uiADUNojs8EDX3
2hJq+BOZLB2J1l4gW/ywLBhL1VfHI0+cwQjQrQXX/dxGclvwO+ou6Fqkqkk1eNHfak7PKeikDKqz
cZs8kRKp8VvX2569KBaP6whPlDHfvWbMnILlDvFDte9pvFlSg9s856zLxOnCzXL4PhAjy1NOLbzr
Lvlj60cuyFCY3/XTeNh3HtZ5O7lK5awFik1yxIH7RwL23b+dH/JfXZth2YuWpDHVg8h9B8fii5rz
aIw6MQzAbqBUEFcyUOwV/kKcvXxQ6bhk4cNfAKKNE1XkTSjW9BnmTNd32DqfrAJc4FTT0Jl9CFwE
fldsNVhqNhzrD6t9ps4PMw+Typ11vPLGfU5tsNUoeL+Aa9N8lBxja+qEJKMxM7vJz300s7V8kkO6
lE+JbDEWIIdd6j+VaztiSx7oOak+yljNqgaG6Qgvr6s7C+KCsXrXjdMMJ3BVp/K/ahX99f7HgKos
E3rIGd4DfotQJfv+NfvGEcKomPNUk0BngyrkbpKitsRG6NKe/DzjeU1BrKu+R65WwONjPbqJ7wCD
dhIEDBgHBlDBblOO9cZpczOIY7JqejxVgnCvObmZojMLQIDM93a6SWtx1K39v1R+OEGYR8CI9OnN
7P2mBr8aNbouubR5C25PyPm/qx1ySWZf7ZumYlC3+y/pXlEDXE1l2JCZQzTunNv6qZWRz+ciWV42
UX6m7JzDi2R5YUec46+NSKGO+u4oVzjxnNUYOtd8NvsUY+GboLt+3053GP/pDpRWDucjXfmEnSJj
1mxObCUs0hsrA1tB+/gscaFEKHD9baSupKZrjU3yRlFssDP9ETD6GhRm/wricO9STl11B6l+TGo4
M7SJC9u+LWd1bt2w38z+yd6G00ZTHrpuiauTft+eJDXCke4s4Y/OXSBfDJduj4jE8WOUD8Njzh+c
rTtH9iWF+NBLunrJOWefYG5EJEaw1w9rMZ7wJuIVJGXIuA7sYDQanN7ic9G5RWJG8Rmy2ha08PKc
AF/RNCiFf7bN7ltDqhINbMWa25QkAo9sVcMP7d4cKsC4rnCCup+SABJLNzc5cO6yRj3UEPQ6tKOi
klkiclgHEpNt07zSYJVN2Wix4sE02wf71aUEyNstxSdgBddfYQeNoKUjUK3wa/e1SGT3cC++E1oL
x3GbLEiGGHxfnOwqDdueYSOYpI2JKVo7BpzyGofC+Wr2ih7WNI6JCqvK0cNb0wa4i+a+12Blo59J
G4kXZZmlkWBl9waJkYG83vrFJFD6hSzgCJJmZRxY0PUpvwxD/eotg/UnxTpxJwFIMcSPOktK+d+X
UEkAPjHkQ+wMZb6MCMWprA5JCXiHIreug8vYAgWSJKdlv3wmAgbaHqVhgLg4JiRqdRHKjA+c6MY5
XMnnKjK01glE5LGBPC1tcSxyJjTwntJI2WQ0B7VZVvD/1P91kf7ss9ggR2NLFBzGsC58O+V9d23V
hbx2eP1eqqD1pfX3tqP1Ns8ts9r/ZxbIAsfsy3HjUEx8aIigKDu1kqs7mCFESsIzrdrPYamS9RBr
UXNXKqSaT04STgaOzyVHY3BrKFP0P3VuW0SvK2fG0Lv5gDa2znSUTXa4fYTQQfGAd0HAUG4VLyOd
7lsGVQNU38sxnQ7vdh4nBzZBalo4FiVChE3cyGl58Wy85tPfTu2CIh27EW72edMbdqWF7cYAsYhs
m7JlNESsoAytpwPHc0AqWEXewAq/DXcYAZ2EdyGwXXwUgrNQ6DRCqa4x5GcHqGwxVMKQDaD43Go2
1h8RVbC5lf6y9XwX9UxYbO8bPsTKSGlmJwLbYVgjY52CBno8Oq7sgdOcsFGTtg7dTY3ix+YCkeO5
6SWU8YpAhKI1OmTI1RRz1c2J6Cy+dr2U5vQFUtkLdyzKYaC2CgHGIQmpre9W9djZiJbrIBMqgnsI
4E/noQb2qelK+1hyK8+ieeEbSAQtPE6u9U7gJTTgdY2kiuSXeUehJmx75NnHW0YS0UKEhfGVaNE9
T7nmusKSyK2zhZ4uKNtdluyowC+y0vfL57k1vN77q6RwFsU5Jlp+IJMAlFAlUWkL2+6Cb6SyU2HL
hI04Fi43dRaRAz+dKLYvA8yqx64R8Vz6YEzd2bZfKQzkiR7HvedH26xtKvDJATPAVT33U9qn6/Q4
AUsjan+x0vR0HqXScFxitsZ5F438adne4BoTQzn5al0HfBhu5YMR/w/rzTtbdrLzJVRtu5SaRCFs
FzSeviy8MNiymhV6QVckYrILNzjfCUsb1BjI1jBAwjPtA+vq+JPwDp+biipBs8v8ayvmACqAm9Ba
1WthsTNSTxlTBmkrgjHR4yNIzUF6w9Otvnav/AlbrzTrJLfI2AeXyLLpPRfMnIx8HM2QJZl6aow6
H9QSvddnn84iLGkmVrQqm3LOtY2+wgMYISX8OxRXOOWvJkcylPPMHAJqJsLkvOxNaoxQxfGCXQlf
TG9b10V116JCDUYjex79nvxv1lyu69TKHMm6Wyi+LF4dZxMwc1sBsaVnAO4fEGgWSBVcZgV/WRNk
8Z4oKalcZpOZXl4uHiG8pX1xBT5nDz5XZmYFBTYkHQSgAk+0K4tnA0XvWWM93exSIjVTW96eP6Ea
QdstahSn7StW+RD0eudEFnUQEs86etobYxV4wVGnHwXPRUcaPmKgsJWIrf9SjbI98rrBvG5N9Pvy
apdpHQJ/t8HVwj8/AJfS/8Qx0uQndKW/H9ViRsjoG37OowP53dXP5HwCTedONKhcId+qVj9lIZYr
CaMXO+kMOndHrWpLNbZXgbyIjA1k4WITdMcRFy+wLo2dOn3pCl5uXMN5/j0ASNdi5cDobcO6iFma
O1/Z3lrEkZ4gzm9fapPID2lsdSYRrpmQDf165cW/l8PsBqAwXGfUIF5StNNBXIq7bn8FyDbzcXlM
UIJjKZwYqGOOOcEau+Z3IvOZE43wY89op1ovoVT+a4RRKiOe05BaSUpepf81XSCHm/i+aql67lmb
1ykpdbX1AuOt8o3LX0r1eVxBZo5tv9dntZ58cJr3jgHRIJF8Xw1IVVF+COiy7byL3C33ObR7fC3S
zHwiNOFL9lg2HYd4agftRtirtGE55o5a0DbZD1ph/fb/Kk517yTe1Cxdt1YlJliAGv3FPNYbrOjT
m04U9hOPswWPJ3nGUXj1XcHxILxK6qR7DNIU1KfsgO7Zzla8J09qeMgo5NDNKO8IeRborQG24aRQ
xr/c0RJDC3kfqJfgCj5Lf62+wdnQreUOE3Hf+5f7VgyDpXgpVVbHPjkF6VK2ilR8RLH5bxY2SgQs
g+Tiud4vGxEqvTgEjkID+xShGt26e+S1NsIxI7JdNIwmQpXjV25DztqfL3XfGjVZqcDxZS63O+J3
trf5KIuQRlr4CKNAojIDylplexT1Am/u/Vk+E7iBCxeH3d7r2xYrkpDZm5SkUt12JHqm/SlkOVRq
oI8jQ7G331+iqy2s3HOcRIw3DvBrKGlGpyNC/kmLqZOuZPNQe1gO+1LxbQ2G3TKpGhDevl+IWFTS
HQlJTpkAU8LO/vG1HHSNwNFZEMea3NWgz0MpaO4qjzgS8IPyth1yikafgZs2L8dLuvRGr20EIo6Z
s1Dqj8uBasZU9/q1s3YQE2k/cz7Prd6aVXEMz6L95klsCgUIzuTdhZZ+cvsvNGcITXBqWB6chXv1
6fjz8ETgcDgj5NtuqGoHxJM48E5jun0aCMi3M8OUgu2AP02hsTBC2ecXOPTEiaAETnsjncz1Q4Qg
w/spnpaLIsLLE8/8NhWXee7xbs7aakl2fejz8xhABdnKp5ilRU9OcOBPskWD6aEDubWUyL6HCy2O
k0vxV74JAKgg0P1BuIkr2hqfzekHkJWoWK2O6Lxp5XlSwozRm45Zz3DvgrS4sT6wayMIxFJtTi4W
dnxy1Q0UQezCsz0uADh1JxnOfEGyltb0iHgdsJHbfUwBTvRRAdcpOJsy8bvcq0zpzjpVmbTDqYyC
YOHE8OZr0y4al1lhXNi5AKViV1P8P9UEzg6UFeoI/wlyL94bBrNeUDrN90boyRJ50crX2ucv0rIm
5coyyC85r/AHIccx1C+fNgMGFaFUywxfgnlzS3v5IV0jq/5WMazcXXKin4GbMBnBcCtkbv2DQDn0
30ShjaFBEd9DC2DswdbRK/8GnO/XF/2S5+94sBi09xJkQrE3nLh52jRCkzbLhQSfsFUeOy94kWy8
yL3Sxof+w45bvHB2sWd5zQvNoPA6kQWMtB6feXwwz/BKDxTIQ/k57nP1PengWZV6NRtMV//FL5XX
6RqljEDd4X33YBcQHC7gfOQX7caYQWl9qR8LFRbVz4U2QrOfOEY2gXZULLJ/4TOek+nfHIyFumb3
gKR+pgnM4k2YIZGZxXtP9J4OR9xjEbCl1Cst80RJ5jFpoI91EFFmb4N1MPTaj81oW+dq4iErGQPm
wr+b/YPikaUn869PToIh3p5sgUtNbAwlDTMcDl47sehwg7RsCycAA1mJCIYP/t/Rv4Q6oPwEgsqP
x7naeL35leJHDYHuVttFkPje8rP/H+kCewwjaKtJTVr3+hw4+72WReJ/d67ZKSHSN4WzOLcH3iLh
dA8uXNNhG8lHdpZq0byLrMomtX9JeVdDV3w0voL+9gIUfkYZjlBn7GklTWHYve2vCQ3LKFeDazep
dnochA2/U85Swz8GzhrFqmxdmUkMtwAtk1nhArakUq5cl0eYwwrp13/A6vmkB9VPsmmhacSmfg5p
erKetg7Hb3QfA0CX0aXbWTfSYDSvlRvl5faXSCXQPVxY45VUQ1M8loeftszO3JDe2VUka2ul8uvw
7/F70mPxYhuIk7G3X8D+Ce/7qG/po6HBEI4CgJAztVTi9myj1qeklhzDu82AkgxzPTOzpEkwyEzz
RzDbOgi8WWvhyT/0Z4BoV/317F5m7mEIJ14XMpZTsE9hOVL8lrS60Ug2J6vmCa9vRwIYGlMsDxgO
61MLSy0WJIpLHLXZPG48JcBBYdv2W2UtihJnVAdxrfJORimklz9gDWJGeSf7fiH6qoHX1TKqbX/s
dnLG1k14Um6zBxnPqdfUY52Bkx6opH1DDZV2g0/GNw/Us/l0omZfBL1uifKv/3uMsyQVCaWAsU0R
nvZtmIiLlPzNlwuukr6qRp92t4FCaBC6vYbCcy05+JVmqbbDolVN2sUPL6ALUsLnCMN2xCPdgK+V
ztlBZI+MVWvxCBeA6PDgn2b9L8sXphySn9jcyviAUeFzef3ZmrFCRkUBxKaQZ/8kkp4IrYIPNe6F
0K7JMgaz9bclv0kL1R/TgX87G9kOPfQcFBoMmNgcnIQx5DmxQeHmGPa3CeFB8B4h+trCE8VHRb9j
sU8Hf4+FhU7whKC+06vm1aa7eL37vBxwXkw92FXjpbfT3RZEEnmRfMdbX4NK2bCOO4w3D0yVPWhU
g3VYhuBcWXKWIPGwUxbeJn3MiSMFMMjSQKgKdomBpiBIIwKd/HNusnbhdAgZLaWdLjoSx7qkt1Kf
0866K/g9lO6ITDPwHwLm/kfsi0bSapgVNcXFNsBYLAdTGb5ZT0dokwQQjOGcz95vdvEWF9vDu5RU
d0pL9WG+FvxAxQ1XbsfRf8psLth6m7l33UKpvr2rw8AqdG+z0ub0Plsyqa9cSYz2EPkkug1ndBNe
C2go26r/Q2EeRzrx2rfwgEc5PPu/w0BqJYC+JxypXqW26i+dqICcZOMjyFFp1D0ha1DTN4UHdx8E
niqLNaZ31paHchQ2HlpZrhxV27cA6V1F8QUGiKPBHKxZjx9z2fkU1KdbMap4ROyfytwHLRj2G+37
FLxyzF5DNSj/4fVrbmHK33tlQun78vfqBAMoym9vrVa4cD82hP9E5y4TSuy0mf3ZjO+xbdGoGwo8
vB4yrnS8XqqZxtsf5EXlc8m0nWTPfaxRAmLHffwPP2A5fale1dSP6B7OppF2f1Y40hnxGlL4CM6H
a7iDT4ifMnl2Xl+1ktx/TMpNODHx3s4UdyQ014FVb7QrudpdNmfb+8GrItZjlf7a+d1SjzXGwRE8
jlpbvRDQzJokhYRBMyrS1Cov9bqNePYWYXO3TtZItnR5YfHalEw66hkvYOa2TCtbnKynvwAmTrwi
DBYml8p+bbysy+vDAeShYhfusszA6/67TRC089SPFXU2OERKJGv+BFVbRV+/CVvQbmCy84fN2EH1
h/Vc0TnefuRCuZ5kzr6mp02g4yH4XgucD3lh+pkA59Z2Gs662VawPVb2ueT9cYyIrJnBBA29ipHn
RNLsZhrntFdaY/nKjNY6ttgA9MTYLl0Ez3Kn+Vn/3oT7BqkhZcZ86Pw2P3UhwL1SlNUXlG67FXbi
Iq92kxRKE6dC7/HFkgH1ehLD6akFP6fatLEpe95KMltu42CGiGw7ulr4aqbYqw2S3rSRTu8lktHN
XP5ZRdOYOAHWobrd5BACDDIgsHVxCK6jDh6t5digxm4ZigUAWunPOoZmGLswk/LytTQpUbL0ZgIn
vKDHQnooYrBpPFMjMDZ/WnCLAbGcS55e/ITJgOzfSUcv6uTB2F1VQyl9tj+EaDNUnzXyAUHHChFm
OOtV1rPI07lCQJ4j3JqGBLeZbQSKWrr0/rvoLyFkXlXrBXu0VK1kn0piWttxoqU3ZUlVZlz34qd4
x2pnicUBdDIqUlgJaeIXBmBxcucrAKuOSa44JGELkHK6cxyVb6Dx9OpcJJFxL/EJVPygeNpPd1KE
tbWtvQ2Kzxk7ZGLoZoasMZCmTaKVSR6APCxlQLIa4z6YrSIk2xGRjpe0vhhli2y0FKTXch0lPnm2
qovzFEOlf4lfzIJhwKtnWJ8ejgboKVnQpQN7K10mJ31Asurf+C7PhzpjoSRDgd8LZr+77KfK9web
2D/69MeO8StwmIoBRh0MuvxixOBeh3B9jfBhlt197+KDXN7j+eI+yZ2mTnuWs+s0b7xk33tX9MFw
xv5vq5sPTxKD3orOb5ejX1e8eGAw6mEJ7dY7VdgRuhNEwMZGCCFCg0NvxiS2DR3myj5DeZo3Zm8u
4cOUfl0BkWA1Z0/4Qx6me9OHRl3JxWOpozamsAcy/KhLwkT9JxSjvuofl+uLOqKtbskvYrhsJx5J
C1YzI6gIxlVaf+6n9StgrOVO6G12PbhykuKg2sj0LvUbUFfk4gqZojR4mW6asgiH//SXRvxIxbuY
PuraE773tfiFssqyxzKjnt5DhWTxG8i/Emuoma6/OOAfbINtdB/GOKTByWVAeHuyyLd5fMsBaZWN
lGtaIou4pZhulshrgNQtMH1a2OQPYsxFNDr0n698CQ8DfXHYA0HGgn8FF9+xvayxVXc5aGiRqx0X
B1CqoQOp3LIvrufiJ0NW14heWxZzdEWG53h7Jx6+Ovbf/d/9ZGVm646hU7NNx+fcMJgFYp4XMQ32
y4F8FV9Do4cZBThzyDfl+Jvddl+Erkf2TdPUHMhK5yPbtKLD2FQ42hufeRZg3XsKg+9iaBih3R0Q
6X3z5QRcX8t+V97rwWxpUEMDIdfaAGOGXYWGkNX69T2vC3aSrRypxWvLUtJDSS3vICudyc5BgZ1j
2H+2MEQMEzcpkgU5CccWuj7wXeZJd7DQw6Dk0cY28sx/q8vAxh0Tc39p3rog0ZNjEiraWYBxoF33
OTW/Ccr1TWo+2k1Gs9xCW2um3pMbKX2X6zcJAlq1q1dLs7UJ6L5IV+9umL5T2Gk5Cm6SvNtXC/AY
BkQd8c8JF4b1o39A4N+CtBm30EKVXgGMpVbSTsYT+YYM127UhLFaJRkPFb573A7HrCd6nXJffSen
TF/Me2HPPogAqXBXhuuo59zTahMzxzLvQspmSgs4vSLAbxIWz8GOquOOiAU9fEaHZLE4glPZbgTp
brAxfSbNeMY9rx/kPfHRY80lXaeUbyZBOpJgATqPOrfBb6t8tyTolZFMxxkhrFdNBEfZv6pdfey8
rYKeUzIfDAvk6XXIbTXrR/95Vm6e3jY7tpHBem+vH6NNGKQur0z/LfF9YDdGDu8vf86IG2fZvhVx
cNw0YRHHPqBUJC5vRYMSAqcpLzT6elD6OdmvdwXPkLQDclr1bISfKw/n34c7vEGAWjibXYit/098
37hLfG2iK1YLeEklgTKbZHornTiGOLlI5OSBYB6yvSpIfMrAP9kyI0Br4GHQsgRUEeINDivH+vNB
h55A81kYPYT71TX2/6GEUvxSZn1bgI+lIq5hnj95VxWZyoG7pGdQh6eNeWZhHDHPM/kxTTH7JRRv
MitJlHnOiS/4sMUkbvOoKNeHFhDFxx1+SnehumNMiiBb6zKTvHdLCZegbO86ah2jH786pdg7HVuV
nVtfw3Kx4daJeUQFegwKUXlQKDYX1EF37/SB9fn6KFRIUrhaQvSnPQaEqOP3KeagjRt2SkjTu9yN
HulHu7j39eREWmWX4iQiU6pfL8Y9+H+qBMA2cuczMZmu7rgVKvPKAtuzrh6WVmdNBlqm/6QFTliK
E6+EaAEbdcCcdhi6ld3w2vh0VUBCgUVwIInEplTnmshDieJGSFxLcXBNlOfakJYhoP9qSV2geJLX
kZmnhXlFld2+HEdz3Tv95hI1XowYFBE+oVnoxs+Kayoobq5xWk5CUY9AJIS2FqUWc81Q1r2TDGJp
o+kMeLm1tn2QvDRE3iGRClUNsY5taJns58TxvIJgF4VfBvU1Gkfxg5yPVZ4jtFUeELjJMAUsKU7/
SLszr9zxyIVZ2MbLYaoO69DLRNpkDVEslxiTOTTQr+Z90cbj0a/LyIiXD6D5ccUwXuCJBlweM8ES
dTp31O2MLSu2qQeEJddCbi+o91hCKxsZdgoo5ic0MZeZdSnziUumDkUbUseqhek2hDJ28xPf/xNi
rXgIu5SvSFHl04wr8b7Riean8X80s6rhYiAf5hjK0y0ghHKLkY8LeEoYDPFzU+R2w8/ICPJy60xh
aAWX2ysQZQr6OJ0v7VEKsZDaeAR7BnpHPqHr8v65cSiRFF9jzlMEjHNgaOPZ0EgK0OJ/B2SqjQm1
sISCuCa0llXV2CTxtk2nLWC/YCP8iTF+4WSsL2+pUIWaoBEu1rEYaYty3yzi8Nbi8kZu9jZwnpAp
ttGM//L3wsZgLJ7deCP5Mc6fSAnwz2whNSzI2HVlkyXsWnOK11jQPIMTTmGxQKNzs0iCcbdBjbwJ
xvacQC3Wx/B9HVKxVAy/q9xGARfGSnoUr/qdVR2GzvOCiKhKsC02CglhY5lRY51+QxFOwAUDL1Ed
yMXFZgmRA3E9Wa4unwF5lOc6mjABAFJc9CPxizUG1q9HMLpn3xwlFt3Msb5HnNGaBJKUhwQkr3Ir
sCszZfv3NeUEkxgYO/+qDUAQ6cwnfBrUtWc8J8vrdbNeKEioqRAwe8YNIpu1eB8eerJLxh6v/XXW
5j/8coDS8AeKi8/1AEQ1lw3nHwIs87WWtFIgg21pTzhzS12FaEEqZw8KpLe9+T0cXwTg0e5bclgK
gWI6h0StbWleka8piQiLepm2v/ghe6HXoza3TCHvbrAeWezxkYzhv8p9KyYmvCMANhYrf6iQuKGx
ZC4+8b4Dru6qQ3fvMgJv35Cv2ttUuAF7TgpzT1oeosPVI22EF4tRCSIfGbXczpGv8/k+MiHAxj6K
g8ftbfmY0GCXl/bkqOKRpTj4oE+mxU7/BOwn5QNtOEBTwCSHIU2hRB6sdDEPTsnN3v1BKswN9kNd
UpSZnvc5q/FT0xcDAIC7WSeDzBICimD+fhkw8B6ntw+9VxPLBBFyZrV7lcZoMN6bFffDhXeGan1e
yEL+sgObVrTg/cvxxgd77TAnYB9ralNP1hBfLrkzFiVUeypof6SDYnDGRIXgzrnyrT12V3J0DnCY
oJpP6FgCLtfnlRWSuzl+DMrhF80ZYOvMZWifh6TpwwKYS/A6nosRjVO+cGYCFqFY7rrTt69coPwJ
qs6AaGjSlK2d+s7I9EKx/rgN3SRLrjRA0xMZIl9QSOIMWDtOP35MelIOJTgtwXjQFdBRcSeH8QIN
vVAqGkYwsyb+miLT/hnCGlgfT8qSRbtLl8SnzK4DNvRYOEmKCubeJhDZqhb5T6LIbd/QMBebkw9F
l7lIJBgpumo/4vTh3AmQawi4VOLiX9twH8TtSr4bpF4uBzbTJppnfDLPrnLl2YqE/+NfyUPsN0lg
3K0RpEUdEuzoAheEHwhA372wnpWZGQnxlF8yzSj/RBPxFn9MzQkExWS6h7VoFfAFnJ3Gphoo+DKg
SjAy3J5B4ZZT94uG21qrcM/CwAF/KqzlceacTkHleRj4o5/WxBKXFQMBKu3DiLkwuKmR58c/yHSM
nxkz7Nu3FvkRIAXhLXpphVDt3qVnsoRCcLFssrOnYnFzigjGZSUoLG6lJPUW8oSatmhlHwNQLmVO
UQvhHGAyVyXD9Z/EG1ZGf21JJFvhId2JEtQbI1jxt/NCgzBiC8W/ne1rNFTnL/m6Myf3aGF6HlfH
LU2cSG1RCAhkc2L2liO+K8yhZZlfdv4lPXYCqf8GKm5GpCuC3g1RCDUiHrkJjU1jPGL7keVl1wi8
gFwVPIKoGKFfLdJFru+fXB3lM+3+vTAZ0kcKyxEAnNSD91chL/3FGORqv7/sBu9BZ3wxqyvdVQ/g
pEaCTWQYMqCGIvOBDsxHiDJs67PrBqYZXYMeNUVmSqmONI2X9gIQ/TgUb4V+GsW8QapM5zRxHyL+
qKw8Ki6teFRo4AOpSi5EeD3U0fhOv9pRdhHMllnra5Ryyh+V6gn/zVtvRHlTKUTlD/J95uBP4BNP
8P4IJ6idc+7SMvmkNFie51nrsx8g6ZdweC8ZAhuTSo32UQ9DG03vZl/RgMAS2KCyat4qI+s0mvFx
EHSyw6B+kgYyasMNb5cMdLScz+t4jBr7tg26b0P2Ysn9vUh1+bkuR//KTzM6d4nqA4+J/rr72tYV
vqQkmV1QCf5WvSOusyLDz++VFtrOngrXSj/6EvpzaGftNIPvqMD0cqmzkK4cqZiIMRgBgQRE1VCB
wZPOo5rx66hZD8YQ8qw8IKEoXNaqExW9CIkHDI+AkeTGsAVS/S+jvQgd3dGWdceOg+bpRAHqZfdy
L6+DwzZQWCCkf5G+SRtWSDHZOKmArA2vFgWlEqfJ/SRSvxe1Y3a4PXOFQHknTeooU0GSEf1xosrN
p7WnbEPAeHnV4B8SOBO6kOoPg5ebhrDJR+DqZLa99c8s3SfjYDdZ0BzbSmuxt7xRPp/irEg7W8Vf
C7GSKATd0fYIevpmQectBefWZmdzgcC3qp1LnkL4+PkmgoVXzNDQoZohRH8dVNaeEyKRfHjgGB4H
+sVq+yXncw4gSFi/VDuD1e+ywFL2RG3PeZGacJ5X4Y40CthS+eVbUW6kLfouI8V5lRbwDuiajynx
2okDs8I/MDuLzDJp89sUNofqpytYH6SqO7up0GBsayXDXCtKQUWbGz7ucPIfhRFKvaWlhDw5N+ng
LO+adcpy7EGi6LLlCFqCPopeGuCwfkXv3779nmC6RtBmohrSk/LV6j57T+F3JhJ07LnYnz5dvzUK
bJMhsr4H8okAxiJUfEG23UWZtzCVGtbFqWav2tRq8cSuojpFUhDAE77LSXmZ6g0LsMsRi/BldeaJ
g/EasXq4/k7wcuM1HFdzPh5dDo7WkC97EAkfTzvKrxycRiaTRjoMoJ/Y5wfIDSA1678sZPIOscox
mh8D4LMilF60jnDT4eKoQv5BA7KzHU144RarQ8wqZ3ysSKsLMx75g8nQaIGUVmgDR6KE2TDRSXqg
b0ehVYHFgA77vwdOa/2hs2KvDB0sDN9UGKoz7a6PJAOrmX/WTVAcH9QJqKLh0t2aVqeAQCO4aADc
PghqEoHqLRBGN9OLmH3cBYgsF2/ClhtGGLQgOHpKmsN78+92Pw50HJAdt6OdnveMf90mh71k7lsg
b1lEfshTQ8LQKxKuMOITglMkLkVZzOwDdzD6i8dKQFFmONHx/6g19seK3V9fdZNNPLqECYCLnLl8
0tKCLbP56kefsrtc0gVLliu0/kuO32oSJftfihyUuSS3KjynTmvtWFJ1ow2VCp6eHaojD0gq5Ikb
kEHujqXx1UmMPbfRwCPQ6XAli6F48XHQpn6PIg3hXjOF6wxfWO9buo5aBz/jdVN83VxesZ0iD2Kv
d5Hfdq+30+MUqRbDI7L4VKz/yOWosKYpJMkQk36OSe6J9veFiQJJqtJl5dMjK36qt3oTfa6PyWMg
cAbO5uVZR/MOP8bAq5+Dd0epDmUROx0d1OV01hkhqwH4oHsDDXOuDlLcCPCftqdT6Ahr9PMSF1rg
p4X9kBd6ExGa9VjMhTUK8vtpQEwxYd2t3maaqTYA7vNyoWJ+UpQ+futdCUoUlcIXz1MMzZaoMEYT
wU8BrhjgQfwQ3btG7dvORq4UQvkJCEn8NV8fV4oXWyf6WwYqe9NuYNOVzYIPXYVekW0fg5Qa/H1/
QwitKC948smfr5rBOPnZrPepZ/WLKp8NziW8LbWyYFogbviOafwe3c8gYuwWBl4zYUZ3VrlmcYh5
/pgAhRTSyn3JOLOOuGUkpQ61of8BQ8zgJOtTtxxfkjHKiLwvN0yKxP1SMlWGaRDuRJJl0Mwuz1yV
7vqEguXoos+zYswyqS8Mlgk/jOJUvYCSw/S7BJJN8RZBqAWUe/sTSwr9HG67DcjdVwU0G73QbhFr
WPFVIrvWpkCZ+i4o8b/+xNcsTqQgyWilbvOEbZ3selXLfk4bal+DKdW9RxT3mjCUyU3b1bLbmhNs
ZuiVAPZ7Xh6LCX4o8dqmR9680taZ1GQXpEhy2yj9/JxJZFiylh3d6fEMuEl4xbbRQpdcQz9xnPm1
Fa7VjWml886DH5c8N+3uOvdIjLSvkr4aohUs7qWpJ2fwu9DtbBGXWGkyUq0Omq1g8skFuCk/3Kxz
tnIP2tKynOPu5gk438NSSipzzzC3jjCmmn8bjOlbUo1hrOcAjWee/ISNtEwgt/ZmQk3GQl0EqWPx
uzPbaUOMf5y3iNjCwz9uJU55X9n2ToqXWS1BCPVGeDo+GRpRjsJ8Fa+APdZkjMKgAJlvlMYmxOju
NHc5fs0jNPYQ+MnuQ0scLh7xsbeW/wIgaQ8OTKd004mu72rYs8YGJH+vYrnG3q0baG5WlBtWtsS+
dJj5KNQDMolt0FYRk4slh3bEEI4MQplIOgk9pLg3vOpvvE3pll/eWzODgOWU79bolvt24yEa0+d0
MJO4MsWYMmss3mUPYbGzi6dWoaa/M1q9sFX68V33z+LWrTeuvEqiN9nMmEMAMFTJgHQDSE7FK7SS
+HrddbFLIR54/bGrJrN5158dBxFk9knVSvo7qLOimxpHVKMYm2olkzw+QOIbux+JSwTQ3djOR0af
ug3+xiQPRyXuIXhjo/iKYqtFCAWlYcs+fNd/U7HRTPRqWiPYhFjCWAOq5Gp61rCaHms1cv+8s1Lh
dX/pt7+DdYdqf1ycThVDV9MwoX0fE7LF2ZWVA2Y4BcEhsVtrN/PkzGhMRfDBW28pC+18lt5wTv2E
19Trqi1HeTTlg6acw7lNiANUgGKR5g16llnrrn5hqm23RP2IdFzmTWkP6aDsJEaDTZjymB4maSCx
kAh09OHKuNljMViBHdiCObxwbS82+erBAvhy0EQDxOLdIYzmy4MBNMEFCOnAYSB5m622HbjV4RXE
VMhazY94zE2FTS9eMvyj3qwWBgt6g2lDGVlXfmRzsNFcM0iACq3UsE+8t2ezD6cJiYcbC65Wlu9r
EZJllM+69WgMRm5GBCZ+4sC4x2ZQVkogC+ghAJGb+88t3LkyYaGFPh4+iDXXJgWoAxu1XLLOasiI
UqE72KnkJWm0HTjbgw9m4IygnEiCytq5NbVHfL/eYryVOjuRx5jRCXK6qERaRXxm5u24G62PQBEO
TAMsyCdOaekQRj2Gbx+ERLaUYWXJnMAIyGd/aO0O1TH0edqM162Vl22Ro6DkhnmWl5ZnORZOvJAy
06HpBK8YQhSAkJFp7Re4Aduld8VSOv1wW/ER/48nQik9kwTSS0Vrh65FVW6/IQvfIVNOn779soiU
9U7ng9dn6GURfl+K5rINX2kYvUYD6nqA8ox9aSoyDsDPgcJCKqe6vswSTZhbh2r3kli08+9mHwWK
0bWIk5lhasH1Yg50hxcMEZP49gJkJs0PSxOTeGw74o68aKTnDaGT8wVQGhJ3us31qrNKqRDz5qlX
ULyNl/sroffYZWXNZnmEPxkeuUju/nPOchzSgNaIFaT754n/4q8JYV4MIWdVsHiCEC0dKqmRmhMp
Kc05DkuthbKLh/eDhX6FlS7ZGzm7iVi6k4qlLTjb1/Fy0puEMiMtH3qrhDwur8QEkPe2E97JbWpe
aj+nCkmBZTCcmnEvW5MTKUCGZgi2TyqsV0RaCsaxGu+Z9P7XzXvwOaIZwn1X6xMLtuxuEejvsWLA
aSVZw4F0J38P6ZGZnnsogEpkbqJdw9ZKX7KzlVsZALr16q3iNw6z1t5J/LT7uIaFgheFOmad6PIO
CHNS47/uMXyN9zl73rGj40ka8ubzqPpik/NrCHN+i8aCIhiQMis5RPH1sULbkGOIK+aAnVLhaVBg
Sl3KgwtHUVDeCL+bUw8UZhdIE43leS14Wz90lB5QvCNrvKesE6hvucgcyU5vfammgx2BwifcHBZ1
ddG5n6U3eOSk/C9IE15EftHFftzMPn+qKIlhsQwOKiJ7Ou2fxFthkltlsj3L09HIoTybuNIk6D2B
+BWRUqBkBEy5nbB9We67fd55DvLfUiOuSVHEZa9iKCZmLEqg+RAIrRZTsqio+hJb09m9ndKcfsUj
LnXO79RmiTXBl1Z2Y/ilr9VFspzSq8qDMonJqcG3+5/1xcNkBabHnBEbKDza7om6xLGFO0PwUlDI
YeyeeTdsf9kfbOBFuD1zlAVyr1tc/O6GNBW1ZZJ2B+ZWrw01ueVoG+ZV9RlnME4DDwnb108K+0gO
VtDrSw1VxQcglehRsfdDMDTa9G2W/J+GFB2YsYeMZc8u+XwzAO/8fvyEY4vViB6FvW5pL9g0+Alv
Hkk9oi6iEK4ckP8n7v60UjFaMwQF14ILVlH4nYyUbBDt2bjAHRy+0yz2YsGseuCReh8//M16yVyC
LptiFP+jKQAl9EMAoENDjY2sngwX1NEhv8sdn7GJzy1wuJag8V4vlNBoclnqO3D/M61QAyBcBoV0
RYFjXa/tEYXnjFb/1ac+ZFVUwu2wiBt6nqzw6tVnrXe4UyasbNDsmAD7j80l9ibtRzA34lsn5+bX
CyuTTXdKAOfvriwUgFYDeAfDBH8CRvdAwcx2s8zYgoHkaKkQHdz4mC+xrf/zXG3Nk9ETdkJ60s9j
KNYCcge4zanJP4v+kbGRMzfsGmDGfNsaniZwRc9PQfuRiJklwXyk2Ul6HFgikhxiRrWUveZqV2jW
K2QftqKJdixTPVPRA7s/BL0xVFEKPjhNRivFt3xMfyPHeCa4cDz8DDibfBEyP642ZjFnyTYTDRbU
4zqdCvP8lX40C/Z5LhDT0qY/lNUc150jTDdBnZmbc64b8/yYLzmTFBq+fR5qwT66pyIqUz04n+9R
r9dkQkX4z9d1ezWpq0nbox29J2BNQcmg5sOXJ83BBIyO9u8tFgXhA0+wrH8yAT46au6qdyADfnxS
mbZL+z1klVozBKMMRLX4oKIJtPLcj00+Y+tB1mag7LnN2eox5hAUDBvQmEgi93D2WRD3tirKcZ13
l2OP2bQ2hESFr0ji1XwdkquZsZR0PxQ3o67zZeL6JC4CCoTEyPKXAYx2AUOlh0rdVqiSmKhVX9Zv
D1ngjLOCu4ZKgEOHvXQ6OsFiy3XjaR2tO4bsFO2/4WkhMXiASQl8XiQtjbCd07/ukdYbGAUrv4Cg
o55sCd7XCz3vyr7hK/q9qgzMErnyGqkkxqdMEyC2ILv0Vin5zG7UiVNqChNL6ehKBRtrQBZ1zgPA
dmy+9KBja3XKtuY1QaT+LpwMA6JL6/lVr+9qGB1gMZ1JNSnnKo18CpEbgYUuYDG2o++G66PS6qB1
gIYvx7nQi8EfHxGgJhIPnjSAhNkg66MaCEaae9aak12hq4R6ZzkDvc66aY++wh0shwL17cWsolYO
LFr4QAqm4WuZtmrA2hdhkOoF8zBxLvpCrLx/2QTwTo0jb4FkKxsNRVSSPOPT0nWIQl8D6qTWbYDJ
uOkhyo+8dHi3N3S8kLEKzLODmtvVtgUX81AWAzJ4ckqgqQJ8MifoY11YMO51pY55Qu7PW5016UUB
HFfwt9vgslMHVYxgKm3ALb5bkjMIabcBSE6SIw0H0ndh39ReGJKwqC7SwDH6pFokXMw0IC/BxZJb
l9kBGsDDVaOKpbYLdDass6n2Rl+H0T7NRsv0FXc5sCL3+lJa7qpjiIp9R00Ac60BAnK11nY7EIHk
cqYO8mEAH3jATltIgizviJSOXSMGnxFvITo5MClSnin6NYWWe2MnSLQvGDs3uQfOdvurPMNt08Hz
iL2uvka8qCgCFkOwleYiEZVBTJZi1tngdz7aBfNIPHysb4xD07TR6q1qFzS2UHZ96tUK/HCF4LUK
xhTadWjCTvWYuhmTNTpDYK5j4i7pWhB7pzHLdSCsT7aPf5fNoQB2gpztAKZHRZvHInYNi2+M/gbm
fYhKpmMzrwxk4iqrrBelyNzhl+aw+fYYngqQGuFNOCoorz7NFKFyw6o/F7gHKGJzY476UtartnqL
DHrR5ecXx2Bp7UyRrkG0rDd0KJdLfC9QHw/tC+fs241HXffHQhXT4xUKIGIOUqe0+8sYr0UlG9lF
q3nJpgGEdz/DNML7goD0T7LblheJb5dzsBirOy4aD7QlLh4h9zCRWQZta/MZA1x1bptjIOWcbc8A
+SPJBN6rk8sX9ur7EYTFcQfsdkf8+8q4Kg3jwa59QHh3/XPgvdDelXoSK27OQZKTmLqrVhhZJRBs
L/JFwEo9qkB2Z/NcDbFDFa5ZMVxqA8m4L3ofTq6wCzth+odI/0pmyz98LA5seZ1bSC8XTWexnVS4
O2985RWOUF4X41qnduUPil5xK311IxetgLRjJmimBMXAAGTg6NZxobsRqwMjXx/CEQ2YCE4n2ABO
/8qrg/eT4sjKPsLELCQGFkmza+Pv6UDrZB+R1ZpcEgyIjiWaJsyLwvHQRNwBFOW6FPrdXw6D/tQA
JEXE+vc/hYc/SPiLobuK4Fgla75sorhTmlfGWFoyNHYSP6f2egIZillMagsEo0OHdlwOZY2ZnHc0
USsZ3m+CNhJf3buRhP7bdPQrQ3GMJd1MO9Nf/bJ1NlBYYZNnemFObIVIjvzuQeLBOGsaWsF0GW8+
sZm5R7St+gXFT+J8My9ihejGXC7QAfhPAowvJZESHu0hUqA9U2cKfye2nrlQguS9PZeMl9qbCx4E
cda86EeFCVi4XXDxGiS8vQOxjROcupfdyfUFtKHiVTDvFlLYXEPOhb15UEuzxV8WEMF+xTcBlhKi
nzaNAuNot81pLbhxb2yF81u6T/rohVWOVy8vySAXXQKBHyuWBgD0FVyE8C2ULRbQ/mAViOUvXC7a
kjQAdoZv/3Aps9a6ym1/AY1RiATU+0t6SXYsgzGK1Ey/3nFt3cW9ZFw0JRXkZrY7NL472gvat+dV
pLn1hy5ovrSZFY5B/JErmvXvHUFEPe8zN8z+dyLs6yuikULEW6zcnwVjag0ovniF3oyIuFULbvhh
HVfr8nF4leyFCdR120XNw5WUDtdTGq3u0lPz/qLQ9arie4SJPUViFDfeuzHdNMsnOQzrqNF8VKem
FWnDO6hhuOmtM3eyXsmjTmg26fbimiSdDSdZnDMBiEe3nyw5KSBFXBVqEIyxu4ZhnexirZpD79Fm
JY6zfdeIYhSuFR1d6iFcD74NsS6R82IDxT4Bg1cVpCwUOZu0omr7YjWIMjUamyqmI/sGjKB7+rYu
3pR3VFyiC/6573yk+xbqfC9IoAv3F+gF7RhfVbtrDaQo1q/tS74RFe2UtNy+4U1KOaqWcaecx0dL
R0cu7DXr9ywFjaUqau2+OwrcHc8bJJisdh5b2uIXP/1Up2THlXG86c5inc+ungb37MgMjq5mqlnS
Sr2dW6+ec78YcCxVHrGmmdR5bCTSF6P8KT+zecRQkPklreYsEkSkf07pc29pTsm7OnVsu/Rody4A
PG72HBtRsxQgcq3gxZE/NkwKf+SRid7lX1Dj7rwOmYXqw2sd6PM/5R1w3pJw3rIDtmUt9pz69I7u
lKCCArjdQWQjxyXGUDIwujlQ4DHT4y5HipCm8FioPzOY/z6BtDcg/NtQG5cZYiqQaP0xzWQcj4gK
+rJbJLKa45NkyU8+lsI+lTKQKDyMD7245hVnBjSQHqmEpJ2q8HltsAz1Vd9aKBL4+9WF0oPxa0K9
pD+49H5QFH2/B7dznDLnzJmIpg1ihnkmjFZFSUJYROkfRgNZAUgUdN2K7DKqYS/b6HbbT5JsmLeq
SQlDqSDG4RfMrA0pt0vKvs93TyQUBskHb/tWvhciDTdfWYq74pyyfS8FPozXDXzOMBO67/0BOnab
gxh3M+PP+vCtUpDJZpdrMkeO2WvVF7SehB0eOJaosfWbP3s9yOfbSrE7hVvkQ38xKu3Gd3VQ+EY4
m2YBiU3L4awVINGnrmxzDqT9C1fz3Fp/mdn83i7q9eGyXOMUGH3PilRDn1TfOzM99Fi/SL0V8rUs
x6gSFlw+XnXMzS3/XAJs86ffwbJhMKF5vFUHcGjT3bJwPb5nwoK4AYxflr+6+xtMuzhyttc6nRnV
bGGvYDQiFOhczqElGjWheyYq4znKc9s9FBGZewsf3vTJTXlFSUTOqaog3iKkCV0KVhpjQioXCrXr
HjZWMzkkRni+qVlPWeJyYsP1wn+Pu2gzwAsN4+1NfuS21+LXHFViU9gCal8d8g/XH7ChM1I/5lef
qFrt5DM9nFgozl1/Y1as4bhLF2aEmD8IWifQsX1WtzTcUy2iwZDfzRk11ArvPz+b0/S2DS/3RywY
XN/HyBZsRN7242MmhoCzohMm5yz+7cABxZB3cGJhETAwvxQRKG95jVt7BqZ7x+4Gu8dZcZxxtigY
vpvY2mVPkLutmWL7/yd5ALV5FqGA8gqrUhGCtUcrSCW354+HeAusSdXJ0QgdSmbmPMJMCly2Do1k
dMEUa4eAsEbKgPSdgrwZFRZpoJH2J1SpmS6Ox8ied6pJ8oxUHvtIofOz+GzrQ0QgKvaWA9cJeH4J
6O+p7gWm275NFuiVRCT3/O9QMsvpVGeKjcbrKbehHs9nFbuBL859I2pbNxOOpGBeXjvMKnl+hS/+
HvnMII5GouGXzt4CsJsrynIzqvLB6ekoQ11uneO0bAielpix0VH4uWRi+a2ZYHkCRsExvyynv4pa
jWIxJRSyV2uVAXPIVCzNz169nidseH5yfnTXlWoHiTzcPyvkMpKMG39rUM6bzo0OpZjYVjzNmTLq
C6649RQSB+7h7eu5gmAPYwCCJoq69qQgX+CixtFd5hUaP9BC9b/FvmxaYaa0qq9jpccj5jc7pVpQ
wEpKh5LvbZof2/EjtXTwoxCC8hOmTkmC4O0YxuhplxJslXHVTnT7aNpcOXxTjbmY3pmKWnvOIp85
u9Xnd9785asTilIIENgNqyz51VxCWnXb4UfPErbeKDmeJi9C0l8YPDUBLr07WqRUHmRjhhlGisAR
3wJCWFm/GE+1GyH9NA5No9helQbGe0h0lwnSw0qv/OK2dkXOTF0dTcAc9Ijl9uZvBXDnJuKuMBTW
HyuOy9343f1Rm47NRcF6929DQsCsAYL172mYm7t/L2+dsOggfrKXbr08X1Ajwl3DzGv8oEEtUKPO
YDuZCJ4/WMjXNieh+NBXTdR+x7/G2u8e8qgG8gTzTujQPDmi+sEKObkFTjSvRIPUYb7W/YGPb9NK
qcgObzGD9KAPN9PyE9+ih4zrn0E3VZlXZOf8wewe2lZiVMPFVTt1xf8AavmwCdq6cWZw6U0fkTu2
WoESOZwjge6Wgt7hafSCFFYiYFuanFmvrJKhLcBxcmgw/PHop2/mkv5G5KCCeT/ZZ2LyyYUxtLnj
zmOSG+kB95uZIRhEckecqs0xJt+Nm7fqjEGWg7G0wNXh8y2M7QipVKw7ZjXPO1JisNQi7+W0bE3p
NLfuz1YA3ldi3dIXo6Cocl1oLlLHX55cuRnNU6HIwbdxNqIlgvrXgyL69cCeA0yo/h3kvM3SKV2X
G5NZJ1ezvI8rAWF8KezpHZFLHUsvvnxBg3I+8ppil+R7bpWesOWHXUw3XWNew8REK9g8WYdLcUeG
TEWOCM4YpeDm8+l5CbdcbUH8WjojmYT9WH7+BItmgKsPWfBnRCTItungXxQp04/cjqphm+dZGg3d
SNJ2ajjEX14N9pKecbPEC5MzTHXZM+gj4zHrimLCxkMMJYOQdWCoWAKHDvYK0Rom/cKyYAotWEGe
cutgHxOiDH4h6ny4unAPYhIQ7UleQOJac0kwd1FUKEZoJT4F/nWgywISqvAnKLUIbPVwkGvoEn38
6a7/gFx36YtMY9jiIBxPLdxQ1au0RPDd1iCqSnbRR2JFNV7vDMtmDCGqeYX4LMygaCTU5/19Yh+2
m5/Lw2Ea2Yx2VmRka2e7e+hAJpx+n0lxMtctVNTYjAWeqobJi/hv+dguGvoZT5Zv+AXZAa7Ad3WG
UUZgvzi+H4zID+ygUwkmr53Pb6qr7mjeVhogaFNgh1C0YVc8Vpx82QJIdGy2EiNd4sRyelvdD6Sa
g51PlIU7HHNi23K38rbiUgJRW2GKwEdsfHo94aSp7pRRefPFLVlzl9DbY5q3tKk5ue+kKgazwAs8
ble+2Ff/uED650iJiOv1aesYvc23vcyKCyWIqY2ZO2sz3F+TrRjWjQV/NXwpjhZy7P5iFt4Ws1rm
QQ3NWQjPMw0OXOi3js0G0N9r/4tZIidxP/H9GUy9an58RNWwUgQvkleL74bsQTliiDpR+CAotWF6
0Wv3VJNH0e3VSS0McK0r8ezz+LNbRFSFB3JDvhuswqj7VKHS2eAnknmOW1abbW5R2FhsKXyck5xZ
078Hv8Db42Yql6Raz/Z2kdaptumheQNX015wOLpGN8tQQBWgAxk9fzf5TDK6K6SyVARBjtTd+7Ql
jJFlhGp1FSHfVclRKDcRnKT7nIwteiyDSxBl4poo5ngWs2y7Mbsmujnd3D/TCwi0F6GbLMX1tWUk
wm1PhdDn1GRD88LdiYokXnH2KWxqBrqgpdjZR95oCJUUXG/s3YPxnQWQ9gMB7eUmkYSa56Yj9utD
AJXF4+nDF0+BB8xI+znk5KsuWcSB2eUS0ALni5gnD41ff3ygQMNtTITYzJ2Akw2xkAEoSX/O0qMo
EcfcVuGPk9YTlgPQabxdTHjY9aIadoEOo4kxFlOZ3V7rxSqqu99ZZDO3mCDKkMUTIDcfhGhi66Id
r+jtB5IabegOyUMxj6PxUq6rRvdPb6Yg7KCOXxK5E803w2x2eXi2lAkx1V5T6yMN4GlfKf5a6c5h
pb1vKvrqV5gDtiWuYy85TZuDOqpX9rh/jQXT4RXRkZNItCfGQocP6t6iZvzu3e+6+Anuv8wRwFZs
BdGwOXNmmvyOhllqC4poYtc5R71Ex0b5In19y29GVjl2LDK+HROuwfmzH0BDa4TQ9Kn5ch1TpoMO
5XtkHE4X9o9rJk2385XW3b+w97tWnl/tbyXtEuVwlbm0T9FL3DZKelda22asuEf/myYxm6wqCtXN
GYjnDpOn/VuqmIBVqj2ok293EtwdcQ8lSWgcLUk7nOAp+vppjv8gp8iXTawZpyl4fWkOHmPMyCI1
Yu5P78eB/BX9FnwRaCVR6/sf24g1V/V9Y14I/o2Al7W+9B+Il+wUcW3214NjBPWl0IyJZytTnA73
PdWDTJ3aEVOs4pGHZe8kL56dLCeDYiXeoYgsqzbftYxcp41i4FB4KbSq8mr1SMYrK7b3OGlcb31L
sh7WJv4J2UzY/XuFAo0hhPGWgH8IxsD04Km5J+bdD88k2odHbPqLyqU8twMCzvkjVX5pNOzJ3vpw
BRZKqj00scyWyPSAuTeZVP5cudFuGHGirgraZZ99wlwBpu7d/Zd4a6hTqKHAZWknkHUmHlZXB2B+
BwxQNqnEwva5QC0h0qmex2MWiNgwZa808b/lT4YVBnxO9K8JvD72Anbos1/KzfEtGGF8HuSabKas
e5XaMvtbjQuFsWWt5o8X4tpdmEEbvSH55/NNDCW21PHHf9IgysgkoJbCjJxwVSaQTetPcdaFtllx
hLHhb1rjrtV8X1L6vrxE1AsGyuu5VRgKNqRMDrjEHjEv2mk9VhNNDOB+PsnEBkeRGpny2S7pIN3h
57p0acZDVangdtnrqr9S8x9I5N6y0KaUVDj3HhMDtI8bITcmLX6hz7NTTYSvp75R8UOOA+OcV9+R
XFBARs/rBp8ylyNRrOY4r1pci8Xo7tVBqmzLesw8kemunmwsr3FL/vh6b2R8Zo5EagRAdB6rwfrp
yAVV2P0kQETOyW0kNA9LlFmgar4JAZzxz6CA8WLoFpd2Lf+YV0u+tGUXb/8aEwr/IB/MBpKywUff
AcUgvVmetYqURDMh7vMjDn8s57j5rwHdLgV6bsB3LYFQ3F4989nRvt4iewmJLmb6YI+7k5r2Ei8Y
2QGvKp8uPUTaJKhN6PKdo8sImTXxrx1B33FHGmy7+kdaTGTXp9+PJsW03MKGJmVATwSnGGO79Gkr
hFgJSWTg3Ta5SbO16FTbqDknarREBtHJigtvY0/kxwtnr0Xo1FK22omKvzaolx444TshayZxmTaS
zqe084Ot/tmvMeFMlMp7Cgo65NroBnayzW7vteTq41d/Oahs0p890VLHewuJ6nEJfSjAS8K28+vj
ssxECJq8Tq9wh+9EOF2c9SDkz/ohbOUZ69+9iWdKERXvAXLuWZkypw9nR90Mzn65KM5LMasYDGED
2I5uwOKgh1icDYK9bSy0aFVh659+4z6+W0BI6p05G4ML2jczrYOTVVo/451uVjXEAy1Ck5YbE/In
4i5MSyh1OV4xsN7AnZoBYPYR3Bt3zGVic1egTKtaCkU0f6NVE7O2exMqNlvLgYAQVV/w6CpWF8j0
61fO0rZPU+oH2CnSqOK6Qp3yqUOrLuDnTXlBHtm3HVzsk6iuGwhdDFpdlMFBHUhLBXOJ8+CbQGYA
6KPXtjc43evoMY8Sb25ScvE7miLAAhkApYvkydxI93tbVxB1a8K6l+k2Z3Gul+miUzFNSLLg0Gma
yaeJxuYBHRppT/lXKlnzto2D0wMOOq+YUgfb5Kj1XGG348lqigfrswqv4FTqAqa9UyPd2V4kSJVG
bxwU86K6vUUGdYO58OwAuHikEQ7UYpX/r8mAKRR+wT0T3YOMPewIJSZpIp7A7hp2ZDZPCFOOjB6W
mt6lA0oKZFZ9UKvGiTUkcgQZNHTr9wj9JSvIR6PZ2erFlg3Pu+rx+iBK/OA7N4mBcxzn64QU2Zze
Wls96rBKqSyer0+pNv1xjxSIc6yBnD1RGtHBb8lXRXgMwnxcx9NpgQWq33hdo6kYDit7dRnVlqG7
ib6Y9vHudJSapyEuwQ2xvFbxOt0OMeXHEf+ITbsM9LAruNxE+HaUhOD8IPmugwhdt37iJ8QIsHvL
eo7e2PlIuStZ8NmLo5KywWKHQ6xQJEz7FOxN4HnVxu/beC92HWq4eAXPvdUS0/4YGcWrA4BLlBVk
o12q7QUTs8w1W5TVQCmwSTxJ2TALuthOwrhahDsErM1rL7X5oqO3tMX/pLsR08xUOhi6jWzrrNA2
as4YIPxo/ezs83pYIJ/9/buTS1wZWeWvL7elqc1LzfUs33GombOrX+yiDh/V8hvTJMbGdMvp+45t
JTJgkSphZNLWy9x9jU25ZAzJbOeZ6NOzAzRGa6iHTZXcsN6MIsASw+NhW26BGsijYpU6eZlxZlI6
n3G/JAYQJThJjMOnN1eyv+qX2TUjbchGw3K7ONBQtr533l+gs44xvo8ZBm8ouhNyRy2AbxMUw2+U
TDT4NLEjk3pZtgo6pBY6Zsu9rv+oUGg9ZZhQfqATk1t9EqZz0Ks/8tkoynQEaZM9MfUbfPnO5O6+
I3H2oa7GqY3E/ycHnMuFnfK+3cQ6cbhlZn/sl5+zSf4h+1pJhVhA30nOQb+hafP+xvmBPCxzFCdh
vMKs2Trd+GWwbJ+iHi1Sk/ff8C7WxqEUmFERPzFFToWiR7U7bXgUY5ta/6sScTfrwZymwa033l/Y
wz9rY0fJ/xo9nVKpHQdU5TTokkHIV7FVxem7GW9TPNXVNPbL7MVUzX4mjQXUwSaqlVEnk6WI1bjf
F+BFTNdRa7WAqPRJyhYHEplo1VWcNg3VdUehRcriXbHqkvRBVv9eNa8oid1pfZiRVK/lLCmpBnSq
JYjq+GsSagqtzDiuzbWpLTPecM3rijjCv2eJON4Ts/63lyeWKA1QqUNuwcyCk5Im3RQ2KyvTQ8kN
9gU0xJ1iWNwIgYlg4IxHL0G2o0Cy80vqiuiD7FYA0KryE1EdVhp3DuMAdexDB/423358YQNoDMl/
b8bc5Aj0gVY99L1+QWbvWMNKe8iQQJ6KaK1fPKtqDLKpF+ElV6qooBKc0wN+l74RtMn/6BJVURRY
uv3oR85DGpROI+dgGH4aIqyt89OZHNCqdq/idrZ+CfRWxo/wmcoGmZqjURQxxownOuVW1bkkGSk4
FSeREt5EuO9bxGRSjwnlgBlrZbJ8wg6h17g+Go/HhuOOD/KkQq/+Pz+R4OXnILZRoxOmwkv/s97Z
x6/ZQn4XjNLZwA/uVKzTa2o+wu0x79g3/NuZospOMYnuLJ4CQiwqTElx/jGtVlvA1HkVZyHN/p5F
HFJVanBxgIcC258CgKCFYvP1jRpVwvukCn8eUVwmSmwwDJWI7Bt3E5600qX2ximJY7tGzKPNEftr
dESK0txrliPNBNphainETS61xJap39G4m1awTWUx8b1PhDLB4OkiqdON4ZntGh5Haj/WFwmeFYP4
FUY3zgsn78jtDFGI3UcRuT5IOsONWq40L1INlwUNjIsNgZnGcga+dRluysuxNPAiuVLaYVrj9M2W
5R/SofXtGzvzK8Euio88yXDdpOHTct+zyQRwFZhs+LctMBcJRu9+nzIvD6N8HCI/eTKAAky9AvZu
zt4x5aG6xueG06lut6jGunHY4IJdyg8nlQkqWndOqztF9vS5+l1pkcysyZRTChIu9gXzHHWEmgXN
FgbqssQeOeBQRiZrDkeKuQYam7/pDE8KpmOhMAqMwOR3bt66eps7Pl6eIWPApvUodFI3b+3kJQm1
Noyx3Z+HVwSj/fUBTdfT/bKpaAte7rl+FFxLDGvt2WszBdeENIG9BgvL1x6f+YkU5G90qcNhoRNK
pAr18UN9WsiiCu0adDg97R+yd2G6jjl9xyNQ2ThlyGnKGvrjX4q4Xp/1C27aJgwHO3sI9R+3hu48
fUsn7gvp0AJZkS/7s1cGz4wFBBx3R7mmAy11I1pK2qwCbXyKHvl9+lN1OsPFRE5ay9DU5QsGtGxj
H3TH9mGQsZN6odw6d1/ilewZru0V++03PIldIBQ+hwnHFriH1oZL3bksz1OwzMzLNNfpI5P1mmGY
D6Yq7OxriGchPYioK7vq5mCdp/FZ7/H9eJuAVG8DzUQSR6l59JxnEx1jbNLsyXxrNLDDOa3RjFNc
lym2akxoaWBsRRW/2XRojvuQfrovuBOs4ABb9Y7rgj9kGPDq6yqE6Y/H1X1hNeK64M6Jxi8lqow2
xWd9Zc3aav9DRwa1wyOiirQ/U2F65GC1XWYr+T72z0i1ILyLueJh50EedNLbm7v3bbi/flBW5a0M
RPgZiyXLW3zvD1RtKsHEDxKYBao0dJalzAWg7hjyUqt6rRkb8sPcStTcpGiCcod1PEtxXQvbHsvQ
Uc6+HT6xRjWnNcdNNkOmGUp3WDuWN5GXs9H5AbanX/KEtDWKvxj7Evus26CRyGsjEMSCW1DKcSpy
Cr2M6mVbQ4dQHzHhIi7vM2fZqbm+iOehGJ1lot++UELeuD4XPeRMMJis4ykY4AdYZu/2pGtzotd7
RopOG5iw9yrceGwnwyY+hggERFoP2DdTh9O6iVk/poqlwh74KF8qhGfx65jhHQcJfDUQrn5CWVIi
omkiYBaW6BaM3QmoAq4jjR16q5VzFi3ZF7xp5doMl55PMxe0MtgVLLfF/gi9lfLyE0zU/+OOTwDv
Weg+27m/YE7D82YmXxW8F4vZqSKkP1snnWTDJr1GX1Y6uhTMZUTOoBquBizB/4uOVBaZe8tGhD3+
bT2KONvvCRrPjASFoeHj/qAIlqarM4nrVoCJfHMuDG3svoSjdz25i3x5narAJ7rg4xySR84HVrUp
q5HOSInhmV98RbsftWM8MedN7zs5itEpLKoSTKK3G7gbvX2g6bEDi5JsszwH5PnZV8S3DfNVYJw9
hMMVY1NosuKUEM2xFOUHFEZePSmR11KX4EAY9K0GBpj1DCicCtFh+glJ+/2hlZ9KePguCdeMtdLY
EXJiDZZwlZZoGM58RtSbmmCo68kCR/0MEnxPDpwU4h7z3Z0dVZnCNnkWkPGX6gED00sJ3spNnlnv
8vlLakOPYbRPKfm6pDKnH+4V5SZuCH4ciuSVOplLM1GmFZtRSBsd9Fnxgm/msnqp2Hm/0QXYjkWu
XZBVynB6G9T5NySFtNFpDCRq5NFrdFylyg+rPpM/btMEHU2QcMmWk5NEBpLnsmFaA3fnMbnZsjVV
3uMV4H8oZMs0E/LE3CXkqpxETfJ9lnKhELjmreom6GB/emtEL56yCjaNPK4kOWZ1l4OzgnHLdxLb
o7F3nNxTAFv0fg9GP+7YfA+PjKvuwnO8pw3VrEu9JVs7NwucQ5PIjOu01OvwWxn9CSZhT611To1g
HGizdJzWHR4KvfE9pIvPHb1/ptaetSNQdTH9S1r9Qkq0ZNiJ5CYYcycUfG+jk0as8lcnZBR+X0ZA
3u5DPnsIyLFhIvKe1HWKIrBHoKTKU10OIEhOrGcpeVpu4IMwwBz2aKRbWbqu/go4xGoJY70kHdwb
0aWK8/k3Du5Eg+wK8g+uuU2uoqMc9pcl6gb4Mgkrwe6/nUrgzR7rGaYAAApBNoPeCCYQ8wgYyjOj
oQX3tbItfWodvxsFsPvXOL3JAxZ6VMxdjdcseBPcBvEwc37BeRLRSYVepIP84sfQSf6b0M6bFTrr
KqxrRVwfn5XaLgJfjmdq29DOplkost3AooI8bkUNJfmeuo5VqeTIqry1m6soIE2Zm0V3ZNrXQxfC
gKTNJGyGi6H/XmUy+huog072TC7FWX7QMTxyOoKgXAJIsD/ozW4D65JSil36F4cE4NEfoMmW+UEv
g0Y/p9bBzXZhGJI/WsOkSfIBfphIdzRtsR7wLorAtCMXGcBbM/9Zo/q/PdqUqMgFrjYVMZanAXBH
sein5EFYTSPDNq93LQftAxWv5zz7n+nYNy3j3ZSWCkJ3lcmx0bfIs/6g7FzfP/B/+uClAPtWXNNa
ntV35nCIyg0/rGymIrCw4msgQC7+4QIc+5hf6gn91LUkcrsUc831KtIzdyRr1DA8sNTkip1cTwde
bGQovYd+7rdvYw1ViXA+ZICzsyc6NcuLf+nHvvSkxH0xhCev6djwN7sTKBIL2LSyS0n/iZEkdEy8
VQ6VhsMxoOG9f/vcXKG/lz5fCgJ4K72+VaME6INV6xnn13GsWVGTjjwRcCzbOkXqXbXHVV/iqgpw
lQsllXmS3r5xQ5e7noUd+lwJx8C0MBAjQXepddIjrLLnBJjSqzGS/4KCYAG5HneSJxIeU1yOFgao
MJERY625lU2/7ttx8f8wCqOTs5VJy3of5ehV2QLIRx6IH3nOVv1Pz5Mz2Vg50j6f1uI7dVcHy8pY
J8DXTj4bvuTR201Pu8jzD+8DWuEGwl3PFbVF5BxX3Z3i4glS3F9RWk7UOq185iMCXIeGE1YeOtvZ
5iuAL9WC5214ZeohjCOda5ue9WYt8zuXUDemlh295z8C3C5Hg9A58/a8DFEYflLajiDcHITajE/L
UZ77FoP3vp1w0y+fVhYVSZ3tfrEGwtG4HH66k/oyiLs4qb389jk91haF0AT3o5INdB1t+pr1Gb68
lOVi8SkCZIyTGsC1jyArPzuaUylo4NsPr0WGvsDroBJOzZgYSd9a3i09feuCDdWIvnrzLNemifuY
PjgsQwGOz+wKqkISgzcKySQiC/XUUtMUNtYtiVy7TNGTp4gSawUUqLztX+la1OgNt+qhmJej5eqE
Gt/glO3G0YfQgZ5Q+0wmPCqKc14sdqWUYm6t7AnrXZ3Xs/soUTo8WHIy8/nx0KetsPbaCWirATJj
pqcuodxa2xSxOqCARIjVcfN8JTVTVsOOlZAqIs7AW1b3W7BRqE5v6IgDmuj+XiA25EZHZmBAHvHn
lkCSwRC5nem2+cf2cepOBsSzdRPGobrUic3SDaEbcZlf3R/9hGIl32mmfJUOOeeODRDuY7wa089H
ctxIv95e/0twYim+/+yH9r12yG6wObRM5d5/CxU75lcocOAov/YX9e7Tan3SCuB71Uh4E+/Xa2DZ
m2d956UE422GH4MP632QKi+Hlh2HCpKJP+aCm7dVkvmsy5K3d6cgRvYjoabUNN8UoFqeAmnwxrJ2
iu9lSErV8H9Zp4TLA9G4eBFKTy9t8qqjvDOY49keY0XgdDeaO79pPQhzbcKx7y9AYjHg+RSpPYUV
m3rJ4e8Bttn24q/ocD46eTiFKMVlpGUyP1Mzk2gGEzEZ5h4gl/HGRKJA0E1ojQ4dHUwkK7WJ+8Wd
cV8s+RkVRyOrsxYK/SD0YeRzFJ1aIRrH61kFVmODSvDr/Z7TC9FqUKkqyv8vfJP1GlrxW1BIRrPK
d7xxC84pempj+PgkBXUPMPFyxdahF5O4vW35iwFNJ8iYBJqEdfRI6rSu5npNnfw0zNTIvyaLL5mu
RChJwoQxY2ItUzxBR1y1m08DRwMGaz4np8KX0OEaHmFatkfcyGShUVysDpTi6W34JXmZqXfvl9aw
D8D7TvKiY3Z/UUad5mwLr7ymHOLaWybJcaLfoYV3k8h+Txnlu+QAAEB6DqUThCfluRv9krXCJ6CT
16g3b5VID7NJESkEd8hm/PQEV1e11DU6QoM0z0NjEJMKKuqMS7+YVrkJW4/ANtmZWijiD/mqMcr5
Hbx+n2K322mLng4FqaD0RQppc7hxnkAVNMhauhH+LgRzrHQqTZ0zf+o8ME8kvWCZKo4UH9FthBhN
rScckzFjyF29+T8ObPEzvM0fYkLpuOdXKtU1vfh4VL+7fSki0urwVW16p2WClHJX8cypYsVPlfoC
Tf5sc3fhrWhRBS+6UhL8rVw84t1kRS0RK3K/4E7N+4lC/8wWhtXldSXR53hNLwcO7XCWdRZ81GVP
XRyiM83DTmTqcoYVU/WQn1pc/t8ql/G/BJG7b4fEb0WtaGx/YkKMDpyBxKfc2Xo17G/0RhvH7ayD
qzI9CGBDSb0Drhg61YMBUwOLTOhetlUwrn75JavIo34tfJnxg3yUZPCTAOYYX0iHOJ7aE984T3qs
+1Tgixbr/J23UgxbK/0QWUnlex88mZTRRJ0byymlaAlHVAj2jTZJUlpes4AJsSH1PaE/L7lVhuRX
la4SbShADj//fDAQ+c3VrQo3yTc0OQ5TdY9GgQcm6nI/qXPRYwMDkiP8uTwa+GBTn7JNVdIY4BNH
VD11obMRqPd3m0gIyluAuuFcd75Zs8WarUHSO8GS3WkKEfd+pvpEiJ8GBOtcDS9C7ilwNKOGqtn6
70CsfRgoCWRlmXwmgnP+B+kZQ7oPt7kWCsXADYj4/vVP1gjd4ZuGzHLZktKIDUvTAMuzz0NLBUBN
/bh0XyvEb7xN+EMMi+vX4ZTaKlvwj22Mhpf8gqC2teZ0c0O5UA+mjC46fjZkxo+v3mIbcJlgVR0x
vRVhEqIqXC4W69DZxtXpXzDw8IIbYrv5N0db3w6UKYHjGJhJ8IycldBXIurIPMSFdWI5w3C369gr
NLLN5VBLq0SfkUOGTW70ql62Q4/Frq9sdqTE63zivaxx+ScEbwLbICJrHXa3y4TMbpJOVQOJfCdt
tetfTTh9UGJ/D1NeariG+dfylmOy/f9w+iD9cxvHDX0iBYL/6pCFp2VECEb4O1LbUDLrEirz9E8c
qYFHoAmkdX7LyfSzNN4tldsY8aTvRV0HDT3Xi/Z6+yWP6LpwXR+2AoiDmuRui5NpFniH40w6uHpe
JzAUlMOywgOapOmN1z3coyERoV0IUzFvvN1Zw2YVKl6RvOitTO/JFxqes0kUkUKwwo2Jcwfa+gKF
c3qU7gxYmWbXwzsSAGTVepID1nVQYBFvA2SKk1VmTC58o5CStLswwh2Y/zKtcrFtLWLjDwW3aRVr
HGi7smd+f7AYAf1gTnyvdXsE77BzTLpPq6+YR/11xYtGbjWZiEzr85CI3tm5HL14goy+iB2PJMYH
w4HhUSC0eO31Oe35DXYlw5oxxoYAMV5GMBEs1zBK1wTvHOYSA2SwPB0sVrHGInkg23YRjzgoyesq
kTFiMfvLKL5CSjL8vwj85qpEpU/6jajf5cGawN8Zd+vvVySBedHbONdqFQ0U6hxRb6T2tMLvn7ZT
E+If+/+T0qQzogG+2o35w6Uq3/UIng2AaDpLJIWDYDfmS5X1H7JOlCUaTwliuBvzsPV4iEV0pswO
Sc+RjKZvGjLc8gpwVNs6E/NoazUMkcngRhn4Yknjf/p2z3dy6wB+92Uzd2RIDKSdd8aNusHaDTtG
vktg1VPp4M7XXhHt6davhAbNJVCR2c/NuKKJuKl72LM8fmxUoB2AHjSLzkjCmtUN84rInDJ1+Lny
CWfFLGMmuC1B3/mBeH/5b1KSJ+x/lo54xuA/YOaLwDnF/n6L1YZEJl+igTMg0pxGEvoJ3ahrSbWy
Ex4l+C14ftksSidVm63N2x0OPxIeBEkQzFd8zW4YmrteZndjoIXrWoDe2foQKAQJjadziRATkJck
gpL2y9wtt/uGIvzrizaSpL7ivU6js/SbXfFBCtMXLlpv+2gXwRJ79MFufxKJsdiExAho3Hh12Lad
nIqx9gWO8OOn75TtFxkus+uqtQDQkfT/w36wgdUx3YFZyVhBp7EGNp2VkIMm13k4+L1uiR0EQ8kT
YAbhZBEQK9+yivPstvTm/UbY41tVzXAQ4qqHp9LJD06VE5aqqO5w3bU6eW6uCriZbSLf1Ld+SmAv
r9qtOdWc2LKD66CoFwdec+wfgMKTy9dhykjySbMx6ijtcx4QNplEQ8XpmeoLUvkboGqLk24sk/lY
OvJtEyQUkFP9rtFfj0uinrlvUO/7UueasXWhBRyXFQK18F7s+K66bcNJV2sbE4EwM3Zb5bboDUAh
/Gur3zasQybKCzY+z2LEd+sp5CBig1XJ4tjR851GrzuJ6rXTibFPxUfgeNoKjydR9sU1n9uCfazs
OXO96Kc6lGgPP7aHDXrx5VFfrxmi3yFeITAS0cY+umznKNy/juod+wbH+RXxGNlo502f7MH2y7lP
68wEQgZ1rE4SYVpeJ0aLIzDIe9LfEAd+/p2Ydl3cO7H0sITUREWpvqd2vTASQnTYKRpL6v4pyudw
4v8pekxgATskMWf6buCTwLTqyQmBaYhTt4AxsZNlLteD2DpGwJWYwY3ooizHQ1dg9tJ0I+htTmHJ
f/3euSAtHiKe69ZqlgbiGjkXl4U8J5bmAaj6SzDtslIvBfpLrIMTD0XrMDt9Xi2iuC1rGmKHmGMX
WocdXqEWHvcG7xgU7lkffnsTdhGp0UtBd+UEW1IKBWZubpvyatZ+WBjlsKHCVOmFB4wgmWLPPIci
CNZMa1Es1bh4eqeC0Tg4GfXCdvsaxdlD/XYqvrJi6DjmOF5DwQi7uOW6XTK0AbkxEaGcIGYdjPkR
jeHg6yrybS5fWHmlxliL84CgRfCa7w8VI2at45bRy4SPIRlEC+Po36n5u+zfxpgVmIdUTvZxa/On
TBlrNu9D+PWL7AVNAaFpo1wQ+lB3c782g/m1CfBwhGP0d97qR9b8wux325vul0W0M3F5sRKOUtmq
X5nnku++lRv4pTizDDufh46mfHdxyRR91bBvQOifUhU+Vkm++4S2rnoRG2P3bV9yTLtOhX+nmx5R
FxzAKOD89DwAcSwORuKAxpw/WiDm955MxdDjsJ64y95dVU6HXi6n3sd8wBJIT3nVUyifNrtgLuZr
kuG7vm/FRmFleu3pqxrnTmsU8Mr7WBb+x/6EAN5CpmMgVJkJtKoej2bsoWjIXnQ5/2G/3LEZwexn
6Jfyrgas2EBgG46XqqoG77uRNlB5NjRo4tlHnCoNl93Ls5ZgBxhLX41Id9G1U6Oz0IisScjnCwPh
jtVMwuM5lO5LMFpbfpoHUneCUH9/Dr9g97xtQnuOOq6jcrkiBsxBdtkNoaXZgg0jF0JJlSq9HeO0
QGt1hzoaLpse1Tfkwr6rAzi2LfWwgbJ7Bktl8WK0mKCo6WVTIyNKI3rVZhk3TBOMuw2R74YmcMn2
yf9xOtS+uzeAqtNJS1V0+CUU4N3afBLI4Dt/x336dh/oTaGBJdNVu7F4z3o99Cf5PffUUgNpM6M/
xu390CmngJm0KnPwzFBrnfYS4STIN+7dP9WF4RPCABjIx+ead3z250NMWST7C9OWLt6RhH9U9hLi
YKlZcY234oXEpo8SnL5eNbjr3Atac180FH45adWg6zQOy26MfgKn7Y/FkpAJ7y+iQq40thuq6NTs
k93rQQsDTk2R71JEN+iVe1YgIK2gXjaYISFijPHMxgkCuq2CN8aOYWno3CebYW0NLAFv6cX6aOSH
DYHKbai7KorgDe5Xw/u5j7Rf6UBtR1Knq1vcAJKf4MWOyvkTvq70tJWR9EFyWxvG5VCjSg0tWKux
8cac1abHbvJ0NT5+c2YA+ts1xxjlwGRyThyd09ifKk9tUYQ7xR5oL87kmf353/7ZLYGwafhYQi25
7pA47R+s+fj9WNmuk5HAf9DHaGOk6CtvpKNzkXt7cFyYlej7R8qyFYsoPlS5WVCNiaX3eyyqnGKK
ZeUE5hkBQQTH+31CRsGhF9dU9qDpdEcxLxZEl6RO22pwMOQjatG0HYEH+nkt4jpKICZea8QzT/h2
ajoNZaG1NLi5jWvA2EyhlJ6Bf86XAQMxM+MFumjMIrgQb38MK7IXrtjv19DhOAkNtQLHXUhcJDFk
+J+ARR2+A1x4n4mdEZUVYWFBemFSSuaiwzQz8VEztZYCVxuXbMLq3w790EItePzmK02hAnt99+h3
ChFJ9nkG6l3fh8PyNz+B7voCN7otQk66X8+ArJAzc6kTfasRfYsHxAvFx62WYssAUzSUDTW1EWP+
aIXKZ73QFp5Qjlbf56BJQvp9r/NaYJ7tEcQY625P9MFmRJwZ6z49c5Bu+hyoxpzJv/Nd7unWNnx8
O1DGB30H4SC96Veg3njBOwxGY+Tl7OGaEu8Kw7119izyrEJRfvu0Fx+9KwwWqTZEiklhn0K+Aep1
shIYyNwMVagm6G6WyHBQMP/L5TpW1XvUZ6DKFCBbk0bVCSzwKkTZJO3Ae3jnKn9pE6c46cqUjnBW
D7AfMUMmHq/GuKnS1Lzoop4FEGjWVzT9HyyRaXCcvpWujSD7eyjmiBOxdfNnOx46fA9dV/zDbkmD
yiUGYcEpXN7Cg7cpE+V868vg4A63ZYJdWVnxUZfX9pR+2ipmUPS2BodNdS+7b7R9y/OY9fym9Pzi
xujOpeo/j81TXVUayHvjgkwRF+ZgtCQu8+fkvYum98Rab2ScZbZ7jBuFN1LPhViMVC44kYTDvO53
AQwc2NOPs07wk9IiXKOugckOqUtneIcisET1TRBJor2n1u565Xs9TLhQxkYp75SNf48OgvvuRtiY
MdxjKklmXMnns3nobVAcCCeLPxB6cV94GdhLN+YW+stZeeuMedG5lKeCV8sNkWM94l4agQMo1R4o
TV8B5wkbvggkFmvoa0DBXWdIwehyQNrqImKAx17jSgorxtZ2dcFBNHRJTs+svpM5JI/wTjlQcR4G
Ws7FpC6vIU2aHdioPTJxoZE/AsRrs3xMZszugZZYIIrPHbhKxkedgk/SSj2cCsHjUDfFv0sMFKWv
WB6egvb+K84p2VGit6R8fXUc0dZI/vG9V5XArhI/dAyikPumC7i3zoMMD3L/TGhrwS4YIEFxdCUN
ibKtyXIwVHtyx5nMA01iEdFdMb4RcWw8lFvsc4HVioWcp4UOFu6v1G/wzYIbkut3m87l9PjI0/zN
/WKzmu3eFH7rVLfhYqkv/SddVqfiBC3ehYdqy1iXlU0zoQ3jYzS62EwrwB/eAzI/rDzzt9GWLgcW
SMmkwBwn+AuzPVouc3eDm9GOw6rSYMK9yUFgCW3V3dnAYzTq1gGIZRcM1GOa9GKY0yf0YFU2RoeY
bwzBA3pJuXcQ51orZiREoWHvL4H9B0/Gtd6CT59RFSV7TvqSZszlO4OWGxb2FHR7XWilaNZn55O1
BK+r4iRQyxwygWgYKFSWPjDWKMXH48XP+vlTq6UM/SSwzVejfrNggoPq7iBAj83/YmcudCnc2w8d
dd7GFq7OMWTnOTQfo3FzMbFkbaKYCIO7LVsI/ZhpBqS1F+tH6mLiqN4lWngYKeMMPhEhjtxPyjiW
23ge8LEIeeN5CKIU7EHIFzbEcKt+971E3B8x8/8mvvInHKSb4msn515oCuMpHDdFMyQx9jDKDQsH
JJPCVv86uei6PY+hpZZM1sBO7AyYxJA2vrCsk2SRsUhRoKfxAZIIuoHcB8eqUENCSsZohu8ely/1
c2/CYUGQNXZQ3nCwO8hgd1Gp23P5f+HbvgHalahIkNf+0l/IZem7rJekrBqJGKETbjepkaGGoBYP
Oy9vgYd98n4VUzkVrjSPwbQWonyPufb6Iv6yAi2oDL2by9wOpDyYCO9gTNw6IuCrUMwsbE4rbBQ3
X/rv0BjV3HKXjHO3cxKjSrtIoJIzZleNfU/SAZSzeMIEGpJxWCJI82m9hquhL136s+fGkBRMRk5a
sTYOku10BGu5HtIIbZ3+tK/ci/cS//sAPUYD/rpIFUoExAVnTbVY3rGkH+BvkaDzIPZ4No7VwGoz
rolsmDOhsWeyZmgMkXWM/EQBuB+enLv6wiJu4U9AXtJnlfCPpdsCRurvLVHczojXkPA7I9HMM//Q
nSRLG3aaVesW9OkcytogItl/SgUTwt4ewnPoTP98K5A9iakWKIMvN4NS9zqXhZ0e4/KAfqCrw094
IB5K1+RIK1kHCKddGVBbuVmUmSk/EfBVBpvdqxeRW9Lps9fGY0pWvKT0KmPCHkpBZbMdOiaM8x98
JxkgTde/lfQzqFQ/kYUJPXewGD4IB3o8Tbk3yaf9Z7hWlxuJzUM53kb0L98eCXDd/3jM4SGYOFWX
c2LR1UhbgMNqxzQjEjh/7v37ta6s7y5fzoCxnA7BdnusqLawARuV5suwuMHwHjm3oonohslhNLem
yHuaik2XX+3RwrJfiCglgcg8mEZQ8gVb2qBr5oliA7Yff+MWwCQ8+r+kqgD12pEQ0WMiisKDtNwK
MVkeUHk8dj28cQ1VYVKce0YMJrVxKvZhKBg2Lidywl+Os2Tj5QulHVe7jtqniLmO7lD3d0n0xXq8
qRSPjSYQ4BdOzPPrRtncKNuYaneEoYOeZdYW5PnZJf3X9uLE7t0uACXomiaCd9tfS8Dt1sH9qM/A
9MmQuwG6/mjlAmU+lUGAJNLvctZoCDKx3WqhqVfBGtCdsgjRgrN2r38Z6rfsdInybm1043zqVH/r
2mCI4fCY5gEareZ2E0fZz3Y4B1G0xg69zhM6KHEuqPfpxBgPyjXRWB7tDGQDCyyL/TZz9GTiZyPu
FpACZPuu5ZkUMmHP4FtGIEgYyZgCUu06j3eLiakNhOHO2PHZtaqe5hmpenh/n6KOhe9rRwytznvI
vRnWO/LkEfUjO/M1CkGQBwBfhDpVjFQQJvoWdCf4J/4mVd1oYBjJxwtWhwIMET8Dpn+DqxrBN5Ie
BL9hdewKkS+tM6JkgiKJtAhYergU3qF02Mk3KKg6GohUY4N3YlXMmShI6E5pY+Blj3Yna7bSoBHC
rUrvWDq7CDhGkQ2qSg2uNYHmVKRRSAGRfvFxWwWvjcWf7A1sQh1bBEzWlIJL7PlAWaaBG08Thhc3
EbDhBwTzXrsHKRgEjS7oOexK380yMGFWUgQlIYysbeOZdqXaonCkZmMngOwoAP2Btem50gNH2kfa
EIzcYBMyjnSRd7723fZSqmwdEbbysC7F7hiY3oWuNQpBioU/rnYrsc0CJClwAf/NuH+aOk7bCjXr
arrG9sfK9OMN41P1woxuprmVZ1PAq89BVfnK5J/yZO+RS1/tpRbITC89yu7YcG9hBnIXc13Sg1aA
G7wPHS67KU8LUOSiA8ypO2yEE+P+w36TzyzQzorwGmHaADJ3wO8e1Oq7nuk0oLvoRyb0ZwnTHNgN
1pVPHimuFdb7cyAmgDSXdURVp2nY+6b3r6zzcUMk4bpC7C9DkBHpaLcBtQ6fzOl2LyrWOEFX7BLn
d7mROdOSCR/epGA3O8Mocw/6SA/CyjrXl2+M1mUSYUhwPazCriZY3rR9oMzELSayApaOBFeSXoW4
60zCJOsJrzyorZJz1CnGkyUhDAmletKpsKkwDkXotI7D9MUwYv9wFishDMRfoyokEbDL1EOp0dPx
NjqMXtqRsOgNueGRryY4XeLdBe7Bx5gMezhoUicu3Ezv7L209khTyjnJnK6kFY1AQri/0I0Edsjl
662U0Ije9fisllsed5qykRJONmgUHJbggxuUBt1jzidXJnDHQNbotEzbRTjP1aBZzLsn82x1m1uL
s+JbhZr75zK7FMCA3aZJNW6FDDUDz/yUzahBs3iZt4CcZ+93ZKVYpxJ7k5xg1ctS9vm7Ymy1HHJY
DwYx1w5ABr747kCB2xHmFIxeHg4SioeM+c1iBvNiyNo5LBvZMhLYRQ82iv+6SJiyQLWiZI4hp2Kh
0GzdbvAL0GJsIpj1B9hwiWeesUwIIf0G8+jsiP/Ooas/RHW051sJb+8jfQQiLKyrbVjlOr2ieBpl
kpHHA1587tSc6Sz3unJi7Iol2sg8YI2oJU+7oPu0TqC6sMwetVXD6QVIYbhlG7taullfw/K7C2N9
2r/20V6DQxCdgGCW7DmaGufHJlxSjOjsdP0MfbgOs4QeHqD60qHXXPNwE+3uL5wJmuj7PxnLms1k
TYVZ3uvj1BmFU3wz+rEayMQ99esD36AvJ7ZBZDjZ38hiA8bLsqt4iH9nnbtiJ5JEuMhFSzPd0lCJ
8gdQBSUQ+bEOEO8V7++VGDzxxjrQ2r9kmV+fGeFAKe28HERv/0tQs8nPahFeL479D2VYRtr6WOTp
r0jFMJYRdXgB6r+3+6URNhCQIWp877R+khTcFECeU6gp7o6E2FKOqWihxsR/GAB9BMXsz3518cVr
CULsFOM+uXGlOJj38U1eJHBAufXCqOs1S6cdGN4PgCjP+8kZBfPhiK1pduEB84ygELVYXZfxy/4P
+HTkNcPoe0MH60iCbnCZzecmnaEHGfY8myJShSmII4GGphie4nG+QIIRvFM3/hZTPUBnaHzfy8bQ
RsOjB3WloIvP23qi5CXyWyIbNZq2OS79uQZXHWzosohwIWv/urlFALDrFSdaeEkkg4kK6kHvyo/o
4KprtRjWp1dQt062vh191L5W0OkM06vOYPHZH17FFJdvnyViZ+p0LEwIXEZo6mwGTyk1vvp/jir4
QReiSGMvhNRxmXsYqKMZxluZaF29akTPTPxE9o7TlQWHFQ84wp3EXbxTo/kI99xeVjdILIKLOqfj
/guDic/AhCjStgPBkFOrGjm4mc38HGi57XzFUxjPe+3PYp1EwuMBf2eyQU9UHuz71kKS9v6BzYQn
B3BRvu602rS0QPkWZR8fq5EH7UZ6NkDD8yfA5WYFXZyiDIDchO9OBq60GLrmn7bMUXXyHz03JU4Z
2zAtb5uBIzKYcWZFo65lpriVfMa/mVAaGS5pUOOebSZpVP5R3xr/cs+ZSMEdSwYnOXZfO8L4dY2S
r2tqvyltv4fJMnB1Np6+vHzzO90kuButw3MnzLJwIPaAEplQfyxvCWcjOSW+Oupx5hY7V+GaWoQF
R0EV28QaJEfXgFp8ApNGVOVdwZWLtl2euwUFw10aIUnipbVtX0lM3pfwnKsgSBDRkEKuoruSJERE
sCNnHKwY8MdjhrFrHGlx6LY8cYP5OnmkXWcLKVucatUQeBr3WP3bqo4B4LexoHlk8IKydpMdN5ZS
HhP+uHYelbswYt+ynVSDDChjt/UPONB19ffuPuWDZ0hZonnmxX5Maf08pgvpF2YhUZg90gEVRby7
oDWMKy2MLFJBfaUM9DPeb9cYNtM+N02v2mgel8kRGrKTjsNfadapLtC4yZSQgVPogKSJQpCBGo7a
rKl37NLDC8fgeps1ze/l/GpBAtDV+WWfX2UU4MtrsqRGE39z4x63alscREjEKcVZbgvamZjLOwDI
FMCT+4Df2/alKBBddykjMvpj1zgNmtRNbGmvMKgT4v/zIHnwS+ZSBnAY3mPw6cIblSe+z18UDgIO
v2RFzozDg2h8FJfWRLL2D+OfDapABl9Qcpc6+YScXQZEEQA6RIFv3wG7xNppR4xUpDH8zKEuNqCM
idgk6P/I+HACW7MgM6ZbBeu+tQYLg7v56lwTgAvX/bhgZcsmtNKVCnigq/66tuf+qhx/RRtCp+8A
VcLd7ZSEML1h3z3VhgdqlHXFgQhnyDQJBp3oUoF87pQ1sYLk/dzzZh6vn+SGOXuHlUgYpulkWwAY
t3ugPQqUG1TXjxcnr3aIA8kHwXsb+3l/Se8AA9JCuNPl530wmBkaQj92p2DrIOCHRtMnqI7xV6ux
abMjuhN4xJEUCShkIXUrKqZKIkARSZMkk0uRqq0Wwn/Coqrew+/UqUclvoYy6pVFOyoYtrdHhTEj
iv4S+S/OAPJ688EDJfX/c2WwN1iPXkgRPU4RJsR/xzR42hL/4Jjn1NjlUmZ+Y6hTRalNZh+XCb5r
uQfU87oNsQIfC84zHcT4LrFdcGilQouiK8BcIrUielF3WGuV+SqeMUVY33mW2+fSqaA4mi2MmBIS
C/dAeaQgmxctLFIBvhJw51BgRRpaH5iM9Go7z3JZtebiO4WggVhsiuJSprFIpFl2pwgdk6x7QhFK
DfSWWtkXlUtUK6QrZo6dEmvHr3/LBXWO6H6Y1x7HR56zRpR1+o2OZtSlX6F792zI6+CYB5vI44v8
PSz6HGGvkOBH4WpI29OQ82YRXvMdRnjTTjgFOBMJJ4gR+X/C4Oq3RcR3vz0E70DGnDbRyVO023p+
xdxg9JC5xnA3pSP8qWkhdA2FodPoHeeun7lIaJg4cEHV73lzOdVgy77m+vGAaoNCVgJXcidfZaLd
F5KM5kyez552aGHV5tTF2r+TkkhtlzLoWqSEXKcNo8Lm0onvBOEzB6JeNt7aqlSnpkOKo8uNF81H
7d7zWW7tTlrBizUWiih6DQbmpfU22RSlAuGHHZ8emwP1JCjXEsy6TLlZH8l0oGNc4BQobxRarv/w
1DlXeh1PDahwpcxIwaVuW91CRjBpj0q2Ef8Xz8RiEpqaGRy1ugERdIJhYOfOvq7bL7uXgSCWhbGk
M2U4viuDveu+aE8KBPB1oW1pNNw/gMsC2dWheNfRvPOu6xDK/BQyJeCceCGwUWE08Z5U38nwT0O1
/1oQlLMW9QJY5bNd1jEt6Dcj2/ygZTvwXHe82N18V3eXZt7HK0aEnXoSCdhiQCRwzX1Xv4MrU+ME
sVB4C8qlaa8kApJPvuCyPEWEc9tMmSsdJv7lNG0XBEEP8Pq2w3JXSuVOAnPYV/IAztsLSuZwRPrP
jNQToVOWdyKiC+IoSpUVc3ZlEDfGNURiX5AbwK+4/0Ly4sOklColGItHXufR4Hq20lFU8pACzJ6E
Cp0XCh0dVDoaG2pq7VqUjKD7xRLdqwk3PxY2fSlP0aiPARtjIS22uWQYX6SQR/yzjS2HSEfiUuF2
Z+VbUAJr0Ihp/dPm3uQGNcAhC6QIIk6UrK+IgE06tgXAUWCWrcGUjfPMuQfoDrQgzz8rmD77498F
t4wPbXFnQpjI9bcdRjOF25nWITN4+Ded5spGr4hohl5Y5+hTCwWtomkWQDknf6oIhkKGhsk4nV6G
SqPIEtbh/qcdY/7zz9SSLt6d75Dpp7IRF+4nbmLgrYJdDCCVTStJPj0rBoBVuaMK82xFFvAvEIBl
BBZjUih2vdq4FJaB7L8npMkXGSxjsjOul6PDIRoOQZUeUJmTAiqISjC1EkUmCrzcIqk+AnLde5gJ
t/NbhwbLQgFJRfXrj6CV3fmIDojcp5YZ2OM6TtyX8LbAGvjfLj4QCAO1MgoUr2GgfXuwgE85VaCB
2ZjI0MB1vxqzIvJTfD4aJuvmmZtvWTIJMRZZwNCA0QrbwqLdVRZzuKgxxQGp6igfW7Q8O8gCm16D
eJ3D+B5q23moJM/5K9a12Nir/Z1x41U8E2T2mqN9ZturHQTxRa/JKlOVjUPk/VPPpzqnuDVy8sAK
q1EWI4FUkeJlgv6CJD7akHD1ELDc9XgrLIOt9ETXdBF9PFgFraM1eNqA+TvAMSl4TEBrPW5hEZCM
Ylbvl4/P+XgB+ooTNYM3svEA02XeWHZsJ/pG8kDmVcjLTlb2NulXK2OpPiXIEY2EZxJxqlnd/80e
qUyHGd69azWdhmMB+VDnbqQ+Ut2tzvw+HbMg8/k/rBdvPn+wCWUblQn43gu2KALIs390wzFevmHM
cxv5Uz6HTnqVxmKQE4WO9swCJtdR9aTy9wsIEFSRcH+EPMI8fDKTruInNIwjoT0yw/s74ATrF7Gf
sgIqvqm5FothvQfdyKPPkKPhPmBto6fn0N76FgWB4h9Aam/Ssv+CxtSTfOJW0Ml4CsnXKJSBVCRi
poj47eAROvY6BUGUw4iWtlVPehjvvpAWZfoZsCvWJsl1REjxO/cNTDmV9v11RJyyd2IKbSm/bjIM
b6Sho+HtoxSavwT4l+16CAfpkpTzZN0EsVTq9jzWeA7g3BU+TnwwgTCK6hp6ZVCG/P0Zqt4Jh+8U
4t67JEXX+j/b4S5IXY35CVTa0IEsv4p73+H7nB/lvTYRS5RuQIfBCmjqvOz4r+gprP8SOlLowXH0
Mt/GN5L0oJzNQxVqAYtzwO5TCH0PzKG7mNsGip+1y5xHEgHWtymwUN38ccJUQrzQkIoxf9cjPgux
MNSSUWPI4xAzhppAGnN20XiKC0SA49/2ooRcoFUij+Bv+SiOVJ/ztvmGupQDdOMIrlGDTSzHKO4E
OFmI7rt0FV2cnT43NdJTNGM8ZDHpr7IYCYIVAMz0Gb1qkUYNlCGc6kMRQ46D7x+seIohkilwMnQb
gKJj7tsRpfxrhkwNCXg9iC6IcjmkujI6SVUI+hHeDwKNp6Y6kBxFLzOas9Kwk5trDo03pbh615y9
3CfX5A22bxopAXIfdywtrKGSrt3umTM7iQubVH/hIbFP6RBz0urm7n65csHgoRVXmfuQXRuHNipe
5ItWAlGQykLBPCFmu7+RonoZwhlor43cc3KZgSGu/RUA/Le5Lcto7WU5S7IdKSURsF3G0sAtByHy
nY+g8t/ocr7XOUMkpB/uNe1jNSFwZnag3EreojF2UEfpiB0XmVYxZUXOTX1S4kua/2mFv/mxnyrU
9kk76eRCFJFuRfashdUcYIHf63VW5YAiyjSsDT5Dnal5wWEI3lHW4TxUsAr2KvwizJ38Z9eW+8rR
I0PMrRd9YI66TU56ZtV4zhktfSThE0CJATxrbTBMb2Sy9Bhw+RCiFShksydWg+d+/eshqZv34dTA
WPj7dTvhcxxjd7tNRYjjfp4CMX71NKKbMuEQc449CmQ9VpXUT8mwkNwC6H2r1eUgROHoGkKMPqpM
aOB8tz5KmxxNEy3IRPoPH/yVsDMVv963iPq3wqaa6oiSOVECDMhvgDRgnp6vtNx4HgLUISSVEWxL
AL0/MGME2+tAy/oh4CvZ+Q8yILLa6QbEBFyTas0RwblCzQGxCFdQQgni61HQXGzLdv6R4v15SCOG
56Q2EzLCypgAtbemw8IxHbWXqMBZpd08Z18hASRQcCZQP2MoZYB7Bh7m7n2BBq1kNUpSwGzW/E+e
LDX/n9kTS3naXh3xyIsERqo05f5AWYSvSAYBVOIEeOO0b8wRdeHNMmV1rt7nCaQk/bl/V2fS92SP
K/lPkiRTu5wPcMp+oX7xqQdL8uvge14e/jbFWizSnaNAFibOU6Yv9NAUxaBArBF5MD8lsUFZFerw
g7pCq4T+wjWyb0l5WT9TR+qmRJBx4DGno/GSuiFKgtVb5Ebqy/yLevHd6KDndZdOi3PXrHT9stPk
fVXKtNA0aAb7QDLSot/5d6R+5Hf0Jbty3iCH9OEI/yG6faZplqZLAe7gBXlMANfPBz0xUdk+CZlC
EJXSFJQ6JnxBF7nEj8SVHEcDgVONpNx8lZIpWOajdGPVkRN5eBgy2xyN1BP8rBJeU/NuargfI8z1
qlaJZYfY6dtZXIZNiB60DmSusc5nLNuzd007Mt4MVWEa7YzHozCijsQVybl3J3ECqtC5H8ZtjBff
xcaxat5Ri/pnJq5oNoLaKOhdAhb7bDnQGREzgAG6oQH/Rs+NUa5k4APuCexmVfUKkT1yisWb9Oc+
wKofZvVGQnx6gh8nXu92rHQOdNfifiWG6MLsAq1TAb7j0bax6AKnt5fZ0b98ffuN2du4xb5LSK/n
vGLmRqNsfrixKqg6PIxmmera6bH2Sy1Pt46e7pIWP33xe2ukytZC6dO4xZ7zqxEH9fRwshomOVeT
FJH1DPRhq0rnNdesnqREwes/xnol5mV3WNFSDF8I+H0HEiixetB0acMQY3tOpy9gRruPVd7qdQdM
CVQ4XCYUs+b10Q1csN+95FY3UUqEGGIlnEn+xx3CF31ENFHGrUw7VrN+3z77PSyAPgw5qEgVNnWK
v/mmwjG4YjXLYLzFm6ll22XKQGNbrjZHzzm1xtppWHolkmWGTvpgT+GJXKYs8JmvUDO8ci6q/Jzg
E0REJ/7vi38KjQbA9TE70aJ/hWi5t8qDMaZ6cYZTVKVcLAdV4Vz90wYOjGhu2PpLRU/W1h67Nfcf
zAis0TjEm8onbReAQr40yzb+Nq5TKduW2qb2iS8xV0HVKrJSRbZj7ciglcB04q869Zma0aISNbwb
rMkTXNoMUn7fFYlDVDtf8P5vwPSBDHebfN1U1tETUeKaSeK0theCplObjAaXnsYs/7OOxoHmiT3q
YwSOo0gwuSgVsH5l2AgbnDsFlTofLXZtuaQ5KEugrPHrGrvwvG7vceJobOaYjSq8or02YX3M8Ptx
LcewPDPeSmlwrvcdeOZSgu4A66YA8vRFeJkT1RQ6d7jr6ZRByRa+1os6HXzlLpI7xBOS/2EijRcr
4qZEpdVWRGmtSxKKgUH/7EqdFsbNuTG5XR/RXT7/4nzsJaHYPWfZkUVfiRpR10LR7LJ1E4K3daMQ
swiydYL7vJf5wNKs2XJyO4wpssZu1VM1p/C1FBTWZI8bllZYrYfsVOw92lnlRk7QDArmmNSX0YdW
knJoSOd4zI8KVAwtyfOsJ8X5zjfA7+2tgG483AIVIwFXBlH0kMSu1m/X6CnVmKhwrh5qwk5FUIYz
67gr5TVo4CGSePKdUNNlb+SWEXv2pFOTfr5AZRKLWmxmqAgxokl+H6E94gVWwt7gEaUHw0mR2NTg
rOyfqpU6mLZgesoUje50VRFXJzBag0V/AadfH9euLU0DX1TeeXF5j/jEbzJf1+f3BgApKydYyZbs
EyCzGlEtzwn/Yc5/cxbbpyhlxJOyAHRslVgfVvaZM+B6Iv/S7sSa/Lx+deJ1oc+44FRqCapm3yrM
ozf82xAcosk5zVozklTeh9jPbKb0d+JLBBpvo7xyjVjbCFGK9VH2iZ8834rPQXJL6QivOdfKFYki
26D79RCizJ7n+5REWkUSHQg3lPdaIudYRVg11VjWVL4Fcm/70awOmcoCCzJRYfZdRr92GxdCon0G
Ov6Dt9PLmYGT/mSXZFrugSeNuurPYUmWFBnLLZW6ptaMxRg6nbBS7zoKoFWZ+F6Wjw2NKQL9xhM9
eAWZVZlYV8vtv7GeN6GrOcoa+I8buTbTVF0G3VwVAAYjk6bbI3WbhI8KNraHcEiR4mUMRCrwHCKE
7T7+znxE/6tm89m2SxWqdJX3LOh7BACAFH0vvBoor9UO4KlsSoF5j0ufedlzSlATgFXlIosc4tJR
uktAn8Fu38DNA/wseyTzCECiufhUG12q1Dpn6JqZzQwfllD/2WM3dDV9iTnUO5yE2iTbO6K/kZhb
DduZKscjexIhXL9z2lqcFQjivBEBSLTO53KUa9GT5WoNs66w6wGPOoPXnDAJZ9HTq4HrTvpD/+Nd
mOP46N2bJv2tTgvaSXNQZNLdwld3v8iCq96ZpeSBy1GOG8NDh6sX4MaXfb0hzqw1gPvHJfu4jupm
SF4nBFcpznaSi3aH3VlvHUWKsvQDxMDeIPTa4XYijJ9mcOiVlcEiL+kXHIr2wWBuK7xvMq80ZgLU
4K3ZsBKN8LDSyeEDwIqH20WdiBiuQbw1ZYzA/PCy6DLECLt/jB3ByyfGOdtCRqxjanag7hiTV390
TPHOxC5RJ9sKKu1+6ye8ol2Gp4Kk1MtKA8wx/kiXL1GwfHvzaF3oB27o6M18cAPz3xmPy+tQHdw5
yWwnlZfqezCHD1WOgG9vZNTtVRqhLcNRqajNOcKcpJpBDdkyTHgvaMlA5OlsFnZPH3ZtoZWRENpB
WBa7AmlOz34Kky5vZ84siy1hBxMXSfofJiRRg/TOfm8Hx47PJE5oa/l6EgmDuTYCvzNGc3iVS1Qi
fOdO/7niXyMZ02qe1t7FTQoBvtxWSCp4Hs+EPuU/n/w0z5D+ajR6Nx0sh6fOt3gveIV2Wn3oTlca
T+HQ6JEpSpr9Qe5sBhkVQ20GYYUJqC4aHZul+6GoUnZlZov2alZt+7s+qb4PAdT30mA/kr2wRi+G
GLdOiCNxQWLWvS63r9cUu9+lkfGvoUHFUx+pNq67zDS9Ob0zkoeNInJKxdlT1sKt4tSOrf2sU8Dv
bD38n0ZjbQ+6bvm7BG4deDnFljLasBkuXpP1oxMpv5sDgQIEUDpSz2MpYfqNNaG0IM83tUvN8QSX
SPlRZPSvEHX2SbkvwiNMaU6eea8rnzU0E3MxPTVBBft7BYuj3E/uisxqdfZFef0085LbVt3h067c
3nOP7V00J10toEO7BC14MiCV8TkRYFisdpeJUOonqX/4nNHt4oHstr3DX+s+0Tq5Pqxdonn8daL4
soF5zkmjQj0LpmwGGQY0N0S4BneGr+pYIgpBcaQEwWdIeowdHgUvczS1zINHQ+rjGvs1SZVXpB++
AHy0+4xAoJy2cv4SebDRs6YUwEHvhnoR6xd7g/f8QcoOR1Otxf/8TDQsCf5itgtSctQWlktU0yts
slxQiMUI/nc7vRipkegqoUKQbaOOjO8YDNu1zxtzyM4cWzQOQlIlGIKuGbQKyI649bUW/hh2Z7vr
+z/gbi7tXjzA6PdfAVEMTMVDH7UjND9BZElZNJ+0oJbNgDepKnpj9YDSuK2nVpFM5epxZUglfFdi
KJTJRaKD3Pov6FbWjo56SyBMvCRp5QIF6ghvDtdxbLmp5M35zS8hnIzvK6a4CyUZM4LSYY8Jo0UA
kKdQ10WhSXuu/V8SE7mmgDzAP2LgYTbYGTKVcmNL9z21oZ7pkQHQkE+p9jdzsXOMSPYD1FbzHAq4
GUchJ3TwxAASURZF1JJ0nEYHm04/lkQpm5Njuzhf/h5MdIroAlpt6wUYibTnLkaFM5s5UbaB8WaT
KyZzX1MQUxblPfN5w1e7Azqwwc6hKRY0DeSWRm5SV8kpXD36NydouropCMoTpAxBm7GNzGeO0G9a
4HmLfA92D0U0dXlDFJrXl1Lgt91sN9isDzrzVpPlTktez/EK3Ben60sAyFMQVv1kqycwXN/hu+00
ARVPpmLVp6+3zXLJMHcHTU8YyKNR7+PEcbQ+7xH1fqCeUOIOO+Yw4duQAKo1bZyj6Un9KcJEaEjC
kmI7/50qLGV4nZ2XG7zsrjRw8J907YeU2g+BkkHbEmtL23zpLHVRQBqcdIMJGdIrwq9+KUjAHatf
BwJEAUYt0Nudo2j1MePPhQmfXFUDuNqrfIUGs3uvMVxlymd2y6gmCXPXrvd3wHVPaRQLLQCQyRbj
5knlVf3arT4x+IMcH9FS8G71V0QhAs1O2Ox5Vqp9Q2Sg1EsaKP8yKKkitHSjNk0ANN0ge0GhBWHb
O4geB942ETePJ1cuyI/nffnTucmFrmlqj0Vxwe1YY1v2b3WX8yGozeQr8tgMu5/1uvgKsvWWTlXF
RqQSpXYlkrMv1ZJY1xIlDPLLcASPTq+L+NcqWFeSe6EmvQO2gNtN8lVd5TkDmZ0UqAlbh6tV6oXh
tpPYyklDy/p+5gi2KvnIiRIrXPBYiCQRjx13weKx97ibag8MLxC6zqLv8oaxlGMzGAaD1UlgiO+7
bQ45vafIqbABHljvNdKeUus/Xhue/4m8HJ4Yfn5KfTuSJ8gMPHixTsEasanL+fhn35OHD/HhPE0S
0d6UkuFDpN3VVBsxzcZZMy0AcyNP+1lUUgTPKd7oF2R6Rq5mZ7In1cVHuXvDKtCBUukWgUEYOCzW
BY7vxjD7jm2UkK8nG3PeWtkP5qXp29Vv2ogeSR+EL0OPSCJxVaFpgGiLt3ZnlnepoUY8cgkXl+c0
cloOvdrFFyQiO97vTLjgTV+GmsQPKGrDDorY6Yehoze/ENzjL7qpkId2SbUc4PFwVzDxIqkLJtzU
YXLuONZWHiu7HJKqYJrevCltDRrF2NIsL0e7pXzJOnPp3zzEMx/BB39BEMn4Gx+H9LCxMq1ngzhr
jebeWwwl4/+QV/2+govi4ikQmsb+Mqt+B088whBOc8Ou5L9sng5XkBWEpMLBDvoWIC4YDL062hii
W9qF7j5R/7cBdFLRt6oxUOFszX+qDklN3sUbeO0Ipqgdl8UszrFHcM2O7LrhyOE53QqnTkadO3d4
hLNWBaMIzOQB5bn3VX1w6pCamSdbV4mvR2yqZYE0rzOI0NJ27lCej+r/hXBdRnXV2E7TcAtgOD2c
5bq1GhrdLXkRS5eAymKHv7GNhnELE1DIPd8QS6Th4d2GFgjGFtaaSUJIdtHth8sFXtYuAfucqpv+
7yO2qqbkmZ91rd/ZehOjzB4/zSKB0fHClsb9/uPMinJa+ZFeTWF5UDO6zZJcAQkArpuwBGdsmEln
v+tNyhzRTMGSV0i8eh1/pqZ9C5XwXAESlzX+NEIKAW5LEHGkWX7B5BpSR83CpGirUf92gcCJ4mWJ
WTwJECFcgOieek4WQV32dH70DHIL1S40yrbCqfHZ2Gbtks6Ocprf0pErfoyVGVI87tzcNF5Ddvqm
R/UJnA+00Z+FI6VoGMR3W95mPg6CE2ZxTrnDjWTumEZalbEL94AYop7PfPtUnnTpr5f4JaMcHLHl
BbX86vewHTm7cjXK2Dd+au8tA9c1IviF5m99OnP7kC66PtbXXWVtJM4mxvICZ7AiS3jkf2HoYRZt
3jYnbqVDAiYZGk84eaIUHi1D2VSGJUrrk13XTFV1NQCX+7eXVcb3JfDTU8c8xubr/bqL3XAodqA1
YWPkYYPpCHf+CTttVpbcSRJHzdTMMQSUXH+n9tyEptnMGVH4c4HAUqVoGNqeSD3XKJDud/U3+OLu
yuwx5lUc/xtkSOnqjCMfx6XZr0J8HBa7rR1Rn78VHm+Vwyg2Jazylm6elPrqFix1msyr4uosBDzY
Hin8tisP67GAVl5507MurJzCMaL7NXCvFkfMxw5DdOiKtszZ4pB6PUtpadTcwK532niYa0TzmJ9e
x62fxwXgIfSqiyAgJSZNaAEOgEyWoVS5nB3XeGr/30gUzhB/qpNF+XDb7C+vnDQGRjUEpUMN4YU5
Xk/KqA5l6CjB7W3uQ40wPUqFZQo1xHG+7SMtpN9HEFgVNWZzEP27gB+KYXYMgSrSUQDZ4/BDez7f
jLq4sKv+Hf2gZhF7TwonVq7/BZKB2G3FcG+0BiCf9DaLRCprbiPC2jfgG0zvtP+lTLiXvNPRwh7h
mken0SSlRDUdW94O2O21WPBKbwF2nYgkp2A0D10dKsxvTd/q3kWiK5J7eJb+WWQwWV9EQTi4h6Vi
znL2sLgdt7Io6sDUE/k+nyKJ0m2CVRxaEKRvMdVkX6WOmhrd1xkI5Qu/ekqHMlui/E9dg00zxNGS
xNxea0nX97iEDuaxNXBlo6D//jDd/FGwpWoCMy/kX2dKd9b2cLJL8y9nfTBJu+bt55e83fSRQmYC
HnFTHBygpAqgnc88As/YpVtCSplwHESBaqGNN0fk9YtoiVOShksaHZjNBZxiJofwmkhjMz3x6SJE
yxTtZW94RnnfoRmBwxH/cdBcGrqhFNYF2quOWnFn2xE+290Im3pB/2cUkDQDS6V6pvN18l2v5pH0
yV0z/2DzlAGOZGW2/fIvdKjP+UZicz8gnuxi+Dibi1ob3IluQst0AedN4c0+8sSHPB3s/eHAjAeT
6cV64hbZR04sOJ0KmSwcggvj1+AS+BlgQEr9xhn1A2dEjaYgT7ozZ8Dfh+UziPkaPtldJijbLs/m
xkNDrFVlAWNDRABeh++LeB5+a6RRYdsFhORsb8ZAivYaCX5sIKL3wGAxRX5/j35p9i9nEjC2vZ/Z
9IUdmugAA74QuBskdU1xgS8Kj60zV3pF0T5Ad2R9sFGKfQEzoL6SCZQ1+g5H0Ij0bzJGBgX1zRH+
1AKx67XtORxuw3xZal+At00lGgzA+PGmHyPbjn/Uch2vQNIUZf1FN18A3bdie6o/yEWYmbyrtmR5
J0p7jpVOt4/SPKrPzNdEtOovsgX8c5sJz/u15a3/EFt3Uilm1+3VUdSuiE7WI8hPzM3pTthrDsAS
+DLML04iz/rUHYrDFEJ/1VQcf8C1fRistJgeZ5Di+1CvHHw+M9Kq5apn45ZKEvvn0PcPLg0oP/1u
M+VnRg7sj773SEuwn4lHluB4Svx91A3Rjsyg6bGpn1qDm14LOtJurc9Of2cV5Wj4lcO/JRO68QgJ
VP5fOrOPHcKmyUc7E5pOdLLW7Hm7/i8CpH1WQ/6zJbITRV7bIS5H46Z5MxPBH7w2IzZSlf090jC6
vAcLWlpTr9DwQAPS903qN+xMmjnle0oN0COEULJn1yIr4fLOfBjTFjFhog/y+Mn6EmfOxUhgH3OW
QwHWkD4HxchOWjEr/tsHRvnxXwqBlnmWk4qSQlqt3ZFs0D5f5scyFDTi0wJtfeBSbJ4YBN9iyYZ6
bOwRs3DKFhQwv2KkSGgi+xLrTvkHCzUGiFf6xpaQZsRfh28CYK10TPqcyJ/1jTCvbC0+Jx7CJuyc
ubJzchQeFf/VBpjUZYQvHhHHYS1EgfGyO23j1fOJDryc9wJSl52cvcUG4ufWv1s9+uVnh2ci5nQ5
CNhomW5yhA6BM6PCRNJFcbqQQqeZe8st5UgikrjhDt5MZk5e7wTEIs+wpQqI456zAE67ud7NAftg
7MaiVHmr0oVCYS2OWGKsAOtteX6ljD18fJ1CScn/repvuNU4Ft2p/cav5nHvz35AZ/8bY4pMc027
aC7z5nltsXdO8Qz0GcNbQKdVWZtucz0f6TBvtYiUq0qle/z48SQC9YtZc0nFfV34MAgBWwCg7LCR
zGChVL6q8eGQFppK38Wf/lrpI5dB+5QGK3vKxIomUnbzlyCgfRr49jkQakP5WDA2JJQjMJLap7K6
ciHNAvMjpbaV0yCWpc9JX1i+M7PQCmNzJ2vCfXTVUu3RHBt7NyRVckgp2dLKnc8TyQUy0F8ZWvYG
RcGz7al8MYBm+Xl0M8riXA6IzZ6cim4tMifcI2gXfzCMvfKHWeEG01J45V/7/MishFx5FZdsMS7K
YpCSjqtR55erHIf4sIVpbzwghjkFyh1J+y07B7FWOUH/JWygGLlv3FWwnX3VNcPENIqYvrCcBceZ
/eS1FLS87rIZZSM3L5FHewohyFlF8H9pANbvVDOM2jN+mHQSvXiS1PL/PaCRUhVczm6O/8nF/SdL
zJDIbddm0tIYp6LBgIOqnpe+Zbv+pnu2Xb2PG5x1/mO4iP7lxGfvJn8Huo96Koz/u5pDwR/6pmsS
nJFRphQlhQ39dRQb1CTt3TkZjZAb1RUBTe4Udv5kFX7e0HpqffwFTGqFsH87Aj/A4tqV3Oca4/FY
+yo1vKWmz+ji7KAAC8sVYmcX6rKWlMNoBu47u3SoO2+GxU5PoknpT9S/AhZb8uMat173ZqbgQO0S
YQG7jsA+wUZBbnnAe7wVuOutu90EHTydth52Y7jEVBB1DfpWpjQADzIL2ri1TGIvSIN8jkqkOnxS
gequ2hl77owWkAqhUv7PQDTjjTW8TowV9fItrANGwLEgozjfL8MKWIVxZ+yHGX672RUQdwwJEkQz
7+ba31bmLKBDCM07alHlyfs7+1nv2iCSW9F99Y7WbZSpmfEdZRXD9GOlgUR+O2B2PEAei8z9yfsQ
yAIjAKMDfeXs3yqV/ZXJLTWniNH6CaViJ9W+NltBDXPNTQ9Bjem4d4QABLbnmsIUkVE7kbJbfadk
vcUBRvHS/JDrEUMYBjgWxfDCpuc9+aVruKhO50xqKj41/kALRK/XQM14piAAbmm5T6HqRmcUkW0y
Fxmb3UCLtmqhpAd7GzBFN6k3aWxXQhoQHS/TJE6cx0cOlNKXeGoiTY1pp26cflQ1BCr0SgRi0bDY
DAKX5wzK0oiH9MmfM3nk/CiSD7dCkBbXfvcyg86xm1YzWv+DGk6Yz8UMzHgdnFthb5TE7q9qwU08
LuJ/t0m6yDKb+sfggqyLA14iKHaoUAxhuXZLJaE4bEXRLgBFnLQGy+J1xxMSCO1teTkddDBYMat1
FfyB1L8Lpr08OaaRDSqo3CJkzjxSa8K79BXRToQqvbOVPO+DK05GCRg45gHNWndz/BR+BkPNCHoI
c2n88p/sCZdfK72+Ftt2c1af/xY8HHOvDwfNIHEpSnp/0yRCzpIdtSiet4gkJhbi2oWXBOIqB5ub
DkYH6sk8t2vZHLMMvsLcjGHjjl5SZyKiLkk9AOuUdLcAezcTmUhAP7Dl2u0gvtMwz+hEO8Yf0PLq
IdzxEdSbu49jzHwqayJkRzU15EyBKSFMeO41M5gaU+sT0ljT6y+DUrA/h4FzufKwGYLDLYVtVmrQ
1lJDbXolEZq4rwoSEnM1vADKWH9MPVAyl5VqrcdKkkbW7FZjgUbJcx0E5z8cUpWobPm4bZKgtcvA
3++K88qk695+G3lMSAWbq3fB94j7pUeWSTY/VqyZWCaD1OWl8bXHoPZJIHas8O3jJGKRSTNLq31M
n8pE6RxHLD/Sy+/9GyYKAoW0m/7++gup0ilAY+XZO66RU5FvdFYgnRK9PDp+/M/2a6A2ShwSwlyu
Phawl32H4CcCauvBG7EkCa4sVEX8R+/JoadTZ4veS2KqDHg2t1qOzkmqeSbJ+cd7aIrNmdC+I6Or
RU0TOecsmqEZsPN8MvGBVQNLrZDBEJBZxovuKCcc/dXGY4P4mZaZXvDodC4rXWtu+wtjYZhBcFe5
BxxufJbPbCi16FxOosNjzb7z9jdcKiTA4+amYi94G3ETUpvFLCBe6HZpxrsjRrPPzKKPJtmaNRJu
bKu4SROB6nItR4SP3QblCQq1ddPcpPHLzRagCnDXvR1I2U7KdFareP9+kkeuqvkqTe/b4RLdPuA7
AUr5YwI1R0OSk89PdS0lU4L4pagZIVZqf/KhsxW85TyW0jl85VLHAVkFZxKLh/u+DAhxvRNMEyjo
IC5Mzit8cYKA/kWcBqOwce7RqYIrb+86m9srYgy/QKunHLVSLm2xPAihDWaPRGPSm4gGCcP3pHeR
AJ17ZiXKZqUoThIVCH9y/frhJOhiEKXFoq+RkSsDtvX17MRkJhY1fRSVYKZr6zJ7d8nt9CWBeOtX
Y2KyblaWfVDE8OamETCIRPfRcDVXa15fLacppjpiQUXcM8D3jJ2Prmv22TK888QamD1OOSJFC62U
IyAOxMUDMNZDi698Q7Ql+vUBKSEAUkYXiey9mTejbJSrt2CMwPithTuxjE93IVm3bthTDXunNhdW
OG+vlcu+qyViISY705N7zR75K9quda0EweIeZdHmxvKiYGAWK2Kmi9Hsse3x+RspHvpdt1itvd41
o5SphHEubQEJmWpCYaTcxjunZwWrv3G2LQS8DQZLkK5w4ok1aBKEGWfggUZt0b4gzhqmdoE7dR+k
CnYs28IiY70lJbsuViFPck/csKzaMIIvNs3WGd8nMHenpK0Jn5wkxKufmN257/nMj9ZqPxIhhExS
n898LilWG7yX+rdYeZ6oOb9u+DngTQ+iAQM64KbJifo9OKplKC5i2w0V1IVWozO1CBsZLoy/yN8a
zvwRMZHBQMGeE7y4GiCy1Kom/VbuYPQRgo3unIXStf2Wchxjh5bo3FXvyLtCJftrJ5vZD/Zt+qpn
iExY+6Ysp/nrGMeBjw3+rpvQSMQVddHd862IbxqL85E+5D4jB9mvqfHt7UI7drsoGeXZFLkoKkI7
GkblFcJjIX9exmeCTp/gvQvCBq254AURler9wsmUKLZVU9VRkPWTaNCyu009jO3dGpI/ux8WQmyu
t8ymfg4PIxim7P3sKSA+efA7QJN2ZDmV3AYRxsDb2mcQNlRp4ZiLiArmmO2qAF60T81q9BIw4kkH
CpJ1AKEkwnyHieuJXJjD2xxYh2UeUQZAS+sJC2ChjO2H9RX5rq7doHg3M/zD9HPuzOu6ODlCTUrj
ygXAlFGVFOJej0O793qUUiUwmv7l3L6xPw5LC6HPENEOdpYYYh3DYRSiufl0Yy8xk2pDCQsGuFEf
ADlo5Qs7+c7aGiTLAzMue+xY/vwTqAwk6amhr5vCDVeNU4goHJMCks+abMXcUbuNANntO4D/A5VN
BJrAkw0tNkE024vPazdzesodNmM8TRbeBDeja/Q39YJMHoemdGIF2t5DuuyjJgjlWQ1FZ3NI+bjH
5Yv84Df8FHvckE5FlPzvw58B/NkkdBUi2fx/kDH3+QL2ZEFRp+PY+Hf39O+qProcz3hrM+IJcZ/5
ZC7KdT4mK5b5qjVtXi7YZH8mR9NqlMXTi6AqGeHrew+PN5V4Zvh61XkNKWFAlscWNwZrBYN4SRMy
pwhAdMabBOnhy9NmdYMawmzhWVBOlimo3on/JhZRVa/M1JuyxYaOFC08GHpF5gYtBcd2U2/67mbA
V7RgGrJXR3YX321w0tLaTwQJyFXMemtRw2Pm0SQPq7tC5H0qlruRwTu9HHLRRNcpeqWlDbbLg/1j
Hf2V115eeHYeGivHBzyPabGCM6k0olPje5yxafgGkAYW7ghddZpnjH81xAjOyR/2FPe/+Sn+3+OH
/EjRtH+RkALgtGW3h760NFrfEg4F8TdzfggtR3iSr6emFQASgR9t7r4argsxV/02H/Ot+RpwONr6
KeKAVNbPSVF4CDzwXFSmPVwBiQwGMihoJIrY9iAvqak1NzU84627BK2N0uuhnJeVsGJs1pyYq+6y
mJmXCBAUxud5ULKaL5heBZyJ11U/pu81UJFWNf6/G1SAPu/uPUVeAfzBw16kmrNM3dZhpNH7o7sI
oRwjQ+VE45ZrW5kIaObDJfYkRkGAQN8iHU8d1x4NEsdxm5KUCNpIYQ6RdPd4d4T30sHFm1STAj3I
S45BX0kjX2RmKBQp4bohqwHHb/u45sTywnGMETvA1S2pdaM0o2yavP0Zn6X3BhWIHBd1/CmPyvLh
b1gDFAie7QVmqR0tvoyesJUPHrVypKsxYghloh6nKg0YffSyZCelGSkd2/hG8Gne0TXkLx5FHVgb
mKXxWejahlhgyiw+P1o+WFifKVHrSj/51oxUy3Lp4pgA7+lw0oupg6FmwmG94yC8EAL4r1aog0CM
60hInidb1zM/LChIV+LFvsaXeGnXq15ZQw4hTWQBa7YvKHl9LIbzdEs3wYP/aw5rFhg8oZag8CEv
3nAKwiwYVtcOBtJ+BuXFRBlbImJWNaE934lRjZz6tDlcR8Y+Frb81ZkB6vDiXRxpZe83IpZf73uP
lYc7ABsbWe6+HtdOVF4kY/VNzxIiDNUnbMMJ2YjetyBoHMubqkc0GuAXwjJbxlHyqbgIk3mKnDkv
xQIS8IBYssBfy4jmPgAvS9ArNAp+6OsvKIVuG21Fqq1xTdi7LJ0boEAZDYgfRVo9hHRWixUaaW83
vhMkvGD3KarZSxoMFokv8lvLjJ8h9dGNGOgSMLymR8gdlW016Rjw+fJlCmlZSuRdKt1cLlh5M4Xv
i+vKSM/wnfM4YYq3UAPKNXRDoeg9ppaZW4TL/3is3t7/N+QDVBVY4kxHR1bouo5KKsTDYejyAzBM
qdeMYFLeaTitRaIZ336GDeBXGOEdDJKhthXMAg50k/k9lVzKxYkxM43D/GQOWX3Y/jCwCbOGzKov
orGox8tWBIamfzUMJ1/rLG0U1HuKEgNWUiaQnEV7g2MENeCapUE29jzbhVAgYbgsIUpdRyt9tsaS
hqKj9A3pHYXJIAYgiEQwGqBP2X67IFxGmT6wBE/LsH4c2MShSxngnxG1fVgnOWuFdXgLMhG83d+B
r0wFgJkLoX0Uah2vPNFnpLqYJ5fZhalv/inRZpt2J7wbQiS7+eyoyudcXcgR5zInxTpFHW8cLLmr
z9a8HmX8WeLvvcdkPGpimYbZ3kgPfuJGJiuyF0W+AxMPUJ3EGYBt7B4TEssgoikjT63ReNEM7VK2
pSSUJIjKkKW9bd4p//WKo15ypOsFkEmVKc/0G/92MVK+k/TQdW8uqDdy37iiNwOYdIPeaStWyGEg
Ph5aXbtCpdBFjLAbaKzqiyeWxe+mEWq2iA7RXLDAvuwFQhmvhbBC2T3q6+SowfbSQYFL06DJH8sC
PSuvGdRORTkkSdz9+ScOYAineIm6Dgo7mP/BS88uergINVCyhbaYV9lq46Qd3/kX4YHetf+3Qngw
b25pwWFpwYqOBtneLSS1oL9IzZE71uNQYW3blEKZd25IdLg31AKPfur8WKU0EZP7RNizQWypueOe
sXTnEAZPBX8QsLQ5rToz7V/0IUFCe7lOhtAeT/mvQQTW8MvWlkvKbEW+/fx6Jq6v8HSIVKXtvBEW
bll2BjSErmpv55EfVYryZUPZFeEtbPj9U78Xkt88+MgFIkn83sx6EKCuvIzKzZ6Nm0qSuWzpIKNj
QMKYUWRkD8ewKZkopbAb7ggOLnY1dm++KhgoH3KGaNMW0sOF9cHgCAtI1CJMSD+VHf/wJ7N5HASL
EwitiyK7qQMKKwuHiUaS21OIumSxFKznX6asjMsq7+D6e1eeW3A4TTOkwxYg4cndRsHuYoQJoPHu
gbVTb4k5QKzgmDD+PbgeZTD+BsU9S48seQp9TMUmCf+ebwlnlkvyxTlBih8uiOHWglMikSYt3RHU
tJb21+0ugmVeT7AI1JhnOSPb7WFBnaaMQue7nW6N0BH3V2FF7fnY95A8Ucb3IZDCD2dtZTtWeiEj
RJhex6UkxjQuIrlmDkc5FmmwdOpzsMBQrnjo+B7w6z04nbaemlFSMxn/CdcNIIW4SLzdoG+cmpOH
EU7Ju4k14VTlOTCYCP7apQ6/HPdgH35/ZB+lTOdQSYqgJmXrCMXu9PvNMrmS5ffw+I+8Mk0436Qk
E05ZzpgRC3QeWkXz8eDPRziLLlthWmlWvMKJEsRybEl9TutOYtNkcXx3Zdev3Zr5Nn8BRJSXuZbR
n0STMBmpEOpu4Ocsq6knXVD1EouZ51NX0ERWBnf/8Ha/nRcT+endIokLXWZ6zDkDcqMKprnzFfHm
E6WBBsp+XfWBta+xxPURxgIQSr3e1ioEC0rl4+8bgryTWksIDDRmw1LH22HK7W5YVH+cKdyTkp6t
dHrcLDO52bOoRyUlYGjy+IXR705ae+HRdUE7MFblv3Sze3EHoOwxNUZX4AlvH0JAbhN3mCrSJ59a
+bo1FmmMtnehLJXg3rVJw7k5Os4UCfW1Pz75XzhMjMj8aYSzys3owP9A+0ANINXq1agsPlvKzget
GflzzNNUlIfidJyf3/x7fFV7Jti8IIdB53u27v74DT6ugrJVRrMEXCHsdPDShzfIWXgZ/ZB/oohC
FZ7Do8LwVfjbFRL9zLpYSEbLJa5H3XlJLI3la8ExDcTYz2fjYIvO/S2IoUnUTXeAd1PmzLAZkt0H
6EGOX2a8p5o2JolUy9b3tB3puGsjAEGlo59EUXPiO98vfwxhq32wO4b35I9bM8ILR5Qh98TqeeAk
Gn8vQvkYp+R3HzU8ghtVkjfz6wUsRcYrBkSBkXyEFs3liF3HEoRBCu9RdGOGWTPjtBRd1zkIQn6W
RfeEqYgbtLAk5JgYgeGyXi6pCpG7vqwI1vPgbEv5QgGvDt4jhCTvb0W35YnE5mbLyzTd4jqlfTcs
HrfpEA2fGxK2MUtAE0VUk9fM9EcoxfrVFL/W49djb0IqGtSbOZKGre3hY1NeoVTC1eI74lI3PsQZ
5nH0jL2llKhjhg1fIuyNGkHhiKrGE8fPPr4C491h/qxx6lCMGk+1/wua23Z99VIVLCakn3erVvMn
QjEMHIYFUEHiYdnfFxD5CDghohT16WdhBGEfefMkgbzesm/ZsT7tZ+HPoeWRavdyYtV4pSKXXPuU
j30Ra+/umUpZ4EzZllGPpJ2CpssOtQJD3iEZZaWzZi6zbC59W4lwfM8g8wJKQqJZaNihXruIGof9
9X5BeMMyWPTpX+8t8/z4iIzg4buZCi+d9DkSwyJdO6HPuO2EC68lHPrsGDPCXQ6SSz+dYT1C7svd
ERoQsrW+Bc5Wf3cUP/nXJDYhuy1qEqxRONxnwcl+w4cg93YU2UjIp8WOA3Jkal+Q+Hl+LX5oaSp9
VeOB0FAsr+1eo47S/e1I6dEAz1z4I8BSXjEgErxRtFe/Q1FhNlLXoTqU28BhO2oA55Vxv/euSmo2
MF2qlZpWC0n8Li212m5Mo0fk8R1Wi7rSSGS7HOR6jQjvnV9B9yrxguF6QRjfguBdNmY15Jk3MTvs
RaRnK0wmZCMhuneOz4gqq1JrDmZ6kqxeO/mPmxKo5SzgfJmE3wRBMs07BUb0V/noE8rH9vPUtTvo
LoIQ9E98WrimbpuILW1YdQBnWEObdEGzVMR570qjaXP/eZQwr2lFGaFWI27wrGUnE3NxlEqo3VkO
3gyhdssApXGsncSII1z3nK97VyvRDY1LbRSNw80xpofNhB23Iu5RRpStTI72Ef7EhX8LDjcr15BC
LNty05ZacAkAGPgDhVNPTp0qErNFF9ri8lDPF/WJjWg5jYmd3PcIoIOwqKuJH8aMh3zd6qQICiHc
cLg5E6u5HrMXYRPXJH1rmu6hL593wVSfPSmXF+5xiL92MabSRKjZDz+XoWcRdLCXimCAHhl3jqNf
8PRqox5K78bD8lir1y5P/x6jsPD5zNz8rKMwDk4QWl4pQX4XZFmEnoYyyymSHC/QKwhruZJN5hIX
WumKYDmGWntuvOYole2Bdr2y2nUYX8XPX+wTfxwdZp6reTg52lS+OwDpnNOQPMIpuZOCzuRD4pgF
EaQEKFbIGFDZiSHzG9mkwjegz5Lg9x8ZZFya65zdlgogYXpcrt1u9RVszPMjsyH5VjB9qBOAfNdL
4g40M/jXoEQDVvggOrZP6h/w59BU7HrUovVc6H2JUcSV5rG+E76exF4UT9OZi4y4Y4qfoLeqT7Rh
mq3h+5lHrVXnklS78A4lplqaOy7fdzQsFKvCF686xPOQNeaLSE5CHzHMCSb7fG2o37+/+5Nfxn/X
2rdMNgJvXWr/VfhOgN0T95JkGjx30uy2WvAG9lFfp4dFcygbysHfrGPzLH5lAF8LkBlJ5pu0qvIH
WkQVL2Re5BT2ls0saMx02LBou7LoSdeJ093E9GQfWPFpui8f3vVo/nsWKAyVMYAKd7ra85o2tlsi
+yet8NhZiyf8//OILPYBK4y+aDvh7UP0oVYVtwk6at/O2oOVoS7zn25MoWPmebziWMQv3V1Pzmgr
9d7EiiHSXDMExvnPlXKrNsegvwJhxppRYZqM+m60cON93V8ioACZONMYtCqm4Xa3cYf/r+g6zV1a
U0fZXCYHPsJYBFQCmvJdzU1Hshi9xVIdoSrqqBe3uxE00fMgCULW6Hjy4IAx//7Hjv0eh8pON1KH
oLOU6OhhSnjD+WBX3DMeimRDj08nr/WDJ+Vg4Q/g5kUvML3BiGX1bDXnBe0sA/7Wx9l+0XkzO0bL
hH+CF2OssHo85UxeOwa1DDn+lNbXVFR8BO70hy6S61oIQd/UL1mBR3LZowaU53O4jhAXtp1X0kNk
ZgQBn8RmoxMwM/xtZ5amrpvP89k/grsM5fq1ItoX5Ypee9k6pTFrUeiGQvc+rkrUzp+ujx+q7+cm
yJwsyhnxMTNFx7ZHVnFM0bQHacGYagUmiVWsg9AadbmqE8ZC5v5EIOfac5lWLCc5jLytTsCj8/t+
clbYCOubeQ7ipII9OPc5T58ko5+tMNidFy/02dCqwinZJHHiCdJCW2/d0GuyhylfCEgQxQhWH0cF
3TOf4elhHdUllooslzYcdbIWLHK89sLC/clZ5RCq6N9h4V7nriIyv5JlUMgMpLZRd80LBgndVf+G
fA25M2mrFbsGkBzOeHY0IbNM1vzt2uMjbcn/KQXIhiMlTlVi3Vj0sr18y6bOolJux8iz66OwpCI5
jHiKpk6pJiYYjIC8TllQAoyWnOqB+VajQiETAIJUbx18J097KRTZjdA4cGlRXcXEUibrF8J3Ah3b
UroUplXWbJ5EgGUMaqikdwrj1LxJe0lovZEwuE/0V6CVYpl5SGCsHhuzMeUgPDhlVu8voT18rcLX
I8+NCT8zUDisJOf78Bg8SGosuq4OAqbZtRER9FwOh4Lr8YfWPaaS4pcJXLjEqZ/ZY+EMPXqOCdIU
+dG/nIQN8yXcnxWCwwstLQldTT//f/N4QRXUCGV2b8ICnnN1Gf5CD1kiCoCef204NGVbgkIaOkJ5
1LzN2X7TVh0ltFa/e52Wlb3DcKadS39mnsJ/PGs3alFmXCekjjrqBwGtbSJ6MGzfFk/idDM36w1u
4+GUlBMSUFRIQXZL75CHuDyNOlHxtWs7jbIsZ7OuT5Pm55LiHfzPjgZumctNsQ4d/mWo8xVshASQ
uVfRRo7NplUnasK/aWpft/EclDKSzxpN0ijj+d7j7J+qKu1Cm/KL+qnU1E9Td+D35/+iY6W9+7My
Se0fADWB8Ju9j88AJoKZ8q5gIAv0C6e+ib9B6fdszmBIHKtTxmF2AxJdUaOC5VQ8uVMusz0whbN1
PKWVxBDQ9Jc67vjdr1GMY85aaiat2jUREpcMhOwb2DaA6kkgKsoLUZGxQONE4a5NNg8f6JS90Bq1
yw44zHWCecNsIgq/XMWU0M8Gu2Mz1E4YYBERNZrMFhFQPBrzcmlRR1PEdPY7tyJszJc+c95YNQVG
SnOTP60jRg6naSIT2jc6u468uAKJHkzP1VduWzwi+ICq0SYlrCKki7B+XPdM59czsfdq2JwYONQo
CjkxejNBCE7u/yNzJUbHcedly3sTdA06LjuZBsWcVNi8rDDg2hNYekmd18VB9ORtVr4ncxXjkw1u
BHAQEpshUbx5ysPNk3Xe5WR3/tCvBbnUeurCUuEecWGVStr7zlfPlrW7d8J9uNrWwpDJBl8bBiej
/0TuowOGKML9yHEL+1JKfmOfMzu0FlEodT+Vav+DM2f0QegQhOUGRxKV2Xate6FXYbrDh9eLeHu3
4BlG3xGU7jcvXhGCZ53Qzl65r9zZl0XAnJo0MMHs2ycih+Drrjuq0ok5zz+SnZ0Md3d9G2Tm7oXu
qq0loRyTE5/McnKk0L6iSjeSpd4L+uuyt0m667jUcFQoziBL73GSXs91KMfS2oMfqpU83tRp8Nnk
W9wnnshNjBUxGcTFtBW7SiuWz9EVaGqNgYDJdb1qZzo1qof5BDB7AfPTSm4hHdJ+6Ko04X9IaoN8
aotOjEE0I/4w8V56UVGhJ7KHEELvVEpzju98W0Xl2UfrG/Capl+GMY7b91VlciIQEXjEYOJbaun6
7P9YEeePK9rFbqewy/c+wCocQDTw2dftJhsprlAzVhFvZZkqgZQZ9yI533woIMJtFg8WX3C/np57
zscHRXp7JGLVVvx2uCG53x/quMbLrz+mF068S66mo2yiQp2ju2K1EX9ot2CzS/hjGQuGy13jf5ie
Hb1M2Ghs6OxNUbKlyi59Inlmf/sDF/XQ8wKRzzIsqf40+X9HsD08gj8Bgi1bBn3IgFybkBbCiM/i
yoiJ7fb2RHG7JiX6VK3vaRFwKkX/wJ1KKl8AHD3zg2xfhQvEX3qV8OcliScxkLxz9/4RKCta5Zih
DAAwas3c9wG4DPFVIcsFh2nCJjEkvo6yrE1CmmoXCkhM8c5p4dgLbgTSM/SZgQuVteT+0pSlot4b
+scQ9pWyri7qJKY5osdxwruX0EHbsZDCNrQbUqdKccwA5Fy46v/rfYFPJhh5VIl8Z0MWdqhD0CYN
+Fnn7WjmwpLQfeg+2RROUPgu9vq3TsLoBWXb8VcqdpJ42UQG2vOj+efgagmgFMJ19bM3fOZ9wenn
4wOfXPl5puxy5la5FaK0OJRhRuSsTPpMa5U4KzfsQ6UbBRUkpcSGlQ1GV/Xk/NTE4KWwfL1zX1za
bo0t0cyCtyTr51PRXyXIfayaoGTy9vpIhUYGocdIrg5cUUmQ1jWu4NfMXxVbWS31MAF2rf85by9S
+JGebPC6CWjXwV69LXInRk3P73KSFWE7NWkis6kIjKri7Vs2QrlqWNdOXb6KCxSezaESNEYJumDh
7p+qrgDGkbuUPjRU83o0FpQ5RyH9RJhXF9KUPQPjXcoXZtSTxQbkWboVdORAyy1ghc8x9Dnoxohd
vOwhqrL1Icf7fsihVzaXyrhFk+jXbErqnUVe04zKFey6rm8UZXFDpGgr5qwcYGxd3TAq3x5Wzx8z
4KYWrdVqehHnNobEoBFaBDnViapTwpHtKPqD++2ENLr/1QoWeWb87yIYmpK8cMBrDZnG8wanN5fW
vrlPRWG+ExZB+iocfWDHRJo7y/gfAFdpRmng529rmcgB5a/RVXmYafzqCW+FZkr5D8cg/CpMdH1J
U8JDXwT5YKZoWOXhANz32TXYTDK2sAa6MrC8gEBnsHffrkGcjUTGtEgkGdp/rq3jL7P4UYmeXcnI
v0ihN2P/VwY84Gegw8byhYKIEwaLtAS/JCStRRvN0eCymHbKzV6qxZGxOyGQG1nTaArljYbxYYy8
Wmhq7KPxFcgfC4XMRt+kIhxl0RbtOOzJG1405ePr+IdLdTuqfPRu62UjcQkbwFXHPsCPu0mFg6v1
VUgqMCGiaCL1v5LuwzGrpktUlOtMo81vuCRAudZ00AjFhx44HfAqjGmjQq2o5KJP2UrGaQoLMXi0
K5DPNNQ2x9RPqpURI7a2KIbSjqIbl9lRujejbo4tTWWWuIMQCjOAjb/hM974i5VZEFqtGicFR4iU
DuVATpLmAzU+k0i42fENKoDe4qepq726+D6zX4aMH9WhnQev/DFmzaKOxsm+Et1ss2aqmhqIow+B
GON1A6SwIp/0k4/HE57Dbbu2+TIfmOe11s5D/LPTWe2LyehIqhTKdUgQ3ywUOpo4OGG1OwQHOzS2
9U8D+GcPH2Cb2/iQkqkgQXXrRC/LpdwuKGbN5kmY99M56Cb4kZblM+j7BqX2YmqoL91+Wf/JG091
MG7t0VjjnR8Vtmj+y7/YjcNh6ACjyNDIzMfgiJ5QZYw0UqcY1dFaVwoioj0s9Bg/sA3MLvCuoYy+
ClLeH2yiVE7WyMKllE+oql9gClgupeKTydicZVFPZzvDLsTPgOR8ba91xnub+wzpPA4L9xzSzfXc
Gm47WIWrCtbkHMlEmXo24cyhcZzS63qZJgpLGqjQiw00P5y7VyH7v1Q1Y3TZvURs1hw8oV3TsJUE
LW7v2ZoD1OcoRunyjzC3gXEX+N3RkwTBPTv6LoWg5pmo9qKMexyr4+2fF/RdKClHOEeycEDp79rm
L8Tu4T4AhRjwvasPcOM4FWLhOjcXyNkU1nYtRsdovKPOeCw2PxphRODcd+WmRswG4BGPRmsmhpnM
+VefzE6i0+IQfyqhJ94nWpdhSgNQce7u0nV6jbS7a8aqmc4XBo87jjBA5eAiccWz6RXN1i4EG11G
zgc7B/XXAHjCOoe1u243tdbrSKp16hEu4uxQMkpyo/sdW2Z9OnwYJbu8lSzTvt84omMqnpeWd1Mr
s7SGvOOtjA1K7uQgMeyj4q6x1d9rXFtWp6VSyAXqmbFbZTawhxSgy49k/LsisDAafD+IDE9qmzIr
ZIS9FytiUwIgsDx/W2n+3R8b0Rbg0D6n+8JG4Jgl8qGg3Bbv4bLXO1YDsUqvsMXU0s8kJG6UeEJJ
sil5nyED5rIMzjnhLzBmO05PFTeoAFEvXwrhXNM+p0Ya/866jK6PWKhQq+YEFVbO0N8o22xW/IR4
UQfiTRbaf7iP3AHHXwBs+r8djQDhszACynS1A99HhxlsJe2AcjJRXYZhf/xqxdCI4Dbh+8lCjoRk
FeldtcScCy9rCF4q0fDkcL8uHzOqQKklRUgFderFiiRdCaSPKHTPmzYd6r7OppXg8wlt3UNYo36b
MAwZVEg/Bnj4lRJUVOPBb8vHMqt2vAgqEGhVk2uaJsFJRpQyxuFuPKxVlk80hGDvpn/llskdc4hk
e97xsuildeDCAPzBtkd7fQpf6+UlSxo252MiWEtR2qw7J0giOP89yuFkQsLBmTGVvx1worgHH92m
ApISoOFZV7+DtDutuDbpjMCK8WgLzA/1n2CeWXcQyia2GzbFqaLf9OUy9j3GbB/Ql7U5KZ2sNm2a
ObJNx50xL/oyA/aPKlFU9dlPQ9qjGS/Ck1dh0SNZ8IJbJ0sVvqjUzISf4PUKZn6Ij1UwL3LI6diL
Z0SDIbH/sv7jzYIZ6kcco9Qdn1eqeakEnH9h3AlK/9V+khxLqfbIOfv3XRYlNCMpSHIehfZNeilO
9TvoS30n0WX/CAOvl9AmhrMGtS9YYkutp/3fjh4H5TGZqiq/CJx3z4Hkzd3lhTSrHbGsY1wCVWdZ
DCk+8PhEZB08kK1MbDGtCVE3hEzJg4zj4oEyIU/KY86Wwu9iApwKHzq5SoFetsc1O7Im7HX1ggX6
z2NNoNOfLWXQbcoJO5m/oGcCpXsYr5LZn2V8Auu+3d5P03uHTjTqqtIB5q4sTBkwvI09qgOx1+u7
gPgHg0rJJNtN00doP3MGcMhH96kIuQNWvUQsE2+eQvQF6ZyYq73DfLxYX3eNbPY9QucGO9FimQnt
e52ZhZvZquL3uZVorc+ObfF3X6YhL++5pYbix80qnpgLbtIJxBszONfLMgqKTdXJF4/Z+CcT5/Ph
anxqq/cOjbl+qsv4SxrsTl0g8HEKXmASuCfu1et6Tbx/gq3P5GIpAHONVHnb99qA6Ix3W8rYYiXa
QAR/gP3fcuQDpE+UxSJdsX96cOGlF+gUm6KisI7brZuy9lk1aCx8l0/DrM9Z/vLaP/Zsb/qFrauI
aV6elKSCJ5S/ZWl+VqrhMKNz0+4+CuQUN8x6WKDItPNjSQoW8NXviz4Tv2ag/FIVI4db2a1imT4J
yes1muNVWmCfEI9ipxd/JwQbtQtjEe9em9+UU0CuHHh9BLv2oSqLlfQA6mmRjhbww8UO+i6uKgU9
475d9WAWP6uuztae4EN6Ef4YPNz/sfLrLTYn0QoINoG6/jSwfvQKJBxIzN5cPUd77APnYpqSN92x
M9IA2+TAZA4YAZcLp6aUeHWIlKba7i6lRQEFgWSKQCphdsENsDlJoPHp8BK3U0zCCyQWD/ISic8E
nbT+KgmOoExyu0sylc9t63UDSI+i9yEOMLESHzaxHAnRSahcj+HSP2RTzwpj7eST0u7dvtzYahHn
5y27LbTKdHMqRmfBBdm299Qu6zQPitir01qRkU0DJ17Dkhr8c2YfSvmihYALY+EAQlArLwa4Uo4V
J7jRpB2NCsQ3wIwJ44aAII6iV8kwi7KGGrUKIHo2B7h6ZMOhqeNZKNBgdq4tD+aXRG9EbzA+9vcB
YpCpyoOl60cDYKDc6E99ApSsnokA9hNfsoh7x3E8G6AG/l4qLMIdQNCnhVskjDufp4MyxmSiy0IK
0s6FSqFsIj7KXIxM/c6wkAdxHBYejIGO1BvZtIjksNyQ6c34t+9uj9lzqEt0v9asj/ajWL5b2ylz
hnRSPVUgpq6i5wFSIVYoRk3HAZtlLIpA0aILpYv91tztMbx+FLTCBmEGlq+EhUMom8LGfLqZvLPG
Nfn66f+LN9IV7nGfcGGmlcRh8Vo7lhfripFf4n1FRzG/nngrClQnv/14R/17d2vq9LgLcL5jbTmo
kk/LDFNHQ58WKnCeJlU419F2jrObJohG4vra24kqzdorxK50/jh0dBHc2E3iL7yFAdS0H1bGgex+
m94zHQz/o+Rhj+LUCN+wR12E7H5bJMzwbCK2Z3dVCS7bRwQE6vf45rtWlZ9NgGJhvlmQUkSB5Oho
pSnbmnAPygLeXWMTfStbXA+IYzVFjbRMB3PN59qymy049TZKFXEXux2t5pQ/SYQhazrPwvSgG82S
TN8PJocBNy6kkeD4r/DlBXHyAo/0vEW11J9YMP7cIh2C8714kxypy2Sk8axudRUtZnsHm0MRQuRf
tihUO7koms3A1GnIjKPMc0hvvlW3Mcs1Qv08xI04AOlAW3amhF1nVL37iISP4X6RSlkRKXQIDfiN
4OWHZtKwfk4fFpSrXwBun7uE8OxwGo4PNrtIzJ4S4NravjRBsotqdUOq5jSi0PurUP1Tk6mzmAZI
MiWBRJ3e+olMkYfi2JvFAUMEtw9MFpcuby9oRbi3CwEJcGpruCMG5p+CME5Yo7XkzD44u/vb6rt4
hnYOubBkTams3Ldyx7S7+Jc9Z68W1cRdEEc4qh/abKMyzEB4KoO3L847BdhFI7y8p3HU72ANql8w
j81j9kerFKzDYhPG3/mgW9OCH7ONOIlvHJyNUEl/nO+t/MOYMwU9ExioeYHyuw13NSe5QcYSv7bN
or3rcE+S9b6SCMEAVJ1osl6bwobE7OO1K4PjslW+8p45tTRhw+VRtaLdslX1UzYiHC8VTlPfEP3L
ioWP1+nosLjy/Y7mMfCr1ZM4kQHmtllD+00JFEnF0oPTyurT8PTh6aN0dHrrrIjr16dA1r3VOM6B
brWllHzCycybpg7zbAewWg3JEiK3bJp/u66wz3Juojq3V0Cw8oHjTJqXZyrsRu+ZN/AbinVwjMmR
nzobVyn9+sFdctBbjQ4BKrmAr9siZZFSTAPd9TIlWRb6y8yRge1cVxXZOatlksxV+ceXVrm3WZaM
/oPTJSun2uQJVnIK9Ri2CnAnimAmOSq8opbGseE+7qENwcrkkniE5GPiHRhnoDZh3dSY8kAHfF3R
D8yEbgpSWQEOj8e7MoTAJjIl31B3saNRaLsQCFgUhtuFPT7ng/edhNSQMpJHwuwUQp0nbF8mZ85c
6xUqawLuKoIR1YZ9kej4WWk0sX4Qkgig8Efb+/E6QnoUBkxAsIBCR9Q+RF7fc6PqlXn9Dd5OgsY7
kLKHspyF4GfEHd/XaqdzS5lBUMeBM10GH+L5r8Y2QzC3LNhhh9XwhgQlmkhOEoTORyuq9oiv5FyX
wZwAqgU1H7g0d+woU8oUd3Qco6FZlJkNzeuuO0+gGs3jQ4+4QfXf7neNYl1fxM4qtgPjsFZTTltg
x1Vo1xzdL3gOVnLKwRwAASXqNesNk27y/DK1JC30HrfCxgM7m4UeUx3lXy765laBWzVhBr9hK+4+
PKvx4sWg5Ur+BtM8HtboBhIg6whTP7aUnm26auKr15inHHwjLSV7tN6OTIbXxBA6u4Zla8DpnSud
x7YuQnChFUE63DrIagFWB36/JE8dQ4uxknpsgFFM2Iy3y8V6OZepOv8v0RLCn3aulKjeK5t1ix+V
e1jIJvT2WkcTNk2mV0cwY0cs7dOEy9BYbytHkGUjYtDI11iSo9/phWHfY1m5XrGrZpWibO43FMCp
ncIx0KMQXsbV/KTU/9rPZXwtm8NPaoXUQR0tDHkpEY1fOos5qpx6aAvMPsfLk17kolYtWl87WxK8
aDpEgJpJJtAA7m/1wkLrCeCCwtNHdPKJ16aQWCl0yo3/pgcMEMHzWrhwZXB1ZTpC7E1oShvP9yO6
X46GLYCTu1Dj4iah8aGu0KaYO9jjNgHZl/4tXg7cVjwLsRx2IXSOtI6OVOBYiJjoEmiXr61lHmXt
vpoStO6u5+hIQYm9Xm+uK3ncgj3LswL8uaPhIGtuqfcCqY8OMcjRD6XTKIeMlh7Ws1J1A3b4JnH3
vXaeb2kgRHjQ+RxpiI07xvdFgkbrPrvMJWkzcjvh/Oug/0pMshfO18G8mPbzTepWfPrtKVJak969
WlTut9KQ6rRlOf4X5+ww13iV85331pXOFMtM+9v7bS1AmVCM5JdSSYsylUv9w0E+A6dbc0qaS/NP
4As0d4XquGpEJnXOvjnz/Q5b8WKm54JPMh+Kk9lBHw+72YXiOO7C4OVDJ/4YxIIcIT7GRb409/aK
QOqCeMVKgSt5JTVjUvpuZ7jdUHpnDVJ2vwb7Ogh1pTRDBRzyIYLVJYMAAGFhu3le6xrBgjrPKkBU
+XVi5tiuTggAm1cSBodamSM2U37+wHB2T5QYNh9xBXy9qZy9t/vv85C4Sy5I7uIXPsxwW0u1l5GK
nKBGe9zSbiuEKzSomBd6EpH0kYtS1vQW4en7JC7NJswhGu8Q95QdqNqgrQ6sBcrh07NnBwmVkJqZ
JM6X5op4U6RKY41tHUVhEgyV4eBcbNApKFtOpMOIfd7WC3XbtBt87idkA3sOTA81m29VBZlWEzah
VvJDU/huCHZCNSYqf85oilaAuKySYPMfsFjyv/o0pI/4VfjxA4THZnva7aZDp4YQN/v0ng5AgWwj
CQThvOdscMeGMRfObMCTXAxdMugxpnzKcSBwppWNCCAXzW78W56vCS3edaQmRPt1h/QCFag5ZCqm
eRFrejCALiEfuSOGFulwByB/8Zxq5bmSEfSAB33VJrUE7pC63OMu4OsI90uEUQsWYjQYD6lC+AWo
sZbDE66fgC7c7TjIQj0DNUUj65wMMcwtzHNkc5hcd42wtyU7uvLN9fx4GN9clzjSlJ117R6w7g0y
He/59CZKJvVDYLqA/zhPLaBI2bN/KVabV0/cB+f0gLBc/3rKntlY830JUOv7uvd64TxbvPw3gnxI
00w2z0OA43lg51EsFkjf6AVS1gbpx+vvrWM/zjCgqsn0pJDw9KAgbAIDMHDiwDwnxD+9Mn6sFBf/
1YT82J0c3gGAriIWZX/30yakiJWY8Gm/WBdco9z/kAdrU4S3RWnla1x1YXJqlftM+2uERWNrY14s
EyELB7GIDuTlzA++MiqQr13Sef///I2nRgPJYV/4YsOakTb4xV+12sgtYJsABS7Nn53QYKGABDB0
Ww/mIChsfwczNgC2lD5DqhxoCfrYL+GMnqpOu/eAPzYv/JWqz6ykHlaMJL+npX41uhryiPYuFm97
P2UukH+qFhTXcV2L7SrgqB2wkdQISdqaMBEpyrKtc4XWaTVATJfNDMVE+dHI8ocqxwG4NQTrKPmn
U0Ojnc5KYmB6fwSZ+PPXKkMPCHEuVvXALyqgoGo9ice2Fd0Q1pDPatszHlXPxfnOGiJCy3x9zwu4
Xy9952CzF6g/qf9dj4buJpg+l6cky49BE66+DfUFKfhp5i87aCkKoTzGjKKCEubPiqZk5FMHwFsI
8TZbVtr0JMl5h1FCDx/eCTqWx+6X//3DEnKKQ0lWw4ag5ujPgHvKlagFuEZ8ZDvLtWtRgbPKE/ci
kG2meMKYsNFNm5hXgm9S4MjZ/qiCzhkidD+ekhbPJmtcoT0PSep0oOUaajQl1PFm5rbUIHmSH7S1
MRgek2Ky6FBzuCtxr/45yVBS5DpyQnmRiTxzpI9U1C7/EWg+Se2wyiEfnMgxd7GtA/fEfzOJ8OIX
BAll/SxifUpfNjNC/sfvfHJuLfMaFI0qpzxRnGLQPuQhT6xPenbuWRkIIzr/MP1qjOplSNiYyPkb
q7SeqjZ5wVv2SJHp6eZ6arw1LIvHQOa3Ah0TsH96QmfXYEbTls1haG0jInFZI2pQEuBKQExDtWA2
bPJPmUflffnTBXkghkOXOaOcTCkoJzlKulINjM4Eok7HGFcb7gxY7rCR2aXcMuPBq6FYNsFbOq9e
J0WHiSjOSNk5ThJsDXY64TkKfCE4rXIwqIlq42J35W7Cvwx461Qwk3UPzSlknhcZXp8iOBLDSVaa
yLAWGrCyr/sIVNNknx9aSAPRPsMgOZkawDEsDgQ8IcX85gQfVfpSM3UgLOYgaEWgTa2TedKIX1vD
ogCccmU4K5iE1nAqe7K0Xmx7uwaM+CnijP8pxjPWtqoVCwZ1BpFWM9LEqDzu2U38YDrrf9b6T34g
hQw3STuupXKqtXF+BHijWvn/J1nrAPyBdIYe3ZzRynrY4Xv6sftLIkr6M2PbLaBbI+8UTG+s7IDW
t6ol4JfwQC6bpYbN+Z8wgpdyWZgugzwd++3YzO8iDuHWBOHswECXUr+qjXZpiZ0iMwI0RcfjEKsW
Q7md2HcoiegkXkwHC8PEcXjgpwcWr26MoGc6uwDWg46TWqvQyIBGZ7vZFGwjE3hQVoJO9CqDqefC
iup2IOV8MYeK2D+Pq2O5tWluuGTn5sZl9aLcL6nYbVDzkYMzwna5FoBxMsLV6FG5CTKNUnOT8d+n
QBk6Q0VC4E6aPtTHFVHScl2S8FNS0i9XF34RX/++GogY+ozZ/cPyUmTKH5ZZyjA0mDcUGZ4vfH7V
h7v6whPSqQMGJZ9KqTDyO9ct2mRZyL5diFSD2uVpn2wcZ8nPKpbkHBMop6CPIl7kDrfAIYnQwRkm
3IF+oWzgcukXvIVV6F2PlAzrJsNWQQpb6x3yMCTlen3mvxJr8Ha1N6+f5qHV7s8xoAL+WMm5T1Qg
HaqW4OXo9wL0yUjOSeqQLzJRgxTABNmifcTYNbES+bV1hWDy1amADBuFobPj+z5IcqAUKx4EH70N
rgpy+6cp4OgvQa00HE0zhseaZvAcxNltv/nZ7loaXSvCGzYNEBGmIkF4gmjIm0YsDg+tQ0NC9nX5
LxHN9x5Lc2HYbjKIAEkUNSU9faNlzI/52QphqDZ37X/mJ4bbtN2eY5DlpwrcetYghqdsQGLGBHzu
HJtpyfAyt2FIMgAzApOkVSy83F6qkrLSxP4hN7Noc09WEbIyNsZT5lHa4+3J6Fpkl8ncmjdU3E9Y
Vhl9wpjMzdFzudmlHVzBGp667Qp/zW1QDI9pxwUMT0qWzMgYPkuv70VTzgOKJ3ONK6SCwlR6MF/4
xRfhLpjxyre11m1BB4i+/KE+9/RlvBGpCyoUuT+CIWnkrPyEbiDWw6Gojb5dWZ6C0iLj7JiWkd5y
f3tE9iTEImA4rJ8tmO3BJAbyBTzMUQJGhoAkHHNumYV5x2vWPymwQoAbr7A+Gf/wl+gx5DZg/3/e
2ARycNRSwxCrlG/ybWNlWp4Vw4OpaGUBGznofbSueEHNTPBEmztA+ZK2e+kubwLOCvpamA4ErqW1
VcKfGKM0K/XnrEEyO15BFiRrmP20AxcX/Kb05E5iDTH8RfwCF9JYi4Gz7pKwETqPUzW7xBq1saxr
0hUAwnyfK/Xs1d/gUYDTBtK19/KkFUDcG+vmMKngqoWePrIIkurIKSq/LRxfNYSOnGO9T+gTIbtw
YT1IKezbyhvYpv019lG4yvntSNek6Pw21/N2YhafO9KdbeoTJQRPXPwiZpDmhxc+wwLLBUtZx8n+
Lzkz6ai/LcbN1RC3wvvjAlEKIiHTIt0dbITEXdkvEljdtQ4TxJ4rBgE7JA3cZpxODC8NgEZpgJ4s
sqPpP9wvtOyw29uW5DSsaCXadCn8ePod5hL5+qAeZSaGZ6e8CkyNiq20XjrmsFYAuQIO0Q/q9cZ5
Qk0Uj4KEbDudh9/77nWN1eiPA911owRK2jgylgc6K1mv3tI0N+pJtl5SfHvnLJwsF9MVEnbJmCah
MhChSxTnLOzf5stb+05S//BS8BKAy1jg/YMiGDM5ALF1MAnzXd9mBuqKz9POkDYS8/Xz8+6eqoXb
RJLQrasy8XKIJX8KnwfZL2t4YGqubuu+TaHA5QFlvrvugyxBg5SCtGymyysjVWfmRCmacsx493f3
MJl1h94fztsbceSHLmW+v+nCy/kbhIk6V1NWVXP5eldSGe6vvAk+T0ZMKUciew/EuBNmBQ8YqOJx
s0msmKfHLOcZbkiVW01XQMeqGE9OxgkYLDU6NW51uZSuN6mL+vEaemxcwxDskBF6dz14r9sYMAN0
djrVzOE0nRt3rsOmiETlemfiaQowb2FLZQ1odWBQP/C8gUd83qIGSgG+WTc1rwK2HTVYBmEyNOEA
dNwsdb6ef1QgRFD256FiWykM6jvGjRpNNerFDoLvJWrmOAq1ZXSSHah69cF8ykrYzj/WvYFeFe5T
JNsYhO7jM432oTPp3cHxMbtQx6gTI73tl/gCMrRPw/Ok4NQ6EVQ8SiRv9jW/7GzhKBJqUOzE5x4H
k+d7s+FfSbu0a2YBU2h9VzNQnnzDejR1cZ+cWa2hcXNUyLtz4sqUmfUdVnCYUex1lJw/7Gvj6yvU
WMe55qjxh2ocID6UQkR+5L1+F9SUZrNSZm6DJI6WQl4mam0F4cqXASviIxTP6UgmLvrc/tKwNq1v
EygW2MOw8Ngkm8VVTmNT9RFTNi7Y9yfEmyZMZ/HniDF5ZURFMvsauBdDSic4MANEBOEcsYi639b7
XkLTShMD3Ky9LWX2/FcS6OHFKwyvjKGWyQLt4pQ3iLZVHhDq7b9K3/rW4ySYZiWIwCXqSJkoc1MT
WU5ATyEiRphKptCk0Yt/2w4sHXRA2vN98T95YYGVK4l4glNnrIhKJoNdvW3FCm6ko5ylAjoovGa/
VjKif1iqeyTbh5EFA23mlkJx8te/E/euN76mbgLhv7HzEIEZyAGISjjvvE/xGrYN8p6LIDrURuAi
TsaV/eunj1xtsjHQ3Q0kyz9PDoXsrjwlS1XPkX9UG1T5JkIzvK/19RyN0YXrRffs1T1SJXv8js/m
6wtCZwuYFV8tnxTIozpBLjghJO6GMO0k2GalBvkjZjklIVD9CBf3H8Oc7hD6mMQxPBMa4iSRfJjn
IvqcTjexIliAzFlCFLW8obLhVaY6zPe5xIeL407pEYd0oQMQgIhuCVh78tz7/405DPpvdlfw6euM
v+h3zjPJXZGk9uyJ9PMpyQBycKH34PhLla0kd9zDb9xcAESjLQbMO47fVEjeO/xjpci9FQbKyHLP
pNKaKGqNT4i0AXfpws+UjnnL1C3nfNznB6cyQJLIbO8mfBSd2FnE4paPXp2g7isB9PmHostld3jv
uJbFVzTjZYc9poNQRW15eAyl6kNXmi42Qw7HJXQlH+/taFUhlU+5k0wHlpEbQgc3KpkZ6n0847E+
iEdqC7+DutlwlYqm+H5TYtUAJoQ3DlgSmpoSMMoQFD6znF4ej2DKt5A4B6dG7LhbWl3V/ZaF10mz
6wUWFXvVd2KLB436uWeEkcvUHgOMZgyMuMiE1FqRlARr5ZZ/vmUwf0WqgV5LoTLVofNggSqHz0vy
xlrbliDIIjfnSkzE7fdTIBysygRF7DD2M8ABBVgfq7q+pCOx0a1MqfLQV2FxLEwnjnhDd+dX3iAq
9WCcns+Nl93Jimhn+Z6ZIW/u2JoRlJVOPturqcMRiARWEFEb31ihe4HDxG7agO1H9HrRoXTjgE8c
yd0s58/u7jKjofG5dMwz0AQhUwHUg2kVC6gSPd0or3ag2N6L577KnALEUatB3oTs55CPjVpDW3ps
uU7ozSYmT5aWQIaLYgT+XwAVl9fcl/7h6oHkjkhnpQ7hIBZMDUUNKe+lMpJMiRjux4WldvZPdmNm
dwX3GmXM03TlE+yMg+u3HWjevUByz5vj70hFoGhVy+P2rIcHf3GHWv6ONSCrTWqXPWiOfQcfe9T1
6uAPqRq9PeOrPxNngkRt29QqEpUpxrWtSFuXA8lrNDt92EdR0O0L2slTcVMpSUj/I7hnUSoSZ3m2
JCXZ8qgddXyq2f3imUrS+L/Q8IpAyRteWRQOMe5gFCoj04sLzrBcB3cycRpICUdbovXxFjbYtcem
dlDLXn6fgxfej5mI0fguX/PXJ0Vx08k1K9hnjIIzFCiXtGzh+sRJtbLXuZikUbjHL7Lt0S13wxmC
L/54GaiRUT5oA4LIyOhwj03V8Z1I1pLNoeZdu2MdSF2YI8dMGlGHjTr+pfSat2hPgc6IOCNvEGlq
DPufJqsJRnRHx+/lQnYzoFhfeVNtMpqb3SRBL8/WMlBV9MVN8lBzRpyKQFG2KCLG/wJqjYPt4UQV
ztpxEasTmxowUpYW3la+rKlB7N65qxbE20nuat0Mjwjft4dpdV9IG8rADpXSWiJcvQu62JbemWLt
MHq4YEaEp3V6+NhRWe+n2GayjVp+fP5wqI5lcKXIX/cCFv3MPlEjYfPSw3HrUqFwL5hdfO5O37hD
IpEl1O91vIL7IYJnJq81orL+HsAUATrLMr8sijbmQc9hnQuggg57xGw6ntYhfTnm1LyM6s+3wg0c
vsPGvSvi63fMiNaBB+J0Ee14C7ykMbu3o+9Nvg2YuFKi2b1dAKfxXpJUupdMkSis1Xd0D+la6/ma
c9zGtiA++/diw233YTJ0MkSvQWpYl0awrpcR4QlR31LbkbEunZCb3p9QGZNLrw+0YQIzj2otzLcj
2r3X18mWgQ2nlcWBMZGqJfC4fD4Z6/wmG4jzpJ3PafMxsFBiRWugxX0VoBv6Bc0c2u61sVg9YVVi
munP3XIGzPe/TICfi77PW9Pxs/5ymzHgHHZTmCcH515XiM8EZn52Ji5miZfHTEfcY+VtVdesKcY/
0Wi8bhcAt2v/KVKEkOShtjziu/VYUVScSbJ9IzgZfYkmkZ4SwbMGZoke/cw1v6gBT+2NbTOaycl4
NTIZ7k0D7YX2CWLOEkIrD6bsRnFzDL1yQaP1FlolR9FWlJH/uX82umCeKxQmrccwyJjL5uCxJim/
/Nmh/XpXM2sFCboCszTm/z4HE1QduzwJ30e9l+yPB2/fxIPdQhXa53oDEQR8RAOai9tRjjEcQkcc
JfCAeltwLwYVpy/llLBaZHvwkYoXiU5uo5DlkNr/YXIzedxGjaFQwv8p3cK/Ou7tGONgON0C0RhN
qvOvst8avkvihiWOwT+IwM6MmGm1N74wSYXbQMP7efjvwVnVYhxc3XQ37cGKx/2sTacuzdO/oX5L
L/Qb8/Jv4Z1UceoU/XPT73M4gS28onhU8jjWo0dXc1It/yTQe3NxJnSxnEXavKZxjggN70HT+i8M
w1+dRt9lqg5psTe/sBVhGqc0YfREUca1ih8omX+AAGvwpi3pAW957mJjVQGK7Dg8P/UW9MbNQT2z
vZqeS/lmRObCdN/cuk1ErOpm+/4p/46wXETxynkreOygZdcnho198/zcZDNVpvgKsUcGS0ykt0ID
olwaUYQ6dBOVdqY4B7/ugikZS5EhiDCIh2c/5mEtJr1yqmRg1yyf/QB+HNQzZEduq1SNFW0scMBo
3xW3z2t3IaTH6IrgNsKGQaFYTwGosnjO7XVAYJa0LMusV01BG2tYoOn1FsDL1niRmhm1gWU/Ah05
AEMcO7St06odoj0mQ0e3Hi1M5iVJ+uqKWuIabRjvqj4lIy4g9SRY/c+UxSbrtpHlhHDhGmOkp6mp
0KsIFPgAXU/AdvNzR3lY7qQbMILJEcxeb7cpNtcmQ52WUXbVjuybblpZd/IPayR6tqkCUdUbEUFW
aan4dQPVjIUuqGXYUGpgMWhw76CaI/QxDuNjgZ8IHsunmtDC9jvEfyxhY5kLKrKUF1Lt0hLcIVA8
FhpJ6jSb3+onNKM3FkKhFAQx2+QRRernlLb42XnJvFUx7JaUMbRa02w5YjdAuHH0/APHG7YG0HBq
lLfh7bnck4lX9PfBd/u6p51NjfT0Ty2KIktHgyYVKlWzurMQ6ordokO2UvfKPh25Cc9a/1w49fP8
oH0sZYX8tFbQ2ho+pTP2yIlbKbHhVr+2N1/Fj2Hdvl+KpgvaLmvWSKuSFmBaq722ru3TnyP/gr2U
GgMk2ioEc7Rhs/eKEWiKj/fO44mF0f+aGYKVi6qJA2Heo0hBryDGmKYzl3BNA044hymni8S4nkIW
hR8unkjNpf1zZ6f0/NO45+wRrnUJJ6rSMYyhZBsRHdjrbw6ZDbYdZz6yxgZcbkoFtpltpdARVxW2
HkKs64knSZAqHCfCkZEWAPLC/7RlqLhQbSDg/OuVJ8Qxj5YT23XRO7n6yh4jpvaEu/zkX2K0Y1qy
np2Dd84I7iU/pXYuH3Dhih368l+NJYcJNGKPGhnd9NNtP7/YOrlJrUkW9zFP8rw30UnIOGw6+Fp5
WBon6+3amHoWXAyeAEv/intXnoi6AOfHI806ICrQ5ow/LGlmFv0c7yV0ytBHaIgcLV/GWw0kl3Vu
EIwhdYE0svoNfqtSnRjYruNT2B+eVuX6NgLeXyd/LBSpegyJYLRClSO79HDs36W2wVrpeAavNX3i
LJv94De7wx3QL/Py53/XlOi6WXTEgdaUfn12vjznpW053wu0+hPqn9POAaIR1EwX9Bin0Op2soBL
LRi3BkNRQV42p3WJHlN7NkTY+VHILqSf5O8xGtqlc6+42UPpk8mmvBxPW5dtW5uelDwVtfdZTcC+
IGShoxaFo3YvSHHbG8TcT7sy4dboudivmpKQIzhl4eFWOMPJE6UpsYlZGkTH9hO2b5nGwxQuaZBf
gFZU9CMUtBP0E7JKsd33oekp1GvRRnfocn/s2Rm846ETsclKrI2ocmjP+M93XkgztDIWFzQmtRSS
i6F0i+aqyzajVw8MnkiLRYVJdd97LamT/Z/M8dKiZ6bqyqMwMrwm+1W0IZ5P57D7QB7I71w1/Izc
e2sDKvFjOaF7aFE/8vmdJPOdUEopG6drWcD9dMweqR3YFYtA3BtznscwUkEKxGTsoPIqa1HBGs2d
bpWxmBUj5TBJyilu6N91zppjJo9lAeHgFr/QIaaj2qbbW4oJDLKyNtLW/+mJtKnDCc3zFuvGznPj
r3R5SoXrMPQCtluzb6HMaiX5cnkvwV8PmCciVsbKoFYue3WjuDT+9iWMyQuM6BnWvl5R98eHlFHu
nghADOpFTmzuP+g76EtBUYLmBTkmTcfaElBBrYOXfbUSjBb4hn0Gr/7JVNju92F03V3K60++IAyS
iXWaTR6jX/Uvxf+m+QOkTGQpGOXt5Y8Slj4QnoS5zky0Kwjxc6IdA9t6jNc2Q7amV0GqX8Wl4KfL
PTzdDya8bGWTLkHBRI7G+65Az3Q8/HNzt93DzM8jLmL6vu6WXE4U0WsGFsN4w0Ya0n6Gk49aEvPW
KvTxMmPjci6GYbR1SNRq+mt0n+5VXFF7BG57uqCqUlj8pftwunwCuAvtw8pQky7XT1Z6CnB16EQZ
cIzMneZYayk0rHY1ljfEWt02nDbMWCP1W7NPjP2YjkboY7gV/L1FnJqfMwQriNFO2UjtJ02/YOrg
3f7ZjROp80+OyunP2VJUc02S77yh6tUBuU4Mp+eWDRQ6dlQPVeEkgeA1NAucMFOxoT9FTJW80V/r
ZcsdcLVqYQchqSJgfclT1rxwITrSA5IkR2xDEjBby9Fcp0QvXUqIcg1dAe+5Zr3hRH6uOmXVYRio
joJHic+5eqZeA0i9aoHFhK10fJPkJkHZdRP3ftW1/AYUbE2KrliYW8s+7gRkJTRUDkklDnMET3mL
E1S+WpibhsLdoM67enQUnPJ4qeI2XMjvj3V87sUrzbDy5qBGXz0iU+ibpGvP34FI+epY3xGA+uJ3
k3wxv4CwkyrQRU5aaLizht6TsZBnwXaRxK5otJdAQZz4nNwusM4sZ3F864vv18KPbur12o1hkLY+
3wCOLtF39BrV/eotmR173L1Itu2DE8NUeSjOfWRvRpVYnw9FgAavyuNOw68s+r8VHhKiSAr1cEsZ
aJL0qEc9oLnz+UoRN5OiHQfe/4syxJK6cmIPUopu2r/bm/9Lh3aTSXLpKPiXeLXt3xUzaFv5fGDU
B0mb7l1fJna+kxNDlGhxCbgzYvjhtWhlbidQo0gHEMWfz0JGY/eNmpyQPQcioqnIjfNW9nztAocW
/SIlBqasejTZdPqRR1YVS/1LrRujv2kJl4cUPLsXj+319JCzYFO36cVU5wbpJkesGaS8BUGb+Xn2
Tuwpy7yiMxIR6c+wc0Klg6QiSmPpFGkyt/CsVIzXBiOqP8EHMO8GA7xOi90+gxpr2eFL/9ZStdfW
a++WW08YgqYf9qsSIaygc3NPK9G+rSGXNZXzcHZQ/alseT7vj1uEYYKPMBc4Pti5MF3F0DBD2jjn
1oI8oDP6F1URaWIjewFQ8rtcnpUn3a+IUZpJyuWhE2Rddanxet8+SvXsUxR5i6ZaWByRjx+avlzp
S6ymSmbdLftjOu8q0fUXEZSS9FIHEP6zzyubj7b6U6UXKoRSJG19ZMHinTe/7Xexb7OCaAWOcudY
szeyZtl3Iq/KVW8UilIzh2pLWY0Cm0+QsQbu1JM0hudotRe9rpxpNq6yc8Bug+hq8Xc+o+/Nm4Pu
Ilx+xsCCoZtKA8vhQzi0IgeDWh5aXHdysvmYYanHZI4ukXupuTJjsUMOVH6LTVYEJkXL7pSklccn
MIYTBPS/KVeNeVhXVXKis96R121twd0t+pQ6WI/l6FCUnjnwQGVjvVaVo7LX5c23LB/Ue9kw2UKR
e6B1Hx89jwUtCdxctnbDttxJyCwWfkFArANeEhdgEnFl3MWVl7RmoAq57yIcybQRiABeYkVI5Kwc
VA68sxkMC2pnl88CS+lMUJKG8+fZ9Fw+hK88GwlnQZCGeQSx1wYdJvDXncikUWkjjmuloP4wlkd5
klCfToqhQLSy5gF0MIAmyCpT9Vlc6NST+sF62TrL+415+E6fHjum67LawHT4CawyHWUyOaBUlpbE
y9ArTxjoHoMNyx6lLgxoODVD+LEP8vDsdzd4HkkcJZasLxGYjLC6KksxClN4Jn69OuuOdK9OkwBR
/4IwvED6gcN5Ws8cPOIXtuIqVSnoChZmOc9k8+yqIgWNgKouZ+8BebVDxWKUYSPkwEkgEa1oAJ1i
r8b3glXdo/Fc6ZkehZ2ZOdqWDRScyBB+Noofin5zYe9wI76Q7cmsItLyrUn+z+snyNyJlyUkO7NP
VFP5E8CZQMJuPjV/AVUtKDebxg0jNaILfiLeiZV3ViFnURBduTUSFVBDQLdfSZicXEALHSfXo4dz
fqsxKoC0En2x2XJZRa65smPo5a5A7oGZiVgj+yvoXdWHMnuslUpkBRbh+CH2i4Hj84sKPyytZPw7
bOb1tbJaMt4LsF2UGSyO8pTaDFuuVBG1XqVMeTZmNKoJEP6lSSOoVM7B/VOMcdHBRJP3HP/RnbHU
FJMDyHX+p8DmHjd9eP/UnLYKhPkzc60DE46+ieXi7w1FHxt3NduDdMRNVZM12RbRpT0/22bwFoaZ
A+Xc9VIk9n4cfQhx/kIMUZG1y8k7tJmBG5And7Gxon4YxHO8hbT6ZkGIO2zCe/oLvGbJdN0y+tpH
LpDZFEbc4r2ucfT4nEN4vxRfA+rZhj5PVK2LdKOjF5LNsBvXV1XGJzNe3SC+A2XdXBRC9eVlBis7
ULP0sC+gsuxaYwWifwTMFUtFAc5uWPTmpJThWe5ka57WAmroqrpbfb5xyqQt/w2oPWxjlVZKdj4R
1h5Q1CZtMNPowe0iN6uxO2a69eKK8wpojB5Nzmp9rE2AQVxJrhIYhDFPwPltCuJPj8UXIFqwTpDS
wPnYmjafIURbRImImsUlRAWpg8qkvQVsuu08RWwtWqiGOzACnhyL2oAe8kIlnw/13EZA7+ZRWtbt
JFuFZr9bdzsIstkxJr1cgRiBtjhZ4skTHkh1/r7rAeziXZ8uWcvaWy/nVHpth7bCUzNbhJ15dozZ
3Hr9vvyNfErR6hqN87RWGhPiXGCBLSNYQwrfpBn/B0qzDrMDnMR/t7cc0SZXG8u/6wr3VpNu1HEA
t6HOWC05UVCXwrr9DGqJgrh5DCBuGEmfTauP9uadQVMW43yipKzkfKhpFCpLPAClKhEbFhJbJOA4
gSgGcN1VsLxnojj8XxHdXT5+8ZEK3IlVMmLf9jueQFHsNJO783Q+dEXww4CnakXXh6gOp49GzDaf
HSWC0jrClNNLefLeTfme6glCs0XamuL9I1fW+JbKzVdfQGYRrGbvbYuqUDxAqIVWo4EXBLSr6+gj
rh+1wSHue+QGSE1cHaRcUCRIxqtaItIyg+oNUWJLTjPn2Z13xxvRq5MDDzHIgjyLTzBwoHCLiu0v
R8TtZuLd7Y9fW871AR44riFeGmPC3OmNwhHuRICK7Dw1SdRFKk9VpQOQEy+lK2uOiamkLqxzYvjb
eQhJonf1/7AW6krD1rp8vggWZlFGbae0ESR4RXt8jA+ppSW68kdGtUxWxzb1l0OHG/RKyClo0g0I
R4wd1CCEW9fJiKDJtSFZSpdQ18iq8ptpscRqvLNCCni9QT9mMXxi4ubYATLm08+yLt43ONx8b3Xo
ogD5spM331JkQZxkVC05cgiBMssxPpkg/6dzNb21pz9PhPAl1zj6RIMewdP+Ihig/adYWwCp768H
xiJrLyi6PUReXK3Gv90OUJgPLXTia8j8Qb3EEq6Pj3MeItzVrtUsJRC1dhkk0xFUhEOCcHnbmKw4
H8uF/QEEfXbDJO3fggr4saf1DEywoZWTCsoKK2c5pJybWk3sClkZWCjBJ0yOE0TaS1cy9LuP9JAO
HCxvDadb459oATyH9m16QXb0jRveyffTzazWbcGXdvg2u1emoYPVeiefRuVuQGeQFmPo2riQs7k/
3PaEf/ctZU8aHX1eVXKvz5um0KSytTAPsAFgbD9WvogbHzkbfHieU58cqbxA3jujB/Rz84VoFKFE
9rg1XqJomi0a83BZZyZr4wiw7j1N9eY1s9V0qOYbHqH+JEo3OPkfYFm7lMTkix+gxtOc83ZLdCBw
1mpjNvBP8JTc3t7Ap1ZWiWHrgo95NL3wdHKoYVi3a5a/3P5+zfZzh6aoNykJ1bif8Zx3S1NRNT3c
yn9YQ9qBSRMh/5x9Jh/GycuObEtsLgYl8qTczdjMiC4/RBk3e/0lQq0hiT/E3z6eBJPhAczcnVvf
drFfj86PVEDDL34kTgKLVHBnZ+EvWcD3kbxdIFlC5w1Nl7VLST9XJdkvQWqDkFdHtGNf53lI1Bcd
CcQEyFVIH431PJGQuhCVQi5U3u5E/qDzL7v1GgeY4P5DnvuilZUaQoNsmyKv0Xe91BgssThl4/U3
hkYk/H/fOC26CWGAr7j3LQvezFGzrAr0jZ13dn6Tz8922DR2EnbNmSySV+Abcpoc75EY6tvr/VkN
Gvc6sZKh8mO7vcRztqLxFzM1iu2ijqqcM2NUGs6dahNujCwXRLudZaV5xnU+ofhihAE2vIjlacdd
jgoKD53rOGt/qjIHbzvi21BT7ns/qW3fTLli6YPFs/VqnyTjhJ5vfqWlB6JQhjDDz1SThLCyMwCs
Lmn1cV5/JUPSDavb801EVZiEj5pXmW25ohAnX6Y1jrUr3iZtXrTqOTbGlYEujJy1T/V1CwU6pP0Z
FBrbg7ojEujgv/vf46WDoV5W+rOw9gnGGNNQIcgYleyxxYw5j8hAE48NN1GLYsPf9UCPaHK8Xsiy
EwuuZ4zLJ75HJh1BgPPNpjE0HB+JgrJ1GQMR4cjK37ymQ/BGZxZ/A/Ck4H04OLDu159XDFRTEgiM
AjoXSlQ1c4mAINiotClhjNxaCimKF84FsYJ2X+Uk7nCpDHcWrIGzfuTIy//pCqSGkqMi7t5ZfzYC
OycEW4AS4NoNbbG0+dA+MzvdhdHyUh0gQLvtNwVKFPAZab7TLOHVMasoQZ0GLLSDuZpvA1ISsmNH
H8k44Kxose2nsx+xIEBuNKrxIa6lJHZ19hvLwIOAq/+w7l294FgoJtO4IVm/DxyA+s29M039+KBO
D/10jAGFDlv2PEHpxIEsSKl7BKScD3k6NkKBc6jXIf/TIo6f1vl7QJE/hIYkUbEVFpuLw2gPJ/4L
s1KU/ARsut2x31AdNiFjvlSWbW6CfSrFv3HvfMjmFhPEmLBFGKeBNymBRGajd8A9QM6ClC/vLBj3
r6BMR4jMLkxDAoL1DiVX0kZHw5MuFqRpWHL1Zx9QkNcOUO+HZ9cfbHeHNSV3XpbMwjnfOSGtL9tP
yprucR3E+lSpCm/5a2sgXrG0EgyX2RWLkNDKKMAeKRx/7imrxhjn2oeVjJFyhF/uADWKCjEc0iy+
yrJyOv7Dm6uyaHpiezdCUjYT4zGDeC7yQX2ABb/eN026qmfJ0RZHzxjeJn0BvoMcHQQObSsBTQPw
kpMw7LTyRCDain5yriIlM5+cswfITObym+nY4dNr5Efi1tsvMnPaZgJ1kMJfrhUlxb9HSPRpoGm6
1eldxQvZVCxfoIARG2y7jcaiGl7vqHivdJWCOzxQ6luzdALHUCzsfp3D99d5p8Ewb45M7HjP+Ivp
oqeonLWjfNLOZjY6HwerB3b6xFOoMOZs3MsXYkBhEJ/mGe7I9qXbBvmZwNFWsIVP2NMeV1Zyxtrm
61D0vE1IJXPAHl8FCoOaQhek0P7Ey0YAYElq0D3FT0Am63g/T+ssxAPMCwQKqNB+B6/nPndDqer5
/mBblL47kAvWZkrfhnfN4VUsprki+/seX2ZQCgHyq0fCGPU3Jo/xEjcfn2HM6AecuqrH452+J3Y4
uuMR/JzuCj3NbZRcCLqh76eWkdkRTAaFIR3jKXWpFy4sljkXA0Lm8oIPLnHM6Dw7yTBEG73MPAQq
c1nPd9fKZfE7op0yqkFBpVvcEFFrCMhQ0sUgpiX86IAvg+W5hGSUldlMDPAxgHLYIeCPhHQG6Psv
w5Eyl/o7Bg+w2zax239E319gSxHJr09ebMU5gYeLxjfaBPDk7VOPEOYBdkiZLtNtXrviZYSlWTbB
0CTXzwsHFn9+Rzxlv+FiuKIard1AKIVq8nELYW3cZMfFohcoUSKZUuaEBEWwMwi6k+1O21TGsj6t
CFilsz0iWiQJPACyPGwIVqmVpJnxWNbRHvdYlFnea1cQf5C7Gsqa0R5aAyvgMuQIbwuTzpkpqrMi
GmAHrYTp7yf1P54M+dWm6fvQOSvs4uA1m1yr8WgI04bkVdRTJuyUPC4PrvSVbDlymjsk6ZcZw3Y0
tEI7dx7Cr4fFal9g6OOhqpQt/6+anbKp3c2M7kgnmXimqsuJtjo/EmkzO4Oolk2nzcg1zAw7J2ED
HsvkH8eeVV2Sx8QSbbmNWS4w9cZuYM33y6U8dc0zwDOOrvFIXzzgKXD5t7RoIt/Cb9y87cLJoD/t
Z3RWFEiRW0GE/a2Gl8y19rYdTiPWtA/4o2xrsWoVMjJp3w1K9ikkLoEk6CnPUHj1ZpWHU7At+So1
Ru0LvbgQ2SeWzSLRlzALh46Aw5CP97yuEji+5mGstrKSB/4SfaTx81LhcbZPcfGF4j28u+Y8u0pX
j0n6IEkMZkP293KOt0xdN7sCiInPoLRlJ9mukCa6YV9FxsFswzBZtA7NhFZvx1mxIQ4aafW3O/fm
RRq/BmJ2kZiM9bs4fmj/K3FjX91A3mqEXyLaAqw6Yx+fGFar8Geq38gJE1USO36Ikqv3h5bdcijw
zlVe1ETJzl1fIuVQDxlP7qQeEoJ8BiC3pGCDjAZkYVbVrmVat0WPY9grzbpniZWbdVSWXj43zv3K
0e5ww9hrMNF10xpGNyLzZyTo4oMpL0eUB0+8tcwI4L+/YYDP7oZ1IEePtc39d+AjZ9loeHHKugZa
BUvO6uElwCKf8BeZCsqSSVyXCbCNBtSO4qCC7zY6WkvEnqCHsRaTye47qh4LyscoCedF2if8MJEQ
DGFUFh+DXe8jQGyjutOO2PqY+cnGEnSoWMrbYOvPWmYyGvWazXIVq1EQ8DPZ4vWK54TkTD7Mbb73
k3+M7Z6MwIPkIFhf4k6R7fp3mzcFqgTRkbMNZIuLzH5pVRpBqjFK3VTZ63sBSGhaj4rLeGMs5lMs
DRkqAq6/FfGUrOcudolo77VChu2iJUn+3Xlcl2kCPlpFGuEgxHENyr4qEStLbx6ZiU/YqX0EWSBM
0YipbfD5T2Q9M29omBV7tsqi316zSkeRpk/KIEO0in3UYNOd9OR9DKBlMLF0mcWOQoV+zojc3EE2
5SNorbqC9J3NBaTe4jJZCwAY8SJx8eoW0qfYyJeSo/6iGPBQcmXwsRTB7kFxk6AqVCOaiW3fhhal
WaDvoL+2wsM/c04I9HHagH4onqCyrxMwHAPg/ViYQyLCLueJKOaa2F7s6ASDl7jhs4/JJgG1Jd5A
ykmnrk2/XqyKBI8ujNzPB5pmT5MbBjICnUlO8MsdV09VjW8sy6vxtksgMn4WtaxUgFHPxk6/D7pR
urKP11A9tXLvTqLw3FdQx+l39L45HwYvcOnmuuuGhxNaH1r3JmMIUFWF3ufSdYyqS+9380UJgmwg
p7CzImYVMYgi+u33hjJDwcmptymJKKFbQ60KZ19pMuLznPjyARetUDUEkHEgsep4UG8HqFqA3QDa
JjILnSFWsKY8Q0I63G+p4QDDyRTJ0Es0BcSmje+/YOlqZFaMwRDM33FzlpcMTv0ClIMNGxQ9OJQ/
J0o/JwlEyphLHcB42EO9MJBNKEVF0deMS/t1y5ia7H4gk3xULapvih6tkfsNTK7bonlCYK4TzCsG
qdmX5ubolhUdwlb3TNPqr+gphveyWK45y/0obcJSz0nV6ARODQcldhg4YNHkSA1rcg5RoqXcBxAp
ytTgN+ll++D0NWc4b3ezo5VqvmhPwunQVltk77I+NiwV6//C/ZMPsQcon2J6LvF6hKHGVQYUxL2B
7rBoT0ndoykSEIqxl2pgXkZk45nI8Ai+HZjRX53svGxSlRKTIJtiOFGxlHU7OsR769/ttti8sXoJ
2b1pud9S9QNhb8ZKOD59fkKCExe+5Sb7dpGdQSwFdDbogPCeauAI5PonYYwrP1q2TiOlOMzGD2As
vzkl5/+l+fV2PXw2HNoNTLO3Q68kcfcraMNHMdOkHbOdl2Qsnns7ZTfGnthKWpjHGqANlbbYQJUJ
TLX5E4tb6aeOasHoa9ZgGhFfRK0GNudBfGUuyfpAmfshN8SyFB9oDunI5sDzfpXP4vq3Y/QC6f8c
S61U/uZZvLccMYhZ6lzEcXfDa+V33RLzLlCEpPjrHJ3SGUZ+EB5xXcJeepcC1jxDcC0XHjXZpygj
CV9gqOA80b0PyMT3XQQIxxGB5oqkGZN/9j3+j05Ld/KzE61NO2xLvGEQ++ntHiGM8lM12EDQiIb0
3VJNXp2CHTAUIE15ncAMqFeDVfP5npSmJBx9w08hZzuAUuHLA36FOF+O5xuwjd7D5hUX1M0aqPpp
W0RpgzJ9xkKFD1R/7vmsW21FQeGpdo8zvvpWFo2m41Lsdt2PF2K2uL6DUs/RIg3j4yn4R7W5Ok92
hS7Djpln7eZTBXrBzc4aUQVls7yFtTfq20D/FgKOOxR8JdNzvQ7nkiDpf55Bq3dPgDGwiBCoFFDx
eklDQq5rr99g8VX/G2YirxWAkIgQzIdzoc6Qy9kvuwxiT1VC7+5wRsqAGQKx4EErv0bkRmz68fob
E9ncyvoWaVCJy8pMB/YoLL1t37Iq+UeGCykkO6HHV9AEHHkAN+YaAhpFeqUB1NZHyCgu0SU9wpn1
izYTPhm9rCFItP7hLRuZO02NYjLakNIpdY3w8FRnxo2M6eWFtSUdeDqDLL0dAvATS7OEO4WWODMv
exYjFwa8NInXEmQo8aFlMVTpOA47ASynjGlVhaPR664RWLYpTBiItZzZeANlA4LwRD/X1xjg3RG+
fbupZD2uLLLvJMYmm7ee0zzyS7DqT6IwAWjO1+HVfQGvJ+JBEQJcENGnhD9acpT0OBiuXsI3GhfV
4KIQVtLdgk6nNzN0n8h/DW2v2MlPmbGu2qXW2urQ2WpJlVHvQ+xwK4xn36u+ENXaHDNDiD2rq5hy
000BqRTnzu6BXyr3sVgkRpMHDBsvz1TDeca8itfyYtm2VpSbZ5ONG9CLIYdPadKKUQUyTOCMScCp
7zpS7B9nlLYSoVm5DrwTGUiL1R6jeokO9iuoV3TQGSbFi8eAJBauQueQ5GLyM8JVyPS4mXkQUTo4
0UcvQXnpniCIGYPQG1/vxAqBdZVau4zizzAyWcdDDPVroPE92UEGrtOO+0tlYdzPZLN5VLZ4nD4O
CHDfEHJWUwbAkIw2G+cJy75kNPZtuZJRxm9C4kWLyqeQQnfG/Nvi/vbIjPabAQrLwsR6QpoZkoDH
M7hp3AXSPmNdNTV4QlBRVKY9Nyw+HRNmBIWyayUfDVSrpQ+Vn0bdYhyi1aCo/t7Waz5xvQji8tsE
x9CJlO9o1QaXYI4xjUwyurLqQYo2wfubig98xZ7V8gp/XsbEPpla8c70QxSoTwJk0pR6vys8JFHq
tr62ut8aVeStiReUTyUBQkThKR4PkdIYVk7bfpityiJPSx2cxYwod3wBNPso51e4r5D1H4q5+GOh
OQJISPmpnhiZy35j0zVfX0F604cNLnYThrZcUxqMUePccT8QAA31hQrwOp6zIcMSIFDIE9nWSMrj
EbuASnqWrO5iMwy4FWbYV6DXNw4IOgG8M8Bmjpge2EH7XiPYtmXyOXuj65v5JZhmMGQXGm63tmId
duGJZk0T4EX2GU2hv1c603K/U5GhHhwbqFBWHJZIcIhGvudS26lsw4ddEWDyuxKl+jTI0ldlMCHm
eXZHdkQZuFuv0by4OHYcVGmyzaih75vLSEFL4HkcOkzIjs9OPETm2DDzN6/0kwUqfSiW1SbG61P9
Vmss1wM6bmlHZRoxN7GjoNRGwzn97XRpYkHmztMz69h4KWMYWMIKpvXZRJueBNyS2I406AgHLxW5
nPSINBzy6hsmwPOpYXlwAjQen43ofAwnC633P8R7e4osq8c/mEJqXPemeQjW/1cTuiWO+Ydm0AAe
lCY+urpti10lpUC+3i88pMNjsKRwhbVZXMyO1W0wrfk0/OBxM77DYtlyw4Z0xcZjqwCofNb7ccfF
geZj+1KaX12Y6mwzQR1tFqhq/KLOD1+D9zH7Oc8snKvO9lKTdcuw/5oVKxKxj7gw0HoCyj6+BLhn
bPByCswCvNgyvhSEIoMrp/JhvQT+/AYJBY0aqIZjLUUGeXOAgNzI1DZ2o5QtJ76R6uZ0qlpsdgTT
kcrgjyUagEDk0gJ0esUG+Jm62/i+4RgCyTSPS++/9JitKgN9oPT7t7J6x6EohOkzWMCKsmeuGL1f
ROEB75Z7TC3ZwhOfSlDDhB4F0CYzh5BqpM3hHcQzEPW32hfYAoxTeJGjYBgjabveCWaBg1s+sulV
dFaLJw2tFcKOsZ9UkqePOJfyEwEMGZ5lEaX9cZV+EF5YQbpUdBavSh8w0zN2STbHEdz6qmW2tlAi
ZVi9kcGcbcOY7SVrEiJCjBq83JI6oVB2mrCxukjaYus0X9Mx0G7QS1vKH+Vf4BomGaqgVbzip2Jp
8fGDhIwz4wqhqGiDL2qq7KBiwtepcv4VnLoU7y5N0tLV/M8SjQ6S7lY0Nv5JITdyCPLB/PNZ5I/R
rI3EZm35OVnifssF7i6+ROClP3MSNtPDYA5PrzdWJFHZuDLgW/aAhMjTZm5Fo18dlOj6cS7v/ABR
wIp9k1PFsbTFut1+19fCxXXypCsGlBmDIt7afgr1D49OCVkxZqxznURYLCXd3hgipeGO1zdRgZeK
ZXciurQ3O2i+zeeKpG4RAGzKykwICtVc2zwkenYScLn0k8vUnTBNV1KOttk3vt6vQj5MPTOCLJAg
ZR+c3RAqrMcMvcO84pnu/zVyTu3Gp2f1VdwtL4JNTKLxAbu6Khp3ZYACIVbxAuSnQU7f5+Iz+RTf
V9BeYeS27YqBEM7ER5XCfUMfLC+b4Qp2U8S2DtyNolf8T8Lqu/oWOFQp+UVXf29PJIe80t2ovUQV
agOlqyCp3cMJSW9XTHVbRUmyrrGQ0tefAwvqX4Y2nNQW/4wtyhZ/057V81wADH/Gd/hWkeq42tJ6
XiqYJH4U5JBeObJVZMZmtCBGd5KRuMV7v0/gae/QHExIEf+eAfdZXhcKMeZ635mlAOP/n0Tvo+iv
42vUbOp7opEBsl3wd2oISRpJ3iKBOFM2NL11WoEYogqyUZpn9cG1n8XCJC47Xz0xB1G7HlAiM3jk
VGzw/idDOslxmBnwnxMbW4cnJJRGk8FNRhP5gOgzbXrBvArIQdB/PPn9m5yQ0IMnEZU4FqFFJUjZ
VG8YSedNvDbPhZoz94UwiBc1j2ljUeYob7cY1SEzCQ2GxYt3u1lD4ONG9uU6KCYYhSqzoirBKUr+
WG6KjnMzhyv6Tm+inBmu268+kdH5vFo3D+dB9D8YZDyjD9vSkPx9vQIJWsOjTRazuOcJOIpytLw/
2FEtXWESkmhex/KDwx2D1jQSUVkED0s2VkFhLghwWV3TrdJdIIZqYLGla1SGfi0OCrbo0FA926uf
Pzhx0uhKrUESU5eX5Mi/JWNdOxv39bfpleW9H7SLhGlE65V7In4MQQAXojU2NXuzyWOq7PWRwCfU
lEOVKGrZko90McdwwPTd2xniv5O/kJQlG0ZBA0dTqG8VYB0fmgQiPapckpk74S6tUQlFteQ27BGo
Xnmx9vI0Bagl7I3hpVrIwwUFZEUZR7rX0VfnlEY4EIuWAW7FZuPRfJ+cE6ZorfVnxZD40XL3lM+r
jTVtphHorNOCg7U3/vSluS84TytVYoAkVBO8WwHEbDCSrMo0h/oYIoUl1IiFzbIJYfDjU4psDKRo
RUQS37BqzLUUyDnx0uEnpao6VmF/HgiTnkn8rjv2HQk0CF5YI/NmX1B/sT9wCZ58osfQYjNUTn1m
RReaZRZsSsltYAAdku5DWZ7PlUohoxE6JjsJ+pPxvAWixGfCTr5SQEJzIeBgPacrjt+ZtXwpFzL0
pI7mupYF70lSlGhWoyc4yg2ilmAsfpGWReKqs65cETZUJghAfmkd65OWLnCnFbeU5FueNNhzsVPm
7bMFH3C3e3rIC8+z9npT0Qm7beEnfTZgh8sSElctN5kPHfWAIlZu3KXuo/8slrYE18y+DHTocXEm
v+hl9RnKQqRi8AdWg/kXnsL9cb2HPhNHyWOtNWPe8SKvbEnlFCXeTU0qy6eRYxHv/XFQbE/pPmCw
QFQbFEuieyqyRPAmCDKwlLoOJy69wUeTMsYugvQMZd/1kr41NMLmWECrIg26HKmErTdJE6Afk/sv
pL7QAF5yLSTleVbd6D75Ekr6vCLRogoWDrJaFdM7y+wwRT1v2+mFJb6LyUKmjeL1aYFwT9yrmyyy
l/0GAV7Uy7WM298xagRwlkWa1v+qkxlxQuK2RG5EEpiKQLBRfvF7FXczq13Up+zSSE8Py9Pd6mLp
XTFQLv0HgDGGcT0gSJbi3HJzJqDO5P1EuQhCzSJf8D34DbRv/y2Kcfk5RG5t7x4V9THkQoXIDe8Y
XVJXdb1b9EtuhBhksj3BM2l570l+/tLfV15u8u75scA5jed8kf3TYKA42ECx2BRxTFTO4oED2LWL
VTEFQu68d/fslogryn0lOF1ZbvmyXtJEDDQcrH59nqie9nxwk3MzCmlRsLp17XpX/VWANArZmY05
fJBEP8M77s9YA1qu4XXyaDz+4iyDa6ApMszWVtQIhw6AgE06gcXxI29gJDupgkz/4Q6RQO01qGXq
f86hUtDaSeJFm75X6oWRpewnBZ0CVVK1xW7EExtJ0CJYUHVK8QqKk+gDtn26zvKkDx5BeNBHN/EQ
vBMn0n30aXlXqyOJMZ/BWoPfqRuXWo5C32ai65bKkfYTeBQZA+fTyDaajQbukwCVyBfSJu41Y+sM
ZXD1EtleO8O9Z1u1QpNBgmIa0DV1DO4xF8ARBI+fxEEKxRLjh4FczkxTlknTVpY2ZOkFhg5Au4KN
V0/TkexyDvTnFK+FBREIjZo/oGUKWdpWZWPf2/sKyrvbXatgUnm9yQFBg8TqZ1o8huM3b2376MvE
6xni++iYvfxkTsRXe8mVtjgurqWAHbEnpOOENFL/GI3lt4qbzVPaTi1dgo87nb79W9b2yhigZthh
5qt8bA9WDyaraRZVSrZQv8vJx4Gd/AQ2B4LQ51qc0sIypQ1DS17qkRSST5+GTfu8sQJMiDiLhadU
SD9GN/6ArsoWJpqw3fvHU8pNc37H+1gznsr1QsQdeXghOnsOrjtLfH4GdvD0rTOZ2SWRMln6vNUc
uOjm/sU++UYMOq4XDSpstAMnj64K9QUx0H64zoAEpRsj/oTOWGCmchzHJRCQ8GlX1pWkVrqSl3z5
z7Z0k4LA6DkbE0VFHJ1OaNwGv7yA0BVqPuE65/Iv2Tq1gDYatPFqYeeTEW1S1jWUTz2pP6L24VJk
TDDKzfSsC2/gDH3EVjabnquK4VuFtSmQN1MERZ1QcdJjB2UDRG11fK0+npSJNY/Znd+nKgFlarsF
8j7+egJ0264Mkm52kO1QTk9Q1fsvHWlmjaYD3Mfd5HUZLhf0ALoEE86IDjpvJmrvyhqufYf1sPEw
AtxIEncs0zedA8oZHVyfa5b+WQyq83VbXF/zFA+ntMr6ZJC+BbdD2FpyHDTPuIVa3H6olUXcdnYI
qzm8gsMaPeLVptpsnDVWM++SIU2jeovUAXKz5fJfSsc4ksoipCrRepNDUmfguYnYX/CY8WWlfYwy
v/Q1gHBNE0xDT3TdmzC5kDfa2tqIYBXVf7JAyjasI6D1uqOZorvy+a0TtrhOXtUpZEicaMY2fe4K
eDXRNjNpqhJF1/3man3fNC2NnTCI4wvFGGTDm924pCsQQmZHgeVosz3C/wskE3bjAkCm/RjQZGpv
weP43C6zVDPQBwRiCB1Vmt4o0yGl9MCYxNIxTpYfXuI0XbuuZlaJ3algIVao6LSDlKHa9DBLJjVL
Rzb7FrvuLxxoL5jYwBmHBd8nmWaeuooedrF7i5uQn3sKSrpe+oM7MISjjQcktxn62NO42MhY5q/y
jThqfOjhgqAQMqZ55MGw2hvhSpLECrhvL4e8RefKsqB6AA3WjifQXFx2ClcGHet5A+Zd1OBrddBM
hsOwJRr3CCinNwsfTjcHIwvP9atr+tW5aUgV+ajkEaEF8PL1Y+1oJkzPBnXobJ3AScwCeupzxtoc
XVPGly4j0d72mlkLqd2X6b040NIEaeChYCFDUIpXr4abfIL301n/OYFD3vl3TekqVp5KR4OQlMX4
rrRRe7lil0c1gWVok/L59CtMJy+gaDFWT6WhYKMEvkGwD3JTM2UYlG25BgKBoKqJhkJiYbQfF8kh
pgrH+sCGF7YeYVxhjNQHpMz0aRE0We2k+pcZK/dRU8rstmMR6rTg29BsrUGbMfjLkD7+o4/U16ZC
WexOKTVGAYWbNz+cs11n5LQVcKY7B4U2/PYe6/JLsLxUWgfQOLQjEwbuuwOBuUW2fcIjU95YarSI
38Yc5KVkMhRj4gfJ3OOjXY2J7HmdKyjSAVb53ac+8C1AfKajhrSrwX7l4nL0lj+C8FRUKMczECFj
C+obyVEx9ln6dWP/k9Reyjjo5lWV+wGWr7Jxa2KQq1m7P3Xc/d+iLct7djEZC0jPiYX3j282brWF
L1FAFtpN3mOEVLAucJHKwGjonlIfqPsvgcXG14FC3SKYt7uzDE3fkTKQEdN/jMxsIg7HHdfFaUqS
hh9E58k+EruQ894X+rqLrw26OXh0fpyeAxC0xSVcK7TNvq8b+HTYwRQoDoKVSWQ/aB+Cs6pfdLXR
r4DCInnBRh9WwsB5OrqcZJ8W/ZuwAAVz+NFUYXaHcDWzdp8tASYtanEvD9x48HzLowHPoDHZm2Iw
1rvaYuieHNFgfZOeT+tKsrhWejLCLNZh6eJFzR0Mk2AegNknv/sZ3Wyj8ho/2ec64cYXyQMWd8eo
bjaCdQru6/kZyUHOxP8kmgeNCruRtSYTzOwtzsj0ET/liJM+qcao9gfcGCB71iJEWzBdnRpQoWgz
nr6cZXhMniB5XYJ/3hfB3v8GigsgOxWlERil4+zmd7u92Os7DvNUus+Ou8qO/fxZ4Fa0kRmhlsil
IMRqHm9s+d2iae07iLiEh/LiCkIPDiM3DNqkwkB2PU9FbIK8j/ToeH/eg488bar5/DQVDK1cpRIa
ppqXqUsbQ/dB9zZ0zKNGempfT21Do8uCKPwzux7kSv9zTrlqn5ocbgO8YlzbqYTvCaUi82yEh8Lz
bvPaWGCzmTH+XuxkMIG9Ns2VrnWIJuDxXj7awwf8Ev61VG9iOtYyUtv1NVau0Z3jLrgUS2WhmKBv
YHwiV4oisBwNk1Wk3qHJXDIQmN6F6wL1Fc/jZMUCMWw/kMNWvrF2V+nAapRUHufmGdaQQq3znk5F
MYVcdsewoJQ3VnAvFU7HJEs0vTVSG3Vd3eGMbXNj2Lm8Q2stmQnlje0cEOKvb0+c1UHzUu32zVXt
/d43R7LvVtWWi+XodWBAlbFGr49HZ+t15ZUruGMaY/U+8MSIuR50tEHEdPxgtqjwgljVCiScJGxD
615zGTCBcRz5f2zXszZPYfDyG26aZnbN43SZQ3YHvKhCK1IclONA0K+flmHexn2K9LAxRklhyrV6
kZGbWcXXKMETzedG78VldEAC7mncnecTjsWnOpOEsan1eNU2svm6Td8j4AMLle2Ta7QvUT/ibL7/
lKHuYq8ueRkGjnXv4PFTc+KqXBLZpVv34sPvQ9HPw0c17Cn0wQbTvxaFp05/OF1eM8tu1OfcPVRn
xgvdrPsFZHfGEEMqM2okYsSJwKxaHkkoiOc5QL7vFDK3g3JnFQVuc8D9jdXQSIpOE6m5nXXXcjub
xp/KrbITUqek4pImdc47oC0RhxqhDdP94tTVAeiEll6pSnA5yrE0u+cqYIVf4PhL+UQD0+6FAeMl
yr36p4R1lQ/JAQwGnRbdBhhSs9Ni1XJYBGuKWBLxddaKls7yH9kyOFGkYbT3MNjy/ER79LJBMxgp
ddzUH6tQFsoggMPRWjnuktsf/1LHGZIbffUcwoqEWGvkpVsgibEvIA6h7hfi+HiJuY+TfCf+sh/3
lnux+r3soewEZBd+93jDDWFOLcadn89Cjs6HoC/b9pOFhiE7m/sHLLQXlSKuptmeO8DNLKFjzhUx
Q1tZRuE8vxOnIkMSC8KLEGWYyEfU6+x74pFzrIAwbifUjX/PH4HbgHUWMgsnWW4EjmvdFb9E1uaE
iokTFpBEh9ubSvpuvUkdcVr/SjUZY06SCcJb5EOi48rnoNxLLeeE7WXO/kNq0cXDjlOxRdt+dbEE
MnJE3lJvAXbMbYoGvNjXVpHcZVHG5fFzv2tm4TjIVd4GXmNIRTR7gxU+TIItTiavR5cHLJ0HAnQJ
9IKRpDFXD1I1Numj0+0wG0l+XLUXoR+RP6bTwCZBWxzETAMOwgjTiDrGG/aadbk2414kj5Vb1O4u
EA9tZC3/VjMeytTCmoR4fxoVPd/j1mlb1DzjOToeKfbOjlzLFe6V4Jpqnqh+hCYchN/bhj7nOe1O
sxsBxv253W8z1+JIIh/YF3xw6jLNFt8gC9rFfGrIhvbOLE/mMFVtcGJXgVmif3pydflkamIrc2p6
BCRVrKsX98kXmyzYkH0VH9B/arWIiPMZMrUyfxEAPO7C+BNxojKC/Jf6ULM1G4GA4h5IddhiRl4E
YS8ix9ZgsR3ugZJ6kM8oP+LOmn3RoPBqsxkMHKYeTBZhrm/GqG8kOd55l17JeGSUIDj165qk7JXP
yMjXYtvZTmhgwzDkr71xAc0dQxq5Gwp1IEVTln5YJlh6L7WMvWszXGp5Kcv7BxKZCk18oG4qf0Ll
zBINIu5OD0KLIPBzOteSvK0uL+YAR9mdR/syxJkDpIco/ZiP44bp4JOUFG4LNerz5L1mMBl3nDG0
aoYT+5uEGBgEXp04Ir27jIShL4LOr0MRdL63NNTDKUlslpl3/pMyg6YO3qTQJntAgvzcI29ZjDLS
VIMIGejr55ujlCj9Hq//exZ6FPE1/ADOdHPNMk5MaUMcVBSo2LFZG71M2/CxeHLw2/XkjJtAHrOU
tiswfpG1P+IkLGEbd5N+OHKix/2Ub8mBVmXtbZCb3EztHJwtos/E+dqzhx9iYuINlMKSZ8darEih
WDKcM9wQ4zpwmo6pYsfpUEcNl72AEPMDJPNdCbYmQtEqvMRLJmxE+SEBbLIuslR4QAfHeU8M1PA3
Ic44NworuK1WnVQogJwWKrJovyQuz7mVt8i6mqvsW0YM+85a2Rk0OojYDZppf9C6b6fwp+kO5WrW
/AaYv4ITM5QdLOJKs5f6KeM4eHAm4KMtS4iYjUL9CT7jJtXW2WiZVa8alRLEx38Tk+0WIQMgDeIT
MYGm/tu0Be+0fQg+1Rmw4ymbkWuGKxlIQjK0Lk7k9at4jIo3c11lqkg0UMBsd57kgfoh6+aQfW15
Hn0Low2e7YMNF1oy0tdJE+qCnXYOvcYQo28hLhULIj7kt25aXeRHlnrekBHiPLULphnFBZGUED3D
jYiSUGZdjuR4ge1v8IOwyJay70VyOcn5YE52ciZRFJxxvojZZ29zJHd6mlVesAs2l9lYUP4OSnIt
tKBfy+zeXRQvO+ryrGuYyf9MkqCx/3m892k7EE+kzf0qzbNdRPY+8pNfEueGGovJ5CqQfgzNyj1O
u2pPBBfOkjmctK4CkUtrQWEiLR+Vud+TNiEbqlMdVoPN2ADJ/+NUPo7uSq7WgADu0ZcNvNacPDd0
S9G03DRjCouDfnmJAyWBiO2xwLe3XqOygA6V2vUqXmBxGw7Nchzg4yX15T/0a//fqeyJypOiEXzw
lbocmmEhsKuD3gnXbJZMCdq0pWyFMwwFLC5Ht1Ituq2kyRff9E9SRZ1aiSyJv19YP9SFPl5q8eY0
PTVxA6FsM1d+kiaDEDn/HLHlkUzAOnbGV4T4IUba7Jn9zIk0o5QhjX8IB5d4OY8t33ANUEIOumyc
blDawea8+LWGE6N1hRfDD1vIWcHM385PocUGjWrTMHZUtOSyAdfoyF9OEhJjVZA8Ajqar8SvHPWW
y7UUSaZ9ZD8EsR/o0xD52CGkjfW8lwwRKZInlQGMH6BJzwUGMay+h5LdW5z8UKZYtiupxfo5ykO7
suG3f8IBzc/mC7I50o0gNDLoJxpqQVlKJk7W5djDp2a4hn7mqv5QUQ+Wn2sgZ+qaoKl+eaVN93Cl
i4KZuEfkOrh6SQbaJydLL+Arvub4BScG8LR87eyDHrBcfZ9WGrNEKk/J7pe9frSKuAFhKJy9Bzju
fWAil0t1z48zKmDA8g442sD6XLPyNzlB8tBV6LmXx2CPiMV6/GPs2OahLEKwwOuu7n1bkDCS/aiL
2OxizGpgUPAtQ1Vfxu0PHrkHiuMAGWOxfdbeVjhjyoxDu/Mi1ye6A7cJyAB1L5AJKiqiuQizxWTw
Elt+hIe1pTyQzzxZizXNIPa5w71LoW9O/ct3QKMNFjsc+rXsvtw4Dk6que3nWAPrLrtbWpdKXuxm
NSi0I29zK90E1Seg9Jv3beb0kiWl+6CcqzLVypVZN4G/1eAmtPBZMoLxOwzqBr2lfgWBJctgDbjw
uiIl4g+NVp7FwwAVwWoHDb4yOak6D5acWA1u3oo12vdV/Ml5i5eb5P2B4n5tZ88kF/PvxzCLvML2
9+nptKTuMYeLWomqUkiqLvacELKZqLTU1XTKCk4zwRPb1VA/tmkPSM/x0lDapvZk9Y7eh7kCLPJB
stJ4p6CIU7QW4Jj1630ERjptPSpBeQKuUoudvTnMdwPVbe2jspad1NTOx2zJXZ7vzp1owARBswEb
XJ2eJPRV5J2a2TthxeKrdwZ6NghNVhp6dJ688K9k2ieNHO4ceBemdt6tCZDrZH0rsZj5899+DBFu
j4j2y7h+xtt8FEmxr9KlDC9sA9BHzH4UwgwMaupKO2YdjB3i3sknRoOM186P5vCxI/IQz68Q8hQH
5KjjRAevjDlH8iRgxVVbsydgLh1MV4jaVtU2IzunMPL0zh47BtxknBtdsUwYFxc9+vLYyyYmhYJ/
8sdHAznhbr4UKDKoLInCkWVokc2JZxib6iYmEsEkInUCFnzmYlLugkKbLVa75z6ZnY0ylWLqfp9V
excNOPp8LPxrVa5KZA87h3mklvmZYq7ArkVNXv4+cygXhqZgb08r516FUljq76YMTYciyiVW45G3
iOSnu8BhCNpzGL7EyK4wr4G8nobN6Cvb0Z8b6gy83wCS7xpTVCzNmTsCL2PXKNZ6+CkaOFIgLyF9
ZPWoxPsIPAGJv6x5G4KFXGqwkZy51fCsjmJNvvFSDIm4sS8oU4rYjN9mYIY1TLnGsQjowi5npnlV
1X2MdLzoEg+1Nx2nnjEPK4Uh0mu3rusnSn0vzj13sCqdRHiqiGvLdzZfZL+Pj2ImPJD2OxPSmN3W
ERRniOVMb1eB4YO2uG0r7L/XuMabCTl9f0iaXqHAMmU+O9LBdT+ozOH2ifLLrXvMThQvIWPBqbnw
pjOPRJck5eh0XTwZ549qtmccsb/o3kk+wb7ZDG20nzLVaCGhvIgrkPTSo0mdFe9pPbpRMla6P86f
SNI4JWok7CUGNTgiqYim3wuNml9KCYDRYTd6yR+ga5EmlxyJXtDZiAz1DlGSgCJCkjJ/NVXHlsr5
f/KhcaDYb7y+2Sbxjg8zsxkRkbNkU7T3rnoIQMfTSUdKg+yHWLF78ObfQZE7/pQZKlZ1bXJ8NApG
UjIkn7eAi8Ep6ntmnKWF5ddw5dfzKLYL8W0T0gyg8qrUrE61DQGUdemtmCkYAApsnWgzias9xaXl
DemmkWpDSHhdJaiqfd17Wb1adja+rM2BIpZBsl8XQdsL0rH+zZGSrvyOL5JDCyvMIyjHr8aD7tnc
lsykbq0Q81NriuNDe2cCTAlxBWgo0h7CKkgaHj9LtOTKWA7/2f1yvXk7YZpb3x5sde57LPgZNofv
aOY7baT3I9u6z5LozPn+3BZHi7AHP950k+BlF3flYS8YX0B1MGc2dDz+iUB7VPsL1nknZeBC0avI
QZ16bV6kD5pNVSqtUn51slGsJkCxNHE5OrBUafHJvkX6fHl0tE/2bIsyEhefMluMVfiKqTeAcwNB
clQ77cnQ/G3Z7H0x83xA2AkTPCUKhTjmrXmZ+IPUz37cZlotyXLrC89LfJTnD8kL0T3Rgzv+Jglq
bLUbX6NSpDpcIX1lxfF19OMzNic8LBo9i9YO3MrlW3a91c7B+PauPbermUuY1moq9OaJaj+Doqs7
E/KwVlzcb4qhKtpFwNFm0cYTAKrxTpeUZM81ZHFCjxBTwaGx5YIt55zDUOhejnkTQlUXYF6waeHU
DW7fhPrljO9wUk+qNp7K8q/sEKXgICMUbdmp46ocKdXbp1cAkWU7NSxKCNOYACxPLXWQWPpvVir+
NqVtNghe2wlbnhN5hL0AQ8FrFi4f8aIjhXSjRmzVW5Ak9ZK0THDNBAt43prsHSS3ccg2VIb0Ewkg
Y6Zi/Re36+o0kimOWL/ok6bNtaFI2oblbQSzuMHTXqzKrRqMQoGR7UheODSVWHMXO7rYZzUZzKgJ
JY+jKz3xkqk8Mk6W0ait4Ebun7rAlHC97uwU58LQvXYRzl+JzLNLcxRPZUL37hCcwy+Xk3dBIiPt
xsk1u/6Ob6CxsIkS6IbpBbmQPlTk+fnsLDMhDIkxvTlHm3E/cGKYOnczg+yhSXBLLL71u1EQbs8e
1aotUrl7X+BXtoMP+VQnHVp5Syll2pH0pr3mOvRaPXx9in6jMlm96m6VqfnFKiDG9vgLK3yoTTuL
F6mjXloj+jrDLxAQK0Esj3l7/zuHkQtrCDm1OD3jIsq6JT23L28XOgzaiIrnXK0Jfb8E7EqPk/Ht
Hsdr/yzFOFE1eDFVc75Hy8ebp7jLfr9PsY4IoA8nUNmjvmLEjILd79H3n0XHiIzauFYXY2INn43N
GFGviC4+0kLQFAVQ3c8VPHI+pk5onNVC068zE4MH5rSO9KDBT12WOF3qaezNMaeNY5yzzgVZm7ak
7k+5pIKPf8OA5nGEWaQX9zJKrjQ8yVqMCJM3cxGM8FFqJU0hyUuiCqNCGRPkGWeyEtRUPN4Je5Jp
SOxWoRbaZ7oKMtcZj6Dv/7ivtKc0SjdVdvU9lB+PYR9Opy6c+YyHeb19HUf9OgxiTj7UrC95uhE+
rjxDKkn7Z32EE1tXQG2tEpbOxa+4UgOGcFVVDNqfPeDkDQCEZHFu8r3nqZBYzdEfGWGV4j8yy1ST
vkc6FKNLIekndIf1esKmjp1vd0tgvL8HS7bMrsjbPDJGO3hcfsd5DK+dnqv+6ZJmRjz7olQWIEE3
ry4nZSlrtf/M9Rc/JSNkDKo2xN7fPJm+YNdMHn6N4P9WkmE9G7FRLwfPd8Kfigq8xmZPJvdQ9LxJ
BZ3eKkQlkIORwY4ZaDLotpybLhQZyQg9aY0bBNlBwK3IRWag7O3qeFJ+mLsOZGsKj9SAQFQqmHO9
dYwtT8ZR6seemDjEmZqF5VfNaU0k/WCG9VYXBZ5JNrGYPQL8PbYQT0Gpb5WHJe+vxarhPQ6S1oQw
3FJ3eijKEkSe0Mn8shxTmd+qYetIBf5lhyXJd9zZaW6HW71TRiL6BdO0f6kb1Iw+GgUl3x+5jEEI
RcLQnV3Tx0u/RY0H5df1ARjF5P1ErzdOi/aTZBWrbQEDgEIC9NTSmqBEVTewk6NqE7CBuuKQNCL7
YSDJxvKgGt2EYstLYtmkmhw6M/aBABiBEpKhqleX0yW5i2wrKmvRmppMucwwmW9vINhJYoC9FkA5
nR+P/Fd8iCF1+uXR17+v7BATSNvT/kAsAsLBqSGp1MwDDOVludVvPxdfMdLxTGJM0JbrrclapaDB
k5pn3VzR0rpR7k4GrvW31V/oxYL4vLYHy1WjIMCYS7J9vvyUxFbCw82Q3HHI+1eM8IjwXVcgSX7z
axKeri7ijMjjW8b8eVmZqBzWf31nwyI1AWUkOL2hu5a+6uOEKOBq2iULNbxr8tdd/7k0bYOwMwdr
Jd21DRytMqMLUd7NXhELOwOIuWwkZg4oJtq5F9vWPmjEeysY1MNMOWQ00zxPJzOOFGRSGbfqjc8G
0I+sx3O949dWH3/A6o7VXFcpDKQNXKu1R+jxNGNjM22elq0Eky+IURJyuEtc57VUKUc6LJEQThQm
XHr5kpkw2+AdSrzg0oLVtsDy0Dqc+/xaF/mVbfjL182A2gJP8B0S+Z/vACYpC8Vw9NL1jTKRwTMz
LOTU8wU8ni6E96SEJgSrqwBizMfDfggnUPg5d/t1l02GiZ+QFhbW80fds5IHbhl5sZ9ieepcOj7I
jraJnTxNdQ2B8E7jKGOUxL1sCpJjJOAIOT0YI/z1fBhIGW5d0OVClCSx+5lSOIMOiUZsARUgXqKx
6oyDG5T6L9FsfRa/s/E2uw68q/m46Rk0T7QjChrH6dgZoXHeZEfaV0iQALbp1VRQ89Z93L3L8tA2
0gkckW3qHAH8z1t+G1mOon1LxrIwVpodMjG7ChOBLXU99b7j9Osfz+dxb5roZnsOOqDkKn2mGwiR
pw126yJWONnXhmHlw1lUr5WnYWRE35xgU6Zc1UVh/xKn6ntS+8rK32akaeV+c7s64w/XIwrZNdUn
N35Kpuu1I2q91nQoizfPAZ3uH3aifj7LIspC3cxe/nmCyrfshBe9xf/LKLw96Xo+KdjDX2vVLYhu
vRPbwEZHfrC4zvTRy0E+khs/tVG8tbscE67zqx+YfO0V6qV47xgH1Jax2DPRnU7AGxfIj402nAFI
uev8aSBpIAwgtaj9EsIxpnmuhvr05tMnOie9+AnT0zkYG9tpHCvyRKwRvXA8oa05+MR//NNcPOzf
i0131p+JiszBIX8ubBpT+bZzMnz+YR9zIJHFNSIt43zTFlwcQI2dpIK1NcivYUQbh+quodQydcgU
CHVgtuIoG149DWnsQb8STlRInMX6IxCyDlcpobjDWFhFskXiqv+lALbHiIF2XjsZRn+YH2qf8poF
H9D67fkQMHg5hMzOOcEVCiwPFQDMxNCRZ9MqsWR/ATd/52JWNKoHmAndt/aEXvsO+dju4RGFNW/T
6x8uGkqIcrX+vnFGGmy189UIEXeD7cNS08JD2jTEvmF7iGIiyF+J6B6pwn68DHByVUrSwLGgo0Zx
ACjHRMew4/wJq2GVCuTqBBA+7EvTEAIuMeTS04rWloRiI/fIg3E86FcuvapnSPcv0vyFZAUadkGX
ucfm0XXsytpVCSfavq5NXzNI0smpZmrqYIM0uRxSOIK8JKkBCbNMwje33F1csC1X/11BSqjDXYPL
kdd4FC3FjdA7kv/pemsGBAq7w5YFC03ibZcVM8PZ/F8PuGWHmcj42YZRG5upE0snx2Ikg0d/UVWG
cPTTn3h/g0lC37Jmc7NSyWiZRgxlAp1Gy9Y9mM/7eQnGzTPm7WCG/R+K8vc+1Szl3HadBLy3vucR
l3hb1yXE8r5IhPwdxXNBQ/NCtGSpB16jFJ5hQ18n3prr1ND/ohXG3/fXNmIAApmWNjvbhQwh0yYh
m4LvFWnAKBX8EbweTgoFO65xsKUiib49StjLhppFptunjk2mH8MWAvkHeRt8Emm1Gkey9NWLL7gs
TabguKWM9VFTPBLkWyg9bWXxXH851cOz3hd3BM0a31IgG4KSSzL7aZEeKXowvAxkcY3MBPPDXCsP
RUO/ix2FD+zfS198tiDE0NSvcWKC7W+GCY+0YTmuzAFB1XqfRFf8M4siEV+3wnQP1s/TH6lIxCM1
TIw4RNkH4c3+7wAb7TG1WWnC5TLR69XCr1eft7c9695CGQr6nPX8asL/86FL2qi6A9L+ExXYO5SS
7WL9agYGnfpt2mt5SVgptLwn2hdkvNfMOpfE2vgNAC6SKTwU/Mv8GwOhr32WG4zxBe37clLSXluq
qGJ34wCTWHgycaNK8qZYqpFjFkjX/yj8GhXBSz1GmMXIhDbjaT7mJAHLISbv4W6covjCjsGU9zoR
Hcwln83q//6h9eMb7dkVLQjBjq37Ndj22hCVo4zKQKr/J8TUlTScrD145vkfFHYngmMUeOMKCbCG
qdzKbI9RWD2jFpUJLG//2uo/nozkPiaFmHnZE80RRTOdR++5qFBN8S1PuovJkCw6SRmwytn77O2n
Dz5EyTFWDna64hPBuxnDJeNF5d3w4j224Qd8j2m7A6G+Vh2bMN8P4NfnAUdXlNLCH/0ZGQXDPhsl
VFgNiPWvx9lckGaCTZo6dv7/Xmhua8wF6dfvp/jdy1rt7Z3sC5D10cJIJGL/0Ss//tP5/c790KBk
6JsG8QQvMHidz39P1URCxydVbGMRuZquz+h55lyXKGfTiiLpeSuJLu3CpiqkW7VtmYGfNq/fL0dX
cZrZ9qw8/6BwETrK/JfBLendNrdX+Yw8le28ldXs3ndGUz1zq7R3D5Bl/Xx9xXYsN70qzfYVy5KK
/wn1OoxFsHzSA0flpAxxI/+CXdDUO3O5e/safwfRnF1ezZpUDNFiEszZhx3x5nIPd8DgSKDTu0NG
xnhdCQI1S8WE5fGnQz5pP60Rq0dL2RmTK/t+TSPUglqMv3ccAhQtj5/ZWMgnt5po9LSTiZvibGp9
6lkTbxHze190ApR6P9u6mjggZGrxUGYrJ1j8eGaBBUmhNTzrK4Oj0i68vbymN83on7hvzhAU2jQ1
QX1VUx9+Am4VC81G+4Z0+Q3irHYhKUmZRXZSBCXnzgmQwyKa+ChXLVFNNKCpGqIBuQGfDYsJcYik
gkmqMWqFvnsVtbbjWDyJa+gzcBIu+t+/jA1Zt7X4knT17gHrFxAMfr/zD9Niz3FG6ytmAZydgF11
h+xNRsWARgogN3mnANiS0+NV/XrKoqQesGgKNitFuTholaICgMxUE7fAEOzsTPv0zEJM2l+5lNJz
TcLg8rhFquIjhUi9wZ/7mjh4CJ7yVh9HXf27xqzeDHPM5QPjT2sebRmTNKfWJt6uItA4Z5VKmPCd
MmwRcqyqDVEUqlRGv5nCJ3uty6eIULwpUcY9I/xYQ7hdvaguCT3irSExIj9j/H48+uRM5RHdbo0F
2bnuBN2GCSf0UK3UciaF0nhYTAXyP4UVCh+pBy8L1S+mknJHBvl2lWA8exwVRoIKmKwLmV89S9DN
A2xndoqdShCg4nMJEVxvTZIZscpqUkw3e4dWR2s4c0dCEEQ0fqKs4kjAfdtc2rHvWCsa9obg1qWe
ZcxqUh9oJc1lrOYNa98Ip0aFUYrwlT+bIM28kiFlmQ9HXLeiFw2xrnNgNjuTBH5PqH67XXj/P3v9
0rVjwL3J9iHHlRODc3KSNF15pjXUF7Fru8z2LF49zaRnu1jk8sBDOETZzgVt4bnwH2vGRo485qAF
klQrr3BpQFubvkFsL3dazGOVtuWtxMP6LD1NhccCvQh74bAc9GV9QL70s88E6JpydH/Xfwl/8kcx
577h/jgMWwdW120VdV5luFT5L2DcPZ8AgiWQuQ3R2wCf4WYMAmY610mOqnfhIHqMSFlGvXZKvPms
UtK1mo7fNBwamgeXeZBr0VdmxEjOMmZ91XwfpGB4YRq6QQGYX2y5htk3V2zdHbZ1vCRqF3p/aZix
FuHQfMDTMnZ/CixZagyJ4RvDIV6uHHO4rjn2NAZH3QMF1ftk7KvWcH1ychlPw806J3m07AFl4grz
e7rYFSl3W8mKu2scTDIZBQ37lQOTkrNF0pp/Xj5ux/D51MF/tHBAug/rnqNvvEVBP5koXYkmTLtG
fCoICO39ZTXEhGeT/qk6YZXwRVDA5n7HKal1kCT6Pt+DvuOObzg6b+9s2txgNbvGePIEEzrUBKNx
twmel7C9DC+a60SvEXJ8J5WVnHyrmhNJEWjJgiody6WazWZK7GKwH9t+k9H+JWpdqupGMRhCMNVa
on4lwjNY5ZdooKld1zeM/7cEGbesBIiiYv+J0ZK9dxY4nRW4oN3Xssw+eu/QC5mptGGUGhohqyNf
/CIN+5Ny/WQ7s38NMa16grhmEJ7W7MUg7zuJpm338wv+UIMzlODSF96byZ3a/C3yXGZ6UsJSfDW1
4WNqBVF/PtoFjd9Lk8yemWkBMp6nc1QCId7LaU90bvPvVZm6DYCXE2LwrjaTSjCDgmzJPeKTnzyN
pT6/bfEGasc+39zSP0oZUOj6JrfGmHUgIE9+2JGvP4z4R+pzbAgnAzTDQbCMFQMejcddxZ+R759e
xiv0ne+HmHaaHILk0Ek0phza8THLUlHqFsFNsRLxoWWSIAp2Ewnj3ENq1HE9QFhleUvhFy9ssjiP
VxxunNyP9lEqSeauac2fNXGUKIGGp3vwykdB/vNvC7J1nGRCsTpeDhKzKbgAk+5EvW/QE6c7mgne
gkFB9XqzU777oxlyoLVL8WV4runeiK1a9SEnkmGAHsfjg8Sybgnfc/pySrPDXWku6oYvwGUcncm8
yYJ9Wt5CK81yjOTtUr8DydI7w3CdwOSu92j8DqnbsbNEikVky3LNl1dQ2Vuf6YRV92a11p02lQ+P
8SFgtRj801VLUVW4X0+MMay4P8O8uprhWCjg2YyWGMhVa6c2lgb/pvpx30zIC2NWFBcgvGXN6pD+
xZBZioCGg0Is+sZYs6eYpuph3EZBgoI/dXc4kHrtxh0OijSsOlUcS0plPb8/B51VPqIuwW+u8YWg
1Q3oPhTrFnIoM5ZwC051bMp5aI/fcglim+ow0L8XyJEa61blf2DqP224DuZweTkwLr3PiZ4urQld
VIU6n1Faem9vWQbdn/VXWnuF6HRXQp3ghDkFUpXo3Rza/KnmjDXrt6FCRpRDZgWFuioB0hoZ1QQA
NTh4FEwok6FB55st0YesJJIRwBrdDjpJCtbhIAJKUGv8wSmqmECnG4BJ/HWl4YSRhsyqw6f+14nN
uVZl1fGqOHaqp4S7AJtR/2N92PzHjpBF04A4WApLE3RbeLqe/r3i9z6vbIGo8sXzzbhh+rZdM85n
epR3VNenrF6nb2bhfN83CHVq+tvaORFLyRnKwW49STWRu1e5ycfnxoctljwSNX4UaN68tFeTO/dy
Zmlxj0UW2P7XrLRbHFXdMy+gb8ZoGr07ZYXsmKQx7l6BNShEZl7nLcUld51BvrYukaDS31EogbqH
3973w/w8EujTpKorIBD9Zem4KTAQCwStwAjSOZhD93+YWhj2/r2Hox24fm43+Xgrw4+tx5+gGQPN
yrMaVAni0ahnCWzVI2yKU8oEc86lW2e8O9a6kNz4nRYA17QoND1NrLTpOWShh+3uZ3iW/nist767
Nu946kv0L044hoBzO9wfqypzAvN8cK2kqck98PjUayT0uQUL2dO1FnDu9rw9vMD7tFLpPvDV2LtX
1i7fGOuRVZhtiatjE49TrMGAoSmc5Qaz0ADGNJti+aPPHoM18fnh7Bs9uAXLFrJmbpL+dB00S1Nq
wObaRP3d80XJ+vU2/GtICcmUVIm6vIZEz5+46lTuKw2jVnKxdFO6b5CfZbUlWOBz+jvoGNJ2iSks
FCdukIJQRFHU/gte9aHSsGSiNpGqRBP13lsN5gywwZMrkPzQwQE15AZ9sNHtCYpp+wy2oexlo/0d
vljFzaYnxgxy59BX2s2Hw9QWjQ63FqY/LW2cI/cr5hdHYE0GjyMglZytz1yAtzoiWw8N4dqcIaqU
Sc95qBoh3VkfLwx7/GvcnMYovGhNTs69lefzVMYTV2frqclKKQRWuznoWHyxjxbTuB8N9roQcUxp
XNUDcGRX3oFRMC90hLnq4PcE0FlUZArCYrt2h/0teuuWOveYJz2M0FetJB/7M0w4SXslJLpBw1cF
/efV1da2GPfgwvw7PIqp/dGwLa2egexbth7GBZ50V0Pla1pgDHKFEbb/XNy3Yue8XZF+YIiQ+K1N
0zRy/tW0ZxbFrrmXjVrStBasn7gOpU9bAT6da+OdXSEqK5JddFtJJWyQpIpvBdh2dNuUCHMY6FgH
DunudCjl25JZ1VBVJODkPvsxBuEiuZ1kGt3KjqqcPMD0RncGdN1hYe07MeDDh1QWOlgafhU5YRrZ
mCbWJHKgFlMNGnfZbk6YlSBe3xgfJIURzxlTR41OAOCPMqrjuELrCmofVTztmnMLjjY9dOhqUpsH
9xpsarGA+37t6iDI1qo+W1rSkpVKnkjkL8iF4Y2b8mDJ9U6lfVvWxbsv12J7cVJO4OYz2OkZj8Eg
98NmM+NgDQx/X9l93zy5SOSFS+psbo90gi4JvqiACXIC2sQvCDdYPreWwZniSn6xggVC7042rp8W
dd+nQCRsLejwNHBC1WryRPLPalvPFzoIHfOofj20JnGQPSeXGW4HavSdMgSp963Oe0NbCCFHaVom
sUTPH76YTGzYQsm32cXvXWqDaNdeKdr3RDy8XmA7civG+8IebYuhuGzQDguUivRl3YrG4DhYCadU
sv0EF+vNRHbQrRXlMVjEbis6VtqSPc/uDyNAFFl3vYRgPkNQCOaWp5t1+e9iyvp/F0umzQbfxE72
EQzoo1VS2e9Fdtm7SBFFoKYgSSQzzLMXjUqQuwsQEB/hfalZrRBChPTQfZ3moVOSYsxrVNMDWj4B
O+8tZ0ALWKS7X8gwuCgvliH1+4hQgXHHCWJpGLEJO5UI0g1rtFKssBJMEZ2J1iJ0+gGS8IlGltuA
DPSxJqSlumz7/hXl8JICFKXXlmKBhH5n8Y0k9eRg5sG2r6XObBkDQ8zCfutb0m7ZWdD46sqp+Yur
psjdD37gqfJkbteQWecX0kVvkhIUagaRvgOcncF2heuWWCAvKMI2bi0pjAy0bNTNdyopg4EpVWxh
DmCBZb10aIebfmUQSU/rpHOyG6ANtqGHQEo4Z/dJr3j2f3Fas1eaII46B/TRs/E00BxPXk8d2L1K
wc7K2d26+DX/5jYdF/XOFhZMwyYLs7bWSYiQCPc/bG3yCT8kTr90yDL/L9Hu+0VZIdN44ICDiTml
oUTZTl4m7niXBXTILjv5E43UmZN+Mo4yBkRqYjjsQK67HIQfpByWomCeg3BfW8JjUuaPQsqCuKKx
thbAB8ix139TM1kfS366OYB3O0Jn1T9qd/aWHKTVSpnObJHLpobF+ybVLwte4hmK2W807QXtxAjm
/8JGeWhamSKRtdUBSC+UaA7SQ857ISkpKF7DhqeKM/6LvirTzsxWC01FIlXj+ABIhihjk2+zmEFn
4vlhc96rXFGNEZT+kJ8YSHfidIS3BqQFragNMZZ0PteR0jpPJniq9dKkyCiBWMIYGurHSH2hkbzo
mr+tYT2JwO+9TeO5jTZsa7tFcO+EXuXkK4Qie7XdtFDYFa5hIdlx8l/W1z8jGhPhaCyG8jzRdVGZ
js6DAUdzkETtOijhMZbVFPO+31MTD1vfftr+eHJVpmU6mwXvpjUkdZ6KVYklgV2PJrw/1cYLz4XQ
tWlwUXv7AGoC6lWH+oI48jPOWExvXpfYR/J7zaUK9KWHwzLC/BZnNHiWuGlCsEPPn0mpTqM5CeAu
hpwHoDXfdVRPtZp6+7BMzx3l96yBpThM/kGQCKRUSr+oYurctZor3q7G0830vDXIUyqON+XFiobi
GZ8cCYud81wGUWbBwbIQ7SIPRN16VDBbgDjl2rYgHMZHNK2MxNpBg4I6Dm6azKE1u2Q6Xv0q5z6w
ABnpTSX1VKbs3ZFqvZWjaBznildhRVJgT+YHQ01ZtAJnZnMI0o6ZYQUhVbWdv2MejiUvJJoZApXZ
qXU62mZ+KocgqIFdBZMvYi7bdK5Z3EidsYEFpl0c8oN+cgV0LZybbgH4l3pVjY7xvwugi+bzTwpm
GiBSAEBLW9mv5XedW1ZwfKaWpAPzounKC0D2FDtF+Z7badRC2mSV48Msz6AWtiZEwMVTUZhhEBkZ
zCBrLimMML29odwWkIu+etrqYiAPb0TGkBWIELi8LQlx6iRjYugIlJJMkUu3EeD+XXcTSxRsclW7
eQbrP4kbEV4BkWOyWq8oeDIxLDkBEG02e4DtZX2zugutHx5/JlMzb6vG6NZE0+W//TOb2f6EtG8N
5TcjfPqnm+Eadam10A6TIbfw4Z4tVgtEDh1DWrgfxSfMDLUEBjpxHet1PBisNlK3081n8O+NFwfr
F6JgxTdEj3yv+H1/RAhTBMBJMCDqDtorbnvctjRWlTOk7sdFuOH/uxVeU+I2XLBAW/9pNGjmLvlX
GRzLzVWT0ZWIvS7Momjc5QRlhMUvMrRFjvoEHoWEOp3M4FCZZYKHRfiugRE5l5XYAmWYrfq3JWIV
9FlINQNqtOJ9t7Zp5PZhCBzg/FYhyuRtWjz4wCCoIbBPDFta9OgNlqSavc5Oy4o+jgZYQHBh1uvO
7YvU3hJqBb5QOFY7bckYVqtwJwe1rfVCXzfdxFb9hkl2LadrqpUEhNtNz/shpQPmuLpgP4C15Iml
gwF6MS/gmeNvY6vX9vqOYgMr3q0tmHVAq62fc6MlXH171CdRqPFAw+F/jD8ERDqMg5iQIi+X83dP
jRuqjeipHHXeU02C3cfilbG5nzfyKF6HUgJ7YPCh3Ad0cs34y8I/8m3ZAwPwxPsf4snlxW+5KfS5
CxJ0m445LtXl8etoIGxBy1+qQM5iOI7ZKNgVUK0n0hTuZjSaoJP2bFOiQvza7DI5uVPe6Y5QvwGM
mSbYhLrlQzj38A9H8x0QE+U74/4+g4gowzhDWNOCsujQii456t7+ELfczNZSLl+Ey/M5k1XPcuML
al9pcZrASwJnecWOLr4OpS6qLpbzvLygUA8rLISF0N3yietga5zriLphX2GPksD7wj1Q81mwDI1L
qJt26yz50YSf1seh/tEegPCYpwGvo+SagIWbbn/WPNbZ/4eJ3wWozsbnCDLxRcSIzSnJsUxH9PA9
U1ojHso3juTEvfDMKGH3ZlmFoAQTYKEJSJgA/7J66bNLGyGa/MalGBto45JXVa2VvWYt313Svlgc
VGvIJ1hEJp9YsYEkwTQcPX0y90ZuN3CLcW8RBGnn3sAxvjW9WqGdof+RTIukED/KT5Mc6MyLH5QO
4siz+7SZj7cLelwnTs613gVekjgSx8rtPmxNSqrK3NYC1IYVc6xJ7OrCRTZZdgtz3vwTyQWRUiD5
ZpxM80Rnx8ivDbncsGQ1nQBfftFStU0+bMTuNs9qkvClqHJMqvp746aWsk9RwBZYcDlrQeQFpiDw
9pldbNr5dOjaYTwDV+3U18Y9C+pR6K+/l8Lf5r9oZIhyImIGBYiwdAWmjGmwyLvyfDd0d33ThjQ4
PwM6ag4TS6nY9b+bD+2d5I0qNyEEA49o+W9h3udovyGJdgdNQOexhK+bGBo7kqpljohl2p2iOAsO
19ExNepDowX5WnAknXVHFN193xbhdJlJdLqow0ODu6HYqHYjZ5LgqGyH3E/ek2yyQFhIsu0b7Kev
154qivIeIrqh3DHReEPa9qBZwzQyhOxTgzihoxKGPLzIA+Cfe7Xf+BV5NaBY4p0+LNc0A4oKGMrt
rz5h6q9KDa8bjWh5SVBUKJcPpkW7TK7XY8HJs1k2wchC0DWFu17ZcWaTyo/wKAI5n7Q4G1giMXB5
ajtBbTEd6uZb+3kDb0RoNxbofx/+6YsG6DPAEWwXqmuASnZ9KAzfxliBKjH+/kWG5GAebiRfTxZL
X/2wM9LNv6Fxud995ho+cmiGXNfXAw1hOsTNnarXfLjveTW43Z+KYF8vF0Z+Fx+Ig05OnZkQQcmb
aj88uy4GpfgfcXPJ7IUNZQkZIB5TW7fYlgDjBtigFSy2TXVdNFUpdaXUPBgJj/VK1LXtXRYdFpyO
ZNkX9/HgTbBDN8vEhJINQTmqpt5jCR7b1pZjFm0342kDUHk0PtCh3IikOWoJlgHI6gA+mD9VpFsP
yI9SpU5E22E5zXNaDYnx+yR8QSKO2uaLYEURoq4p2CrGXp4wpjbq0WuAmYmomaVi5KJdaunaj1ZC
VAv8O0aelvQJO0zMfsWuZsdNuGtglxmQeNWKb7AzajtU/5L8uOXic9SesBR30MmOunVlNw5xDaXE
L3W7pbkRck96zCyunln1YMNbjh2UtbW4yXQV7WW+1rnLLXe1/J9AQ5AeIqRPSBMUvYeWe334dkT/
D+CRnut/XHskzq4gXooYSpJAaDawsBj8VUBQ9wMjdgJpAxPoX+MtntUTGYVwlStFZ+TqmUr+aYWz
ifCLpi0j7XqL+VcpHOBU53TRnuaLM9hCh84ITNCDC5eWzr0tMjKp/AY0k5JtD+lf/TVeDmMylMGj
tmEdP0aE55HnkrldIfMtV+zNceiH7hiwn6Iqystwhlk5SnYtpOVL+i2Xn3ZUL9QWWGM9VroYzUiq
5NOaejEzZLCkrRmnuq7yD62O/5saLL/DdHTzi7/uleKzs1FCiKdPOWzCiRf/5Rp5gWm95U61iKII
2YwXH1Ye2aUsMf/dk4GEgxvDBmfRi0JeDsbhAHKLqZGnuOE5iH86Ak/UZVTRXepvNYTHLkgs8PeD
7VIA/HZdIADh9xhmqFgh0CDz47ettkyantYhhPIRHybaeLrcspUxC8tBLesauCiiR97c7aQ4Rqar
u+QDImuR48f0nR4jJwtsmiqaQrjCHbmY042BW5UjKMoTpi5r/xsuUTZg2k4nWdAMiHyA2A2QXhg4
x1orWOXMr9kKhD30XJQR9Ba8DKc6fPvB1zxcjV9bZHoDJaJSCspo3quHjeQSkbZsFhnv2XC2KPJz
499WkC+YRg7IWbdYwG1HaDvqjfUznntQU8zQDm4jns3Vq/yqLF5pHYU2mnscMRKz/0oVoHlgP/+1
hcu8G++SZLNI5Fx9CtSRHoGfqZw8dqL6OmK+5v8NBZNT2+leEcl1u3ZGGGZ2VlX2CmoYTsqndanw
tPim1HGa+STr2GStSlZMbZ2Hgh7EbMrwxePEwaVa2qSfNoGnUMf37nyXMxzPj90D8kJsGpczI2N4
9kUsbE2RflGc+zmOkk6zdRuvlFEtWab8Zo7341mGw/wFCz662ZnqzolXKL2PntlP47AbjWJ/jyhl
K1w+p1HOMBGBAV+XYh8JAuKH1Mh9qi8EDOp7oyEV+QqEiP0k7XXkczwaMW6XnwYHCMTxDq3sDh65
YQcAfbWj5hyJ0oeg6KqrsWjtsT9RKYfEw7sIySt3NPtVhmVvf2xX9cOWchEk4SiMeD7N6J0N1SBV
a15gRgRqMjUIAB+S1ppsludTM1S+/zs8qjPs8tFeM3wZRL4B8FQtJN4t+pSWwvm8T5VLUNC96tpt
6roORqt1ey3Ps8l3e0ITmcNsegduVSbS5Y2nLjTwy5yNR+/yxgzawxdLRWZS+lWk+tO2CsDbTen/
F9zfOD1AQeR2E7J6IpIaql18+dkLEO3GkNIJh5DpxYKqwmfNzQpNCajQDNXF1yaAHPUczVMcsOHK
9PyA6yl0IJAnursR8Dx7sstraoa7mAWpqyo1E554SVz8h0sP+raX8RN0aU2Tmsecy42tb8DTdPTV
vBTlIHlqt7jgmc73Qox4wC/NpL6UUWg8OFES8u0WuI0P7AiOcILYzurYytQFAb7KdxP6nwpp0Eq4
mSwVHpUaGa3pNRqnuDttLmHGGkc45nebXxFY/bkcfn5LIKhLBVDG2qqM27mED4FgXqgtgtzW55PB
lJC4ebV3T6iWScAPDZnA+JuscalxIuiIcYTpgfxVerHscblhITwkeGSSECbNpQNV9i9yBASWW3Iq
9DChkn+iTn2N925Q14Arh4yMgAAdL6ZOcBw5Sz5sRqrdNKqmvNQB/JTB7rbOPdrSpjAvrmS7t4S4
ovTQCBL40xBOsi/Fy4bAC4PgtK3vrOydwThkhQV1xB1IkbfsmpE2I5Peeux3aydvT7VqtQ7FE7p4
YgvxhW9mSy+JNUf3n/akiGlNH4lxWe2DFQHo5VF8/ln2/0vR8DQu0tbj0q3o8+i2cDaLfBHQrN0+
4wMKqwJg+Mxi4eNcNG10Kr0MtYv6HJjtm45VFhRZ4XkQemansIOJxFIULEpN/h4GenN/PD3Wlkic
LL6XIjtzN2nscP3hfK9+IHxQFE+P6NuTQr74gVMGqQyEiQLE2WKAuyLfrAlP+Mtso7F7OX4LEb0k
gZy2+pmXn8n5HaTibQj/cnA2n6lIiMMDU+3TFXVanrBMf7h93Daq1YsIHn0zV8tsSJ9HJQstht0D
Cse6EFusoyrXNdAB7xqBaIsrXevVDpnFYz6UY6C06iTLa/xftAMUTPMP4KFLsWRpGy5sBeLq/i4A
t33sLkTpodDRMV4Vlzxvfh9F4C/TcL/28a4FtZw3BLC0t8jX4XmWCFihIE/o7Lp+Fzk35Zlv64hE
gam6H/z3hZDjiCNSjZnEPVYK6Gnhf06p7kQWCV5KyhjVypdQXN3bIYeKSlK2fs08zplLL1kv7Mus
OTj11pwSTPmNOf0YGvGCsMgthYJrvRbCzTChh4TITL2ihOa6ZdCnhzumW8r7q/ifViqtOt/dRJrK
XDMPArXZR/uzcpHIhegPURHbf/jywvz6V5O4N9Jjm0vu0v7ebtIhQhrLshyLmCerYa+cmKSUkar9
IblT1wUES+7yfwboE7uMHFzfWm7Pg90f0YMRVNOBRbo8VjX8L5g+DMZWt08jD7k6+W8NGk3THdYx
eY+Ml9wYx/D5sA5KBnmW5cS/lBug43Nc0+WK03bJ9ANuQH83kEg3BG3mUDy65Wz/XdYehX1Gtf7+
qROaHLAzlsG+RPuI87NHK1KpfqD8fQdsH4uK/t7+44OtIVoAlsTw3seziMPSjdqOjRLjNi5435cO
Fb+0KoT6SbcxPHGbd8gi0pdnSVy94mj8xX7k7mGtJUaHpEHzfW8QYfk+lKvJPnFQC4JNZZhnwb9c
ai3qWVI9K5D+By5wVIPS/FWV0tW/9WksjvcjuDZkVBBqmLSenZ97XN81i4P7owIhL8Pxpr0HFIl8
2+s5sIYw6Vju3OiliEmsH3AB7aewmdZSKevOwTuV3qDLZ2TFeP+zb2+YmtAS9rPerZF41sSOIEHZ
59/unXS1eNPFrFsdHSwFm35L4VpM+vqoG+IWbzJvRN7+L8+JvmjfhSN83kEauB4Pq/rMD+IPeKFA
vOtJZhLrPed5JABnYfjQlRvVruuMMUDEyaFmP20EQtgoBrFTMgg5e4IxV+4406lNodTE/+ht6gZG
37m8KJ1+ZPc7fg02O1XvCZDP3tGelbJO1eZrL22KrJ56VFUBf9l0Yroja6HGubQNAbofszMwEDdM
8QGDOiJTLbSuJsSk+HYmTxnj8vFs1vOG9wP3bk3dmkkIvqx33hYzCcnsvFBOG3A3IBWFd+hNJamh
aIZsF0fttPwTZ24td7JbtGo/f9OZi1wQBRnUQQ9J5pH++udtwxmkmauCBNBIuD/Lo+A2Cv7WxuW1
PWWV9ldR9uu93cSwiOiSNucfb4A5Fiv9J6kjC+uGgMXe4EzzVfRdorfyn4R60wyTan9bvADe2VjA
4HqIeVuRzb9Aor8yNZKj3ASGZ9atdm2h4/XmIiy+1/6L6CHkd/PydG1mlApc+xYz5FiS6vA1BvqU
5VafXOdKpuuaW4rUzkGqXrTSchM9VBaputDmAXcKfa5cbGuUwWW6MWFusyWW94Z2rDNy3ZZuvUli
gpJ+O3r4oklddMPXr4S7DtxswGdj4SoKZiMjHp/OcvpU+X8jXadJFGG00/5lmEvVD0NqNRql6jz4
wzY/C9PscA/yC/6pJ0FEn0s8Rcuna+DzEilI3xyReLqE9ehtkLsZix7qDteSoIxfJqv1zbJbh6p2
T3FqnyBjmLlH8KXuJJJwF0+j+qjU2ikIhW6fEu+OG0GIj3gjHo3z5tQ1zNo49AtSXePVoP9FTGQi
MH4HV2Cg8jrPUodbIpvEoykLG0qoezClezGGW5I2Qqy337rgTRWPigK2g7duJM4HtJdt5U8Ldk8u
hv2t8zt7X3fwrryw2eR6MI8/1Ty3NdwNhNxjWe6auInPkCZIUi1/FpH21lCQjqde+hkpuVpIwtEu
1eTPfMCJH7IunwqswHswXXhZZKVcZKSkxe6rXB4a0edkD+Q8CDjSSfLXkf9+19n3DmVA5oS8B/6/
KU5oghmGek+E3tN9Lrxjpp3wdI0ER+QAVMf4+Wq7pgTmwLOAuZVQr1yrX5O9Y+gOJlM2glLLU8YH
PeYOKMCrdnL1RR4c0UzFwF0L+m7e3bDIB3DUD02HyLb/A6lfHlEkvrkpDL9U05ON6ht0kkEaWCBw
o4ZSw/C4aChpUW8RligLmC12JUeQgNGhsqmDLnzsgDin0EMLRHH/6L0N2/KIbXio6ItUIC7LAaVG
TKMBCVvEA4AgAh47Ks9je8Au+1kCfNTjiQ/c2+6vimw7qszRfpHNvP5J5sQs2TTEe+9qBRqo3f5/
g1TMluc1otRmiVmoUguGJ0guRGjVKAj1sbA62hLgBeV+AEci+D53Is7HWz2P0PG2Ity0bVmO88Lx
kCW7dlXbhAgYxrPN9bMR18lcpDDcYaLPVmIliaBNfLt+dMBlz8BEaUhkbzM2iedwjCDLVegi+79T
IFEfE4hLZlGE0HO6ueLm3eAV8iZcU3M9Le2YXgsZ+fIHWSMjdIhxOuqIr2WRgaY557XKXS0a82Qb
ryHlIKCgBZRPSS41tmaxoqYd0wGznSqB0/kVIW7+Q1AZpqCJxcDYrEKtiLh2pancm/+wuxKhwklL
iyIIzN/LEow6J2LkMHg5vx5ARhzqfZRcwWJ8s9RefmDvqwUARchfBz6iGqmVSgRHyALGwNpqI8da
36/c5vMehBvbRwiO4DoGr1ivdXOZTObYkAMqLCQ2Qggxt58umu4CzgNPHlERRLhkZam+6givUzqG
wSm9ZD1bpo8OlLEKkqKbTNY4WCXXETjHtaixIdD1TcVO+tiBakCCQKvHjK0aZhzknEYdpA6VM3jb
mAK1mgLmQlMo/72gwWa6PcUZn0wB4gfoZgzaIcN17GXsrddTJJY3Gbog0IRz0iJTYH1hXZj0Mb/Q
V1PLsWH4HlZuG/jfu2uh9gSYzZ0/FMx4VX5z/3U0S5AyxcVUJqB7IdCeu+GmyLmE/wRoG4D7t79w
vAdnKGbiWTE90yeoDYNs5F9F7xmxaJJHgmY0ekVcQ3QBsTmdlfV8GE1Nk/X6Gbq82dlI95yalXll
II/PLImuaeoNydA0Q10xhp/GGR6cm50qFzh9OO3OJ4vMmyI4W6lRRu1Cgoh7POtPpoil4PGZq5bu
ydmeKlLZGq7qfoWoTo3AKU25RhS/IYvoq8kZ1kVidYh9MKvWlU3HaWThbh1bzR9X9GuviSWDoZYV
KSU6cdDyZ3uwsUZYJ8x/3kf1IwIJkndGentEO4F9OFKHU1qFGxxq9q4lLgYjsSduhU3prOOwhuW6
X+3ojKmyRNcjCbCPqpYfcoX0+t/p6so7xXkFMSq3AJRTlPiusjMzG27x1NLCLAXGhYwGK+OVcy01
3TMc5hYmMw7iXy74r7yKRgibFfJVsda0os0hJz8ri2Y1xkjmP53rnjqvuh4NmT1NJXDefDXnKeI6
XF3L0KAXC7yXmrAPOyAB49yXjAcmHvBoQelgdG+UPku8Cjr3k+q0bu50rRZYaywMpwLdCYM2ML1J
BzmOS9FTM9bp4jzXOoH0Mhgz1DeFHzoum0tcwIeLbqvQkKCVXGoez5AmCzHQ8HW9OMFrQYPGl1XR
aikbFXxb5Dhba/kydlki3cOELvEciwFGmuckbWLN5Eye5pnG1rS/rNZlHRitc6jc83m49kglXDED
D1dk/WX4V6O7g7gEcti/dKEH9NtkpbFeZxgOiv63g8UZdRspTamwT0d23qsi+kYnHQYAthO6+rnD
k+eh6piAuCvvC+MgakXN38kaQuob87/y2kdd0LTfIcuEQiqUVrCO7heA++IdxD5ZsBgc9ZieLNIX
vmmISUQLIl1olGbT2889LVkFQp/F4itdmUuU1Yox4+IfUmdJvDSWMKKde1HQND5dah8jMHncwx7H
X0Ri7AUQf3W/ziaoFY5+VAD5Q1y0b+QYmHg0PoejJyuGVqzhATbxaNeYzfn8qHrBWe9wQEQ7j9f4
d4tIxtH/qTrvq9MMF4neXWA2nZe479Yz3hsv4COwS6Ah+iT/+jJzvcb/DIAuiTfUbAbnAdpWjHPG
zG+idshrjkBp0fvKPCRaSKmeXGU6STX3x0+amsWt/xsZzMIh/s+7DfjsBxT6mjkgOUunqbAIhdJy
iD3GxijybksSgIIHrwgucb+s3Z7TY2A9fblxAqwkgr50O3vV5RUrEWGHvmlnALjaC1fC6iHFfXD3
Om9AP9zm9AlxBau0iYBaSckrUrfyKrGi4eujkaKyRN89NArcKj5hPn9A2jrd2+N8QAru6jNT8UAx
/VTnVFII2jJIN+ArnPvqsFLXdX0ByC2Xf0eWDqkaCUwyX3FRO4ZKZzKhngNkFz+mGXUXyhaQfUZg
yp58Hp8YEnRaF+XH4HHC6uTRww6JnhLvcsQgB5f3jBHaQQgbQKHGjufhPc4ybl/QCciNNseoE/XH
sjE1Fn49uh/fdMj+KywlmXo8U0ohzk2c0iOXeHzXclCKz7UlQlYlK05pRUYPWebUSpQFYNPJtC8g
kSoab8psB9fBsbORQuJA3tty7RgCj/hlBTkgwip0Qinfy+RBm3bINmuv3clVhEuKzwnBK/pMUNGS
0DuUMBo2ptecLbtqlQiozyFNW0YVpijPnDsJzjSVUaI8Ty6gCDyj8XTq6vl3GgU2b5OMaN4t3unj
FPopZfQtX18Cpfh0pHHx/3+qoOsGu7tPSikRHpWr2ZVPZOY7V3vRFytdNAbBWvOs+OCq2Te3/KT5
VJl4MKBtE41sXUiU3iTqZ+scJJstiinXwS6bcoDshQdcF5PhkwboZ5NWqvrOB1vwSbkMClnhQaVS
E5slkhR2ohUyI3r/zdFu0BzO/hB8FS3i/i+8LCEU547YXsN7GikMaiKhTu3J1adXcUk0RJLhr0q5
awhFLBcY8Y0IB6kOzCRd+7NcPTcNORJOmjmwmc+0b7tTYh4rSHPzlmQvZnnQQaqEnOgGavfOPKs/
mxlJHsul61R2hDXxl+/b84AiB0ZUSXK6kR3oWS/0KsEXq8ybb4qlX3N2qmnYF5doonHf7tOIuCto
vtuyk2LF9kcx9ZRSvWMzpfFhQejR94UulgTsHES5pobx8N3R3usbUdOM3JPwK2TOS+H0nJhxviwR
q7+9OFo0f4c3xpcx01Hz8vJUW76kkzD+CnUAUhuzNQyc3C90cUf0brBQRntXQhgTMcktd0yY+p92
1n8EpUgafTPZ64uiA4Dc+ZQarnugD0WCCgH6bo6LMWT9hBuuw3+7ZpdMJHIg/mnboTNSrcLPKZAr
8ZtIuwwWohxEkv4Dh1ur0TfrClue5sCVntr+f7+w9gBAQHAqbl+u3rwfRhg7P3BJUzILKMDDYFSx
Gs8KviPEyz+a9lCde00ghfv63OdUWiFPrlCNXOxSL1VpBp/58jxmjn5VIXgN07jdxLjqNWZt2ZBo
YloHqMYvXYO4zTtFA+1aKrUDC0Dkt2d+HzdpuYq/65ePOH5Pt2l6ENYK0rQYn/oatg+uryV+bqzX
150LHKRckdbKdaDwZwGTyKJ+HrIhe+jXa3YQIT/hpfxWHw2NDG+FqEaTrASOxwXl8PqODngqVhWK
G5BXmf0al0QWlBZ2nbP70r7MCYX7UgqAzrmOJTycv+KQu5YyqJyvU+toCjLrt01N4IQgc/0Ue66Q
hl9BQlJt8qAOtNQVRFyAte1VcQiyaVvxDoOrohxP26HkSutKPlgIOLC2a4BUu/AUm5gk8jvIgC+D
pQXYloecLnziP2mb1wJjuy2fseUOIimOabTgxPPv2nC/lMnsZ2hVfh6wHaL7XwyQsePu56NWQV2a
DyFuWLR3GJA4XUhKZUvD7WA2uxAaTdWme4LnHMvjhRG6XoDZ55364RApkzc422x5h3iGjmUf5Lcg
e/dAYj0nVdGAtz8b9tYWd1fLVc3iB+oyHiRpZbrnMk0kKdKaxRAEl6o7Bvi6TyOoZ1Rpjw8FBkmM
TShCVUvDeOxXSygRvfmfJJa2Io4lB+snOo/XaPCM62Jtz5JZLYbfkX+vPZfpI55cmu77wv13PvSg
qy0xu98HZSpNpnTj94QcgdIN5A6lDVWEnkDRjezjR2SCXJa8bvXv/EHVbiPrfj8k3Tpxkn36T7NQ
H1eFD6YZL6jEU6+czwSHkWqzEkIkxGC8lXMjaVkpazTUnA3MS6L4oY4zz/TydIbred8c+MKCjznF
x7wGNlEIBYmSjIo1O3PECdUuMoeRNpydIhOqzCeNYzcJ50JPGsadmVk2OGLsaE+ZUmFloBvCr99t
MdhV8fYQmWWLQaefDsy4+YvkjPltudo0IXSpwnh6vf4LOB2uy/snqk4Mubrp/XZOkU54u8VrUPvm
A6JA7oH4OoxjNh6ZPUlswPTxkhQjChAI7AN3IYCeS17CcISeIGaHO+H+SSkUUHUpOpUT/61eRQ/Q
oftaCYHMntgRaNIX6zxQnJZYVWbR0vM5TYCy4IDIkJY9Ke/xrteXcEtoXJfwyq1K+bxW6+O64jTL
PiDQMrTfoAE3I0Je/oCzc2FnbRefD5ZVSUwMRR6d7hmvfoxGnAYBWMIRKubBytzpNBMzrVIAmQ4+
e3mBiDvrHUwjoDSIz71NmurTnD3579WaCzh7l9k0hvmn2NRfeeHc5SL9bGg1/q7qr/BThJZYf2VR
s+33vDlAqb/Dt96lp35hhY76COs4dTfSwLvRybuFha0JuXi38IdNfAzMVKCj0XBzGHm3dKwS/aN8
RpRqc3X8U7JufxsLMAaOZGZLLm8cv6qBLNMYk+1O0yVBVRw1Q+yuCeFanXQEC0n/jfy/aIBNYshk
WDO9JMwPonCy9aqQyjoWgXN4wmqV05VW3McER6Z1nm8yHpthv1R/D83EBaRFGgu/bAgFLXwOg0gg
XyRUUxS8jLo+z9Xv1Q+IH5WP+4HofO2aVFlPO4emM00kyksMhmHBwQ4te6wVa2tr0CdFBwZDjNqw
zYqdErHDAqP6Esm+BYwUxy53F1rA0/qD+UN6Hll7X92wSHDYWC4GAAFhfMnR+1EOabcwY8pAqUbe
fxUeUHq14UiJAX15DciHSAhdw4KbXxycKrNhtgrR348ZCu60wjPpbbfelfJl2IVA/ED3hyP6j3zR
o9oSLRLsZ9r4tmjv/a4T8blw6AfHAH8YJCrppiSPwD+HWpBDSH4GJQcocf2LKk11VzT9KwYJHhLK
M6x5ixEPm5bHEV03J4LCjCiVLDfPfYQCVtgAJ2DZ5pcNfcKZ7GxSUKu7SFXQxbPsSSkDfTwol0zj
B4W5H5EhbQrIZZQPjyMdj46vru2peyI+bMcu1bo9ajQxDHCiaRZGqN9zeXeMAlUggrq+oipqtKZs
+N87Vw37poSrA3k/k8Gs5MGPqTGJTge6E6nbjTWoXcPLlh5/19jTZ/fNj73+urd2Vx9x0O3nhXUh
dKP0v4101PnaGLfl9MI7EK5yYSYOxa1S87JY6nQFjJzGluPOPUQbg8cqt0qtwllvdKtngMkuoeMB
GzzkeKpw3gebTIHlp2Oe/XOw8wF/uEQu2QdDvDcD0nIE7WJTazfGvEtpjtM2ao5F4dDzGEKY1qZq
LTpuNjDorbOp68J5IpE1hqd+F8PfNFEEX2sv9sJUxlku4tckTYKUDRKMf92Z2+cfccGfb5hEOrhT
g2N86LBkORNuBFftxn/nG65Awyhldx+W2jqCFXA2at5Q3Pb3tKfRPljS4oyRp7qMkO5YYUWelyY6
XkcSLHCVH1S4qMIcMXrCVNLxrEVA7d/ATpKc/XAUe8MnwUpDHDxm3bMUq0ZhWHLHFgkA81rGCW4d
h2H+kEsIXJurCIEWCL10soTFBFDW9Vj19lyvZGLPbbsVzRL+JXC544TRHVevAvIJIhNLtE65u4v9
wGM62cZG49F7G3bocSSIJYcjM6ydDDlMm6WH19c4b4UgFC9yoJ/MMoErbAI+lmv+T8FdIrugbDM5
IfA4TAvjM8KUHZ+cC6lzlC5MLqCNeEjh/LspO56teOJmag+1lG1MUrHBc5s2b1WsIFPl+sboZmha
AxrwfYQl6KPcpCPikKQioFQfGafaIne0M2h1EDdTYnqmcBXV5Ilkh7kXGYjKZsaQPpRYp94J/R+B
ZXx59+fVam6aZ6LqLW9mGSkFQwT0wDeHs+jEC+3jaAPDoNXyGVO59PKb1qvFq4iBYhQjFi9W+iK8
P++rNuDulpEISkshXXa55xQvXyCKNisuI3Yob2bOpO5xteEqQvSAK4H3oNlqZEJ44Sp51yAAsIIE
P0GjIA8dcDqmOVwpZCXTRsklGjsFCuAo0/7TSap1960JfZWHdXAPKDDoVtI6QJv2rbHNLACdvibe
Li7ttE/D3OGesC3mm1oDvKVFHyXW4bNOXS4UYhLUJAaz6huekh5bYNmcF3UzN/k/5VT24kF7fnh0
ONbv4hN9gKRPZq2KbkMXlIdC69Pp164GjSA4y0BfNx6wl9RR84YoLhH054siIsmQHzbveBCm2bv4
Pj/lPWe1OzUFpU38t7Z4OVOE+Zm7+0xMoRIr2AhNEo7c7fZbzUoGI0/m8DFL1d5P5vNy1pVQyqY/
4uATdIC0UrMWeZ0RFpyI8rMzFhsdQDowOee34exWUi3xQIqEALYQkzyeeZea/fnEhil+XpUlyiW0
yhMo51qt5W2OWC6PElD75Jo4curw5jo1eMUtQUitOcVIRc/VKpLAOeD4tUWJIYRXd9Y/1dogZ2FS
6fGNctAkQ/5xGnKFyEfv8PUwo+A3w9sZ1s91SWNjFqZ7hSkoV1JQmyaiGMHq+CQnToHeO+zK/KsE
YLlKqKlNEtEooS3SauQwXw+Y67ketj08IiY1ZwL+2phTc6M9fq36dabR6TYjoUwoHBabIH3PR3Ca
VSneRKI9HwmAs5CGWcRG2RgRpF/3KxRc+rjiVL5YJS+/Qp0gP9wqkLjnneBOCmzFwUxHy5eXfzsj
dAuMxYoOzkKAoEuwa+h5xAeNCahrfZsnJX/BUsnDx3jeXWijIMnPCba74wXwKROlAlNSRb1ITQkn
5lttMzmB2vtcqMJtY3mvMbCAs8QFWrYPX/BIKFxs0cyXYYBpt22viRgAq1PrbVh1197FMSZ0m+vj
JWk6aZIIsWc42XGDItbOuoWJhmH9AmdoVYEyEyl8wi3OScKX8ukO0c1aZJaueh/fOWBesx8S9AIl
6NN/29pa6pHWyUELd9rijLqw+7OF+SGMGaV4pf2Mmgrzdt9ipCea2daSnNT6Pn1bOyV6LErtUvPC
dCsH4jJE2OWqnWUZYbc0hZJs8u65YP+pflihr0Q2Vacym+EsFqiZv/WB1BD/WmpZbDnOERteBoIK
0h8MvLR19J7ssHVEhd2Bd3yzneaTQEMik2cD6sbI4uBksnD6evcg0YlFKoZoHE2mhGkH6T3LYvES
loRe3FHMaiWlvSISRCCHn/Vs81mCguO9nRMCc+7BLQny8Ie6JwiSD3vmmz1lJzbPhNGSmqsJRD6O
StQo41m/UBUxi1fwt6ZHHUwMs36isXE4LY1MEntlneFibmPioUnG5yzC8+H1BJgkoVpg5QusLlKj
xDD9ktzeDtJoMCDuY0/oxoQHyEyDVhwKPEblZK5pYLqFZM3OFnh1/Np9uObzMyMEOntogFemQS/+
hgDUMi6KitwCdvs6jKVN+o33VfX3DJDe8vV5mQRJlcWBlIzu5Dvlr5RMGY3rCw2NQ1tnVGt9zBg4
5Bo+R4F3Za8Xefy0TIFsi1+vtUJw8bu8D29fwMHZJLqg/+b1v/zbclGm7uyKnnyUxluLLvhcP1Nf
wy0teLxY19m0Jh/2z3Uupr+5YuqIa72YswRYfz+/SJ+aqeYzeQE7snZCw+lrRQzpwLanVzhwC31S
tE55prFIJWa45sf/BfA8NIHTQ2ZPqcsF5OkgAg3ImIxzys0Lc2sd8SpcPOQpylo9tSLPtUS60t+4
qnexJfXxwHkyGPhLKeoC2hMfSpHGvx6gLzrNwgxrQf+Z7fFdVzB9zTwqmfSRKt9E8xNM0AWJg2GV
w+sLFLsjH4/7bgCgVI6bxw7WncwKBj/9IvvF3dyEQwRv5bnnUGjwNFU6WdhY0/WgX2uGFZWlmytg
iBhj00d88DfxWKremLjGJtiZz4pSJXXDN3I9Ekc84urAGfCtwacnH7MMdOF1dDLcnUt7yINDbG3s
LoA48MsPy9kadKFcd3KTIX5BZRG5TJIQqnOHMx9gjZN1+HrOZF7EzLVfQZZw3ljfVfxoBC8JkwNs
PtIg1P6q8aOhdskxUv574/PuDt2+hwCLfkVShtMDQcDLV4hanLp9yLl4O1oVFfTCMVDcXuWbXlm4
r9loRnPgSxRwB6gKORyVwXfDxgeKtggsNuBH58mFnHIjPW5kWR24bp7qsEN19Eq4TT6GJ3f5ex3u
9xMwVGb4WQlUNGNoKk4ee6kU4+yEW0yfkq6WEwgySFAcZ1VnTYt4YVtttji/kVmv9ugYWdXUn/ks
JpXwvSVcikmhwNoW7dGA+HQumHR/qC747aV6YqsABTWRIzbf/Aik6/qiXCh9aXHnnfpmOdNzP6oz
kOOJuzmxPnWN8dtBbaF7MKRJqhU6T0LeLIK4iTRCf710M8WpdWoGvkM0EJxU3gOxLQugkcnLYvkZ
mb94iz5jpkXdMu/ZIQk4VpoW8TeVj8ZPBDvH/l9OaIc12qoDjOjTDd4XhAOB3/H0aqY28KOeA/8K
WKmT7mVAjW4HW1tQh16FiFb1mgTyrbKXlATJoNwbDUG4TzbLMuqWM4XzYdO8kozhdFRObZwtKRFw
18BB5V4AIlW6ymXQsPU3qi3pjNO8S4UTwAaXSSicR3lKITetIxzJco0YJMsu6I1TQdlP8u629CIw
8Uf9eEaal5PovhCtGO7qW+gC8VI4KMjWnnYrNrRN7ozMlUko27UYEPv0E9NLTWyyo3jl2bamTwcg
opzZdK2foVWWTdgeEGPlbYuMWqDHYx+/0jUvAOVXM2xHggzm/ag1sbzrHEBSPug34tvhDZ/sQ/jb
kXKDTLd3n5JT+5IC06V4bnXvPVwgQ4NU0FePQiPqMnKKhYR3K/l5YZ6WdW6R6tAOpgNA/QehwFsa
gWhwhGyI0xuXQvhdwiYtmyb2Wxc7sk3YCaASFM7OvwTj6t+F2LEpZuYNhSiOqXzkBr0sFW7toy47
tEnnRrARUsSm+yfdpMxtO93b+kEZnGC70UFuSQB0AINe+E6hdTpjYljvvdm3PPYXKQCKNKL2PnY/
+HtHUnQuHhu5/XhY6RNJNCSQderH3m1+QC2MsctK0pqZX8g6JSgle3Yp61xuKw0DKJYD3ajpOxYJ
4udGzStNbSb9/4Z9Y2IB+v8fKXbrNy2hcO7DHaOaTvNRwidkguR27c7C8Dr5BPSrwxC/Xw21RgTl
R2P39/8lBz6uYMHJK+W4UyvRyzXn+zMjNvDlaRVN43CJXbLt//JhnXzeDi0coBJlINVUOuNf69F8
d50GT8dkScZTb2+eIaVz1nu83PZsQZVFW1HA3USmadrEs0RcvYFL3bfXIfvwO9/OcnzcVA4VYgTK
if5e3m6MBfzWeGsr/3LYbFI0qXMBaUNOXnrX/rW9LqSFVfAy65zkIgInnRt1WnkH0O8KXdaiHrWr
hcDq34Ijgr0OsFhovKmQrW/1vbPhuUog8q6Z2qPkXHQF+HP7036dJBo0CfHnkvOARghiIQs6X37N
wcHdzJG/i/J9K0OizCgpwtawn6k8FGsQsFytjTmM3B+DIokQLaIt/mA1/+q6vtR4WKG3az/7ZcBS
B9+H9NfKB+g13MHQxvI/hiY3L9cFFE1+x0umbAUNBwonaP3z0Avyd132fb0LtRQMhgHs6wFXZsMk
1g2L5DUvomGu70Zfkh+cznOAIheXKOkQejwsmIw2/rrtoljomAyilePVBEJC7SR+CFU/OKRGT6O7
7oal5nEPEecrCit1mOJHXf1ErjyFvYk7BWPrLvZ4X+5XQ0OXOMM1kUzl6agfllH4eIKStQ05md+o
y0RPYBqMEdQEIM84/e0HkRgweaFUNkGJC98S58o61s90ThDXu7vD9bH/qre2li9nzMg87G51Tyxv
jhefe0bjVgUCTZjx++NFMx2XXyKGwkaGmZwYs7uOs+WTFYPKOWBp2cPETTmDPKdMtFZFChseIBD2
5C/w8yIkMTt+95R9ZCbyqT6d/8qJ25iX8IKZJOfuK+AnJ8Hu56FxdKi5qpzCQ3NmEpyuOXPArAWi
OpEtm0An5eLnh4P08EMlik2zFOQuzw8hvIHBz1XRimMiZJsD6kgqrbjKOA7DIACfcn4liv9XrDpf
Prvlnr9qOnZ3Ng4oH3p9A2eKAE+LhqqAWzgK0aBbwZpPfDFWUVCeASIlkppWbjY7+bAecHvVUXDi
rXJvGr6J5isk3pp1wC3DW62jobnj7jfItBdLKBGS/qRQSCPzezl59WdIO8mVP99nXJ/oZjVCusZL
iP6IgJs8ZleVbdCFzCKAaTZ9Fahb5850Sfy+w47Vx/7Ad7/+XVMOdVPpWceps0PNr3n8BRtv0CsY
4PL7nywLwLJl7iEd1E4ize4Wk+ahjJwB1O8Gg1m/kGpR9m4ZcCNdg4orOPlfy1V/dQ1vwXCdXbU2
raHZoT82/YY7oKNQImMKuCUxFJZEjjvKBbTiffeZknsvyUdbIG7Ud7XUiF8hEcm+sRzKfiwhoi3T
1f56omi/Hi+1XlZUZJxYuBYhvKYO7s3De1HTeGuhFzLa16EyhWIc3EG1c1EeUwZydniiLf5abTM4
ejTGNQJSLuWMvVUv4Q4QxQduM7yWzftp/OOMwiWV0kC3/H8zdxmd/E4iDpyb2fh4T2HGjrJaNfuj
COkKUUYsAIzWxndHiuWalf8KEXuwf7Ht1khRAxx7L7aHCY+uumuQIoQAIVPSXHOZcJ5Lo+6vqLPZ
S4FY3ZOVa+pfIU6jh/aGF9NQmXAohvttIu0Dzmn05eJiPvVn+AgCSqt1CgGBVyttSB/+x09NuQsR
MPLVMb8z2DBkFFbyFc1WWvCFKsakhdFWYmC6LY3+R3rpVURbbH3TzlWrzkAt4LegRj5v6s9N+L0V
0yP2Y+KGLMgM4J4NnJHSkQfTT3Y3E871rcJ+4qxB5zPMzVoPzLFq8fwaf+j6cqFy4VNG/ugD0NSc
FckY8aGmtO9JRPziN5d1qEI31TuzwXNpObcrder0hdelUAL+eLXHQ0XQCQbAKvVMuA7Kp30nF9cN
faw6lwg9JGszgMyfMXQyNjZ6YZPHdlfR0cQsag5hLuNpwWO7a/uF64nYEuLApXVtR0yc5VRpfLxH
SgZW+GzxPbFtwFWLqJE2GU0GAceD1eAzhOJ9IOIuLe4HG616F10VLhiVBU0HXjNGo2haqHd47Fa4
8uqwldOQdWDoAsfe70vyFSQ59blWNd/Ou+ZtoL7XixtAVZJjDKUKFjRDEPwmQ1TaT5XaybyXylCh
vVFNMAe1vQEtrnoX2SrRGM4FW4Mc0kFGpTv5lUc58pkrS7FpeldQRUUfgvNvp2iuin/RPmQyky+d
531sjsTn5aSEVRLaWw6dpSwFDdsN6MSH+MGbpC7m0CPGOndfMU1NMzQMlkABvo/1lv+5ebZqTkJc
5gEwCnBvh7Cr+uYthOnmmYRC1C3km5yBLpzlsqOXcgpMc3ZcvKLXZnVsiTHxz1HlkEeQGTBQ4fwi
1dVvKY/PtlQKAPESVEB/I/K23iBoCBGFIeM/NuGtraXznD8tQhLCAd3mNtL0T88M81tu8jpvZfHH
k9ACmbhpOAKdwqpSrU51H/sk8bPHT0UZ9s+H7B+5upsgVh3h/OWqsSe+ZQo/possb3BEseZBcArC
3tIgfk46Mw6LiDDhtuK3HNfZXAbl4KHIbLt6R8QL4yRjTYe/p6GdFa1mfX0ghjrTQ1wGd4W6vBwJ
Qxfp7jhtZP07qTB/LvJXv9mHbwA3n9GWcPu6x/KU+FwGnRzfn90mZlCk9w7WxaIJ4h71pBs3xB0T
1PhOjtS2DNCW2nG3hLsZo0Lrrrx+ENz9SMK/in8pcqrvGh9ifNX8EdvIJinJ9AyO249eywb2Gc9E
UeJWZgmp8M3O9YIaG0LASPJXr5iSmDay+KwO88CFa6wJwMVPrJvaoUgDHrJJsNY30crIIc1HLF96
YV5k6Y5kNJCXInwuwTDHQb32vfIDJMte93yvs4Yi/kEC2c59k9VWTF5x2FlM43V+VhJGxf3GYj1l
E4sKPbHEzcNRRTBAR3Duz3/UmA6MELF+l8AdQfL1JZW0IM4M2H3zt+Trxm22V430lqD8YUsLQ6Ec
MLmni3ixH/vGO4kAOsTvBYawyLVgbegNwfI/Ohh03iy6Za6VFSsipUlLEcMLq6sZWh6XK+QKSvI6
MksiC6jVh0jqeVaZFGbcOdWf0FpuKqvEfQf6nkRk5pz+xEsE/kT2nE5uJfGjEZGqSMbSHy20tTIs
YvMOM7XJqiTCAgfwZ4QQ1Yn+KNTwWqyKgsKpLAsIKRStz6tZb3TwKXSC1nLWXhOwk1yxyAumWrhn
QdDMfKS7EW1XPXQbJTzrVsJzRWNzefvVx4y3KO48Pq0c9OqGnOqsebuUPcvDN06yTKlTlZHIKFtT
LwHenUMwxs/erY//9WiAo30CQ33jQ4FrksTl6EFMZ2+0D7Qv+sLWS+K6Tj+if8XA222jMnQJR2qE
sqGvmPlkNgCrJ30IEJP5EI6pQMa1VkfM/0ZL8MxuKJtSeRrycc3DLKlrce3Gk+ZD8goO9us3CEt9
0l8zaBHk4SCAjL8SOhcbsUtn4u+tGdobRs3G3B7tlUMByzBhsGPEL3G/oLy6QUFXazAyz4BCKD1d
M9jz/CuZsfiPRasDZBou5nBjTvYArfhrUqQfgxvOIcUklTRAXhSBo3Wx5KqJ/aG9y9oHeCpg7LzI
/Vpxc1IR2/8FQFEkESRmcb05szNtUfSzncvAOs7GEfsLSlPQfmrBn3GrffIjyYqfaDSceXpNgYM/
K9/c1oc0an9g0w1CEOyYI2Ot7vTzqdIbxTB5/QtuT7kZkjrXNkHuHc0XIu21MU9ZIiyyN6UznDiH
xWoxi4QAVTz86GQXsCPiOtoIf7BFYz+dNejYW415QE1ed55S5DJryeT+K3tUNjkF/dlWsN+zq4zL
rfZKEszJ9UDCgKxT0F+Ge1ogaV2FXlz9q1v3AKNScNyJrD8VZoemOhrfHdLkLWaloIBbr5rCkl4p
Agqnq7Tp6ZSTe3zSc4Sd+/O4+2Hcmvp6QyYl8jhPMzhFzUu0QGDLiHfcaGALk8RRG0fklWvScvcj
fzEk1aXwHueyu6bkIoAWDlsXNRkBWv5HUEU7cKgaZee7+FKDZ6gT0C6zmeniftTohGbHH09kOjpb
INue3NHbSls2ygnI3oLuutM3VYKBs5DrF6qFxO09v/BgAMT610ui5QFCd3mQUrn98WCBIBzCOyjp
r2XQBMsUg3jfWDR/3tVlT5AU47Dcf1l+I+qAW5jKv66ovE5WRGcFa39G5FCzWt/YWlHWybX32QF8
8ku7UIoaYel87BpwhRgZ2tTqbFq1JKjrU16nWe1QSSAvjAvrX1adDpbfmJ577J/jMYYSuONi3F+q
u0ypuDCT8f4WXEPiiiQz9Wkavd9GoyDgoxp91yAmFSo1Ve+cVKcWVFdYcbKS1RI3LiKDLtTFfFgz
Rr6CwSEsNP05aTz3SIGvs0xmy9c0+7qOKKGbdMQUB/DPjpgwzHoitkFbFdgW/INru0WkJTNgDjXm
VAo2X6g+CvkSriHOFb6pcb6FortkcN/NP0u9h+3Vj1JL3/REL8GVmUJYkrA4aoj5PF83D3hbBxgv
uapmFvLOq9NNBWLrM8/e73UTNyOeuXVG+xlMjatIPbwJgZXM4t+rUsSzaZQCdLWqN3oDISRdtZd8
N+OLkc9CQ1s4bzr4nkBcjRzEhAuVdIz+8Q8w7gh9jO8Qu6kI6Dz/kuleVj4cajOm97PECPqcB2qD
n7NChVwFYMat1oYk4nnsC6aE+8uzPHZTDACNnZhHBhQX5uUilR0Sr3xPyTvFje1IaLQGFMYFYYUa
08pzm4Xb9WQG+sOcMG6//Sv79U9m2r9YL/dKGNZphsfkMsFUoAa8OhLbcGrK5sKr2+wwgFF4JyOv
Wk8/w3dwMeiqUQNZk0z9042VyCYH5I4q/Xe6S3TR34o67BXjrcBOILogGGxfqxHd/Muh7mig36E2
zTnZAbMMiUU6BdHFq8A8l4qaXoiCgd5lPiNptH4mabwRXMMZ49QZKIRbr4jMoBpdtBBUy+T09iG8
QU7ecPALFmMz6bfILN3x5Y+HOlIWMSuorj1DqTQ3KhoWZqmGjnyofaQicHulPrS2Y0kkHd/g/Hvn
yFDS7FaX63P/czHwqoN2bGP3UfBrbVEjGfDUmehRlgmGbLkrBDHD/spcEskmGiPXtAQ4+WPFAceb
jo6G1KlVc2q2++bn4iLSapYSjPhSEfJFtGzfKoHSusMHnwijnTpR2agn6YngJk5szVZRaHWEzNKm
85GfvLdf0hECsk9eRHLfzPoNkwBAz6oReCnaFTyLi8ABs76uS39ijSAMff1wCeowKLPo2GhL4n65
LkhBx/y9dwZA6tsWBZLz4GZXpLpt+Ryj2zPYU6GsjDCEZci/42wHDkyttJSneIx/jRF6d1ta04ke
j4LdvKfruoM6N74VjvkhOWFeFu+b5HBQW6eJWnfc6Ji+pCjHXAQyVIUDYySZaNSxgGFiqUI4Upsv
30ujWvt2u7jvN9BKdQ+5Is35IiIPKOJqAZflIbuZit64vNs3xRr2MkX493C352epLqoh2RH7PGNm
70TOARPV57mlvLMqBCKY/SWQuxPqZKRUrgSE2jJBNJuad3ERuWV0hvoJcmEn1FMW2DH9SO++HKN7
jhcUuxbquGS7001qcL56JPHbacWBY1pPZ7GIsREiZPJXgnrAhr/uXWO+u1Rp7IDfvcV5xVBc9T6w
tzosO/0o/qIezK7QEtiE659IBZiWDAPl4QbXTnXNLghvUQ5RZzj6yYNUoBNmqOH/OW//pxou2pWe
svOS1mQBsxErFG8uLyNqi3qBQp6FqyTtdYAFMTq1jwSljX+viS8bfBb1qQ04Et1oNMcPcvvsHPf4
C5/3UBdmp8KsIGRB6yKBZ3CZvi/kjIi07/dit1fJCQ9O/XAhiYx8NXHEFh6mFHO6f+TtGgtQ+xYB
igS64c4LfjaZYSmbMPmWX0iDso5PcbtJUuaGVeUC3N+RkkHOyXXpTVOyFbU81aih7yfa3t7Pyr9y
s90StzUydSy+9csUNwRqDj2EoI3C2Ed9QflYQREcyckxs5na7kM3OnmqfQCCCekWP7UNFtuGFzWt
nvJT3e9IG0zBVfz0cWW3ug3ew+nk48WCsLs7UH1zbX3FTqcfDBpRFGnZShGS1xkOWzq98PihEQLs
2AQyQzyZxCQBE29x0BfdLOCEHCFAZtRFPVlp8aLALVPOpK0WRnbJdKJeETnUhS7KT/dZMUjev7Ip
Ifce8b+/Qj1yh1FpMXvP4oJkpnFVdBQ7oyJ4BDKH3/FKaExdp9Eo+rj3Y/CTUT4UxhOwGDiijnhU
V+P1CwtMaEKy/9/K548wWvCw/FHItJoXX3peiLnTTo0sMQJ6ya7k+Kvwl1+2Jzq3f+cOLyTlkBPK
EGjxWQfxWWGUWABPWBCTrR5x15NfO4j2KJw0kklkA++SaB5JosA+SvDaOeGx/OBW2IhZ7+ImX/dt
iAbM2JkToPQTKEjzVY34iU8MZXe2WrbnDOGF8IbeHI3kqm18eLCTI8uzjw5VnmfgYnJBB44yDnhN
G021CY60laVOd54h5HLjDwec5sataktuzCCGq+mKMhqBfEjBIr2FvH9LkXyN/49k0DU9g03MF1WB
4F7b0TjpP1Ocg96rbmCXG0+qmgMphYNHvISLiZQZXQDdO9bLqsUCH5D/Yv7bcCe0ttesnuHDZcUU
Lga6f9fLgjgUsEt9iw93y/2Vh3c+NRh6KZGwXqv8pLEotvu0A0jPuyjZCZcYWjcTaKZwYQY/0uZY
tCnEP1Xdu48TOm+Rr8krPUHGwuhroUXb5kLJaQFUxvT7eO1gWtDx2ATUOR/spcfuEbLI8him4oJs
oaXNuYmNLK00xvFSFHGzm9n/Z0nERe9+hUlXtPue8jwOFdRK7aRKP/WuoWOtmhQaEGPSSXkE/m0o
4aPMoEQGG937DNVybwX/BDY/lUw5a5AcynZ5WrYUekkwRVZqA3iZTQfKPuVy2y9lRjboCGlamH5j
tXabIlqPqyKlAeMAjK569q9x+PPrKQnCDlbTIBOtSxBDrU0zBtXCLYo+qpnmL1ZrlmHQdb3jobgm
5QLI9yAMeSDg38u2fMYz4Jx/wuoih25DmhVA+lXG97e7uLr+WZQPvm8FfjslxxFRLbzIFgEJIvnr
yJ6ER3pRv8K6UkWb8yVpp0yU0+99TNH2rs7DxbLN3uRJmyqQEOApPKRd8Kjw4MEENFTALkTCR6Ci
SdL+T84DBjUK5qYpmkMCEFXoLZ6kn7gxCmhxLyrIlUyWnVotK/c1nfHxow4RNkMXyHppidRDtvj1
BYZLYQCkM4HCXbPpgulHRJA5fNBu+jyFrkf0WJCR3QURI/2rtT40mO7rtVDGpCY+he/nGzNgmp5N
vQ9fTChL5wU5mRBha8R6Szfo0C341xTAGBbsjQgzl2rSfHCSh5+f0ko1CAuLlNcRDoEaO23NPLCR
kw9MGRoNQMBkoA4CmnHsJi1PPCE25devHd7DruBftSHAnZtYcpWh1wXVYHz8ksTCNEhC8AOXj1qq
e43b9pfOE3ASSwCRaD4VA1H2M/oMngLISGgtfTPNMKv7VlPEpoHz9riRZzsKP6u9j0Xv808e10Nd
/A1BLqDNxA/qdY2lGlMBI5KxzK4kPZPUyadxVHk118xzDVHHPzVCp5nW7mjaimyWYaoRYIpigPpB
Uu8f782jp5icrU2yAdAOcWz3LJb2twTGjX1kwSFgB9Ga98t9CArFvzIgCfM9dFKQuu6la2Cmj+U4
k9c4Z8k1pGf3iSQ2kfhnM4P69ZiO3L7Y7uHfUqDyQYZrse3Iqs+nH2j9ajZxFO1kVR1d+NJUuoMm
GAOsyMsqvoBnAw+GTaIND0GsCH9kyomMqzVwiEk5uQ/9luY/RcSZD6jORHuiUSvETfVC33sI5jNT
fdh/1epN843eMqqvVtIFjpDddokNL4CMNYWD2UGmPi2n0zhoT10tMzlcOtxjOZsPorVbxhqmu5k2
td/rVuXHRokvKJGorfHW2pka5kMt38UzxnwbRm3/g7SxFPmqBErXEfmftOLfULspl2eyjsy7fSZO
o3saPEKL1UiNobtjlxnnzkSJAOn25Dav/Y4iWSfNFIvlv/5kFH84wU56dzBSjnNrOWUeWSB/cLVn
gSBmgi5Zvnf7nBiq/HLGACZ1FP8/Cp/+ESaQKVOgQk1jPXOEWJkn6o91DZaoGHeN5TWlGmiVRkPm
SZce5IuNVW43NF2zMn8L04+sAWVm8aG6FSQSwopqCdkPWj1TthTooPAo/JKLKkLDCabLfOflSm0v
w2ctgihLPUvEA+3AM1fdeTW4bAf3ERZHju0BX8HHFxUfwB9/EEVoLtqlalnTMh/npPMHOXbkybWW
QP90jbJzTA/K9PXUPsfW2fGcJNnn+D+c9Dz6j1HZEbDQi0npSFpvgUa+w7tRj51e7pVSDlkiPcGN
2wu7ZL7dqbGvpp2wRrZ3EI+aUTXEOIo/i4F49vVIn+M2xempuNc1XNICNLtX9LURmIGjSAAsGcO4
UZclHVuJaH9FouSz58G/sGDhbbfEVLA113TBTaOJ6Q7hy0dOKq21Zbuo61qeAOhL0a8xU8xu5CJv
N5ngZHh9s+QhW67NT8h0BsohqSm9AUXSBxQZ+rAhPZdzaOfJBScPE4uDnAOefgk9wRmTk/0BPS0M
Sdflh1ICY4Z/Mw0O6fL35weJ+vjZ2cuWtY65FgK6Xy2yP5XbY6qwE4nFJZt4uT7ckRlEj01d+COy
zJjitX3+RDe7zCQotnynwPg+bEhmOLFDq9QOhNbFQ9jbfM24eOSksIf4bgXsdPxJNCjY8jVo3Rc6
XXVyxZHrbWejuTPWePH5Ey+8MzyB+KlnHs4IJ1XhJBAB/EmPGjbdQgFXlr4pqY4jrrWUpL0TlSRr
/M7EJvrehxyRMjVcuNTkReo6YlTYSuzvsD/QYTld++ZeR/VER3gylezsqvZQ19Cm2WS29k3qL4Xt
zfXcd1ZN3OYi1fYru76u3GrwigEsFI0jImEtZQ0murTqRWcWEXeaUT7SMe19jarpEEHxRGAWf0MZ
3maTwA/tUttmIDHtf8jUJNQq//GyD20TpD6P2DeMIm/JmaeHVuu9n2rhLpSrAVQu7SZNiYCLn4Pt
oHCkriohWxZK1vKK3u2PhJYAZKk535C4xydiq5fo3JNlXZif/umgDxg5KLrnJBz6jQOMvnornKDe
6Lyyp5NsE4mXQxT6mLjBdwsYlvfpswOfP9j0+c+ZMwYpF+HLf5bAi1YGaknY2POWO+JYy+/ktqDJ
MytfvwfNHePql0okSc8RUxqmmujHtNHOQHp+EAJYHkOwB8SeStoFWpG1CkxQGBtmedC0xdW+/+08
MIC14LLpW15lmMvJMkRZxRfFPK/G6baYALRDOnkZR46bsiOtbllsVxE33EvMBOtHkpWcnaCn+j12
+/8JSqigWmlb7RX1N+EXa8bYIDLTDIDzkIvTPmJfKJNT0Pf0pYT47tOxqFKogSJKWKlYSmv3Xacf
B8CTX/6IeAHz0go7GurdUkvWGyNUv6LGyaSmdQkHeHHG8HeqkUsUkVpXz93M+x6DV0OfhlKB2REC
c/X8h6wYhBzW5rtUdYAUpzdpZePOm3iYat6hYHHFgyh2evbdW9kG80y+ZSsbucF+k9Km0BPYT/1y
Cgwg5m7z5+U7VHBDv4pTx4nfejJmNyV3NLpSdSC5lupyLAY4T17JKMoNt1j52HsXCOHHlRc2gO05
L7TTk8l/AQdXCoK8m55CGCuVq+5DSz2p6SkbCZyJaNjIMOotI2+VfeAbcLScKW2LrhMSyOB6uWXl
9n9awbXrTQGOdv7rnyiVgytnNHfCR6KlNqccb1T8pma41tnJvKTvRVQcDUOA6c9C8+mlwBX0qyUz
8yvRWnXF+sjZQ6ElkoGpj0j4nsUFbExZo8VxGPYbLcgHJ6qfDcmSum4fha2B8nSjz4+G0BlgTSVP
jCDKuq5p4gMzcSEobIfeXv9Rj+XsdYxgbQY9WpYF1jYJ6eFAFm6nrCm0U6gZ7vcl5nxmNRKgBM/w
PJmZo/SUWMOKN6z1GmAiUAriLeEOVjo2sI/ooqOELZJUi9VRMOdbrOQe09+kkXrcFLcuhBDm0ufN
4tsUJyIDfgFh3mo0Eoto0fCr1QWmhz2fJwYXzPXXJjAqvrXH21ANRnBzsGeepaQqhyEs/NIurNL4
Bn5VBoBsA9K6bZym9vm+EN0Ec0jkCAvqbqlFSZXRyDn+aaBj1IxZOzLNi0Z3jIfA03v0WmmY5nLO
O2m3ZIG6qW5YxGrhTdFfuTYB/gcRclhD0W96NTYpyFpm5qwByOmAKwr0GcLHKtSDuditSOlIlkY3
eXlz1aRdrxioNKJacAE80+aDc8fLGKGiSXMdftrm+4uafgW52MFdKCqyIUa6UNe5AdtKIGU5SRiV
Kc05S21X7VMhDxQeYsv1+XhjW6w0XB7DeGUprYvIlLIRo2S10pVZe5eSrrb7ndNGbtfW0+jszse1
R2JIGuDB0n0hpDrJoCKGE+Spzlmc+tKFJUQZdSI/lmd8f1NJtJdw4IfPYDnnHGEwOW7HvSU3w//z
NshlKjHJf30ipVY5KJjMewR83ObuRTrKJN/UO9f+HgMb3/E1rksv2QDocty+XQNoM/mpPWfhkORY
RQo+rYaXWsBLjOYMuOio7aK0f8EiUIjYAhzJlb8pVRhLljXwf3bT2xp+d2r5OvX3p0STj9S0AYel
LD1PKoI/8WC3rGFWyzt5JfSD343c102V1cTs5LCfNQbEQ7Nno1VF0sUueeIzi0uNtrMBluCcgBiS
jm1aBHsRAG5cfbYjo/A8TP3Sq3VINorVYtd7yQ5ZJAtUBLIYm9TLj7rRydjwSPZtCrmFd7+WXhgh
lu+W8q5nZ/i5hW7MmsGDwshben2MQrdR9FM0iOzB5/l9eCG9DVNxpu/5cNsygmxC4pKhRvLrf+dQ
AaKb5osryseXAzZjU6GMX+D0TrmA1wYSeMRCI84A72d0ZF08M7/54vMb4AyCJLBB+tfgiNhqCWSW
Rx90mLHsaCdBZOn4yb9k/5xMcBcsvKSLmjAUxgMALyUbTUSYefW7b10q6oFNG/aq5VTBNIHD6gRw
EUj/0Wl0Sdg75zEFqnZ/QQUrmhOcxIfS7nG+FHqWZOM+/F/Ej2FZOt7JU7Qonjo79145ym3pAoKd
JrIhBOVMJNJEYg6jao32EwHuPaUr3hQgcvoWVaePW+45n4h+AKieTOU3fUqoihKawtJHQQha+Fmf
1e+inkykl+kMl0QAMXA5GRbZmETwJj2qddMI8/oFS3YjCC9VsBy747ltkxmkTdpijgNtDJVrBXeH
kAnQvSaBuOago0ZTKZE8dRyxXuNFzv4uPLNnuC+meWPKWkO5taEKfRkGnhKxvt4tzpDyFGgacwdb
YV21oHZSuK9aE2JV9z/QcMtAENsYR+Y2kvohHzyfP0RbNlhp+YSE8FdN6Ns4L0RApIVFu/A2q0IC
yxSsx+dfSQZjkF2DhnoVQITUV+zkx5KH5dEfnJaJ/XEEHIklSlBaBLISAvplnj7dSXzQBgT371LV
OleJnCfjeneTjYpgz2A8aqLCU9WpUGcu0FPo9ZJ5SATab5N3i/wwO6vRE8Tw5mvVQdKEDrHwwiym
0aHopP0cnqzeARchpRdE+M8Y5BEjF70tXDv2P55Vxq2FLlKpITteXw66SYfzYYj1C7gCXvLK9QKB
Gr6BEooJX9x/LFVQxdtHeE2bx6Fm/D8IURNAG95IHe63+EmSDBF55WS1qK3uYbOseK/nqi6s8EjV
erFlHKqY5HVKYO4THLNAOzkXNx81jxGjxN/peoGbgEc0hHzPxZ4W7ykQAiMrb74M/0eJV+LPS+hR
JLNPqpt1TKlW13ZblNOIU4ojr1cHNVQ8xfwcUNMyyM4uXcEb9ogHrfGUFsszxDkoJaBzO9YmK5Qd
5qf3bzpQrRfrHFLUV8i2bRvSKsceQVjVOdcIr2pAzMSNA0u6p7tB8KJagHZzUPQkD7b+c1Y6ExKS
fi4/i+2GdWczwdnONHOtqfmyBXQYv2x+J5ZepXqfRkZ9VAUgdSY5tPAjqs+DWcYDxXSO5cWx8H/y
XAZU4LdwN3IYQmF9eGEN01NLxf2d71UlRBy5WFoEFk3vXC197FtMdCJG3Q612Hgc31xO+8krhOZz
j9tGcYRn2IXXNJ6UVXnXM69XOV6r6VYXFPTm21jsJRyFFKjDD8AXlberkgBNQeghKzyA7o5Pcj09
5nbl806TWyyKR3xhqGO5gAHU++uIAom0ERzafMF8jvXBAKWrAR0XN0qwTx1f2a/hNvjZo4uxlaYo
coAV3BIEFjFsR89tlkPK/GHVhttI722czV+qUBE0B61WdePITFKpNmVxj+XOv9DqVZToV5wId94O
b95GAQuCDaGVXWW5q1sCH6a0/K7PTng2afPqjxlCZH7QTmVPWmvIgzdLfx7WVfvdy3KkGHp+tX0w
CRcbOkWARdY66nuR4fULmztCfuRxEZYEB+xEzN9bKH4mImDCMYft86hBOr5v6xydxJO1Vt4Pk6aE
Rd91mjRPqRdeZoS6lUoa4VqXV0h0GTTvSOsNIn3T4d7y6ZewJMccbiupnzz3I4MaIdc1il88f5YN
uST9waGYDFTZSbnGU/90hjX/F4sGWMI1F97j+RnTfUpgtvFMQ/uU7kYp5WFIiDAQB3+NFwzTzEvb
NOEiPbHvSgg+QT/295/0vwCekYhTj6pfRsEiCDMzINkGW7oCKk8ASYHvlrjBqTTOCNHQRtRGyd+6
71pK3Ekf8flRIakA2pG5Jsmlz0GTISC3fbKhyK3wsXfQxfQzYlBvzmu+RDAFisaYukvoUIKG2FPx
QP+i4GKBEfy4vIaL16nE+LBqQ45hzRpzLOy3khl8z+6aNyYUuk5oWGiMAnsxumGUq6g8wJYl1Q3H
8qgvswECxwEO3I6OEG5/WU5beMCNRVa20QLHlZnHHErcQpfRTcVatTqfDw9ize3KKXBRQJr8KY6i
YbOLR8zwQd2T1T53MtcKeQf+YyXFXfJtdlkSX6WUU19YHmArnv7Tk1LV7mNg58jtJxoggZU3UeOz
R4ksrG8ULhxrstOMsggaaI73H8CLpDJAYEBa2hTCncYeVdaSabBrzwQmjAl7fJwINfqn7xcg61UP
uVPpkk/mn5aENLzsQsR2X70M5KhiICNpOZBO/o5lShTaauFvNSFN0P8FdV2e2zhh6MuA6VlWzGuw
ppTv2g5r2EaIMBiUj9OOJz9Rg8Rk63hyl+e00vmWjgp9U+ulWBQnUWn/8n+kGNJVEHwjieP1ecni
Na+1Buq+YfUMiPe5786GYfHvpeulmemFdwCkrwUO6wYEB5aqPwThnAZYdt6lR6muX822x87i8PqI
xgNF4d+fuEYzkTbg9KZsMkx5ILUEhxm9UxRd40ARYUrIE1i2CgTzynrMMGRHO3hGNqyG6sXlx+lU
IDu+CidmsxrdTTPPq8kGWsZWZi/5ofPjhBb++vJFJ9h1CzK557ZUYVQPoZdcUNj/BJSU4JVTkp7f
kTynW6X08SAZmt8wLJW1ZVk5prKtvWFp14zBDHSCQ0Xu5CmkjH26BeBXfx12Wne9tWoEkuKNVtQw
I7tntWDUKlLHrsN+AOIZqLmgAUQeGnXvXbouhJwRXi/mdG+uxH/Rn1LGySVKS4QVL+Z2bs5Eore6
4rvd12b7OpD6ySH1l8MknaLccJ/ApVZeadmoWuQ/6azlMYAzXlGAjfkJw9Wj8Ci6xkHqr6iem8u8
p+554nHCik22Yr3Js/knKk7dTqA23WBdGShK+kBE1wVy6dYrC14JwT7GqiR6qF0664qYdlZs8lJJ
tcC4v95PyGie7X7pFgiyOC8AoppjHKMGzpkFQIw5dEZiRTSM577HVUJE8/rYIgYhF58Vw+GjfjKq
l4rNAHw2Z1s7v/zM6YyhLIflsGZ9fjcFZoc9mUOKJQOs1ngMGpujEqWzzINxIgpCQ2LUFLIgMWhl
kORCFqSv8gIwbD5o+NNqwnSXNP9OOFch9o2iqqXPCPiVNcTNibqEPgSDWHvirNHPOgtso1Ip2NZw
ejgvyfVze40cj7S+ANi17qjXHmnF2UTMX15nPkTVaESPRg9RmX9mioZACrD6EKFOo54Nay9lH6ow
mN2II58Hg0EKFEEbRk8nGboIsqiEdu9++8oRl8mbfrIi9g+KlJhRgm0Kxk/XRC/4quHvv3oXpoxB
aFUqnFtvbon7YiK/vWkKwLFQgsDMe3IfkWLLUHhvd5p6yNgzHA76F6Q45ZsEEnsbNbUZukyQVfGI
J5/JOOYPwWv6ceftLlA+jzDNeXKx8EixhPj3MaHFAufXtAlH97zr/1SDNhyMzRzRGrRurY1gUd2W
wlPhEX04rnJyYPzaQUAOBCyEjLCaTfdrIfQ9Kx8Ju4MAWKTKyh/wqnkc99zvZzk6G2eA9TzP1TYA
4jxQJLe77S+B1NVooWaVpgMGhmwLoFgTVgf8FFtuvZi2DOYF31AP/c/T9SP81wOgwhjjjZ0ULMUV
Y/PDNWyejoBNRpVrakxGttCfvdRKNsiTnarx8PzBELsorJW2DTRFsGG9y95nugInf8+0rOlNXHLz
q+XzkgPLH+Y8EYj4Brw8nTut1091c84sqIDVX8P1dm+hlMdXUMg9p9a23b1dlpZoPwv63jZ2IBrw
uy7VSDes3TmMykJUBJL91Qpy5r2Gl9+rrwPxzlbp4IxtFZINzDM7HhqDmx8ThlfYZb8VUU3hnC8n
IKpwsLe8qBuGKJardIW1t0Lc4lXEw4RZebbrUIJ/VoQpZnAywO73Pk+jl4bOmQosMB+nukwRCa1I
emAtrqeOcILba+ootK7fp2P/kfi2Z7rZomjmlATCgrlM9/TUpokg5E4/clElAgCF9T6YRCSLRH2K
Jr2QXIGvwMSXmWEa12tX5hrG/MQPyb0j319b4g+F3p8+0xSK9QQwnOkKZ6oUkspQo+QPz4Gq0L0a
4tsRjHlTCpZTmHC3Vxf1eUzXLwiGIBEm8uSr/Os9tOL9gqE3BaSe1SbM94NppwlBgjGa9MqWEPQ1
m6M6vlf51rnexEOYgA0I9ZMLM0oV8XN5p0whwh7BINR7xi7yXoNdiwxhzWQEBU93c9oPpNnwl5GL
8GSz313IcFWHDqZR1Q+J22PoPcNrhzVt6nenBaSKLa0KSEsecge3jOiLOP871x8YOySXJDbKuJCf
Di/TF2lCnWEKXhfr7sJlHrFULljX6OvBmT/TMJDMSyKRYZsVUAWyirkWgn21/8oX5wMTRoL21gMW
wkRXIMtbfUGHjjZxick8yFxwxhD1JKbo8Zv6qTYMarnLTSfyDWoMo462Sj7UrWltozXxHd1CD2hd
Q8lrMH4Ks4CjMuuPMn06MXe3X4g2JrZkzz88nIIq3Z9BkX8MILjEzCrLwYNz1hvfuOQ2lAxN08Jd
iux/BJDBKyr2wC1LoQ4Y7UJcYjn7+bCsf5fnleNvNw8gfgzznggrcoATN/fzB9hIeZMYpl+XrFFw
9OCThoIu1EyYoNzM0At75i3GtGOCJWkBdS5lpR6GgxVfKZzQt8XiKeWG1X2gJmLHPgRItJosShI/
avP9s5DPMdaxMUlrSqmshA0pcP0rR2sRPGgMjoajLvUjJ+/A1TSOHSJumpjvXZG+YEHm5/mM6uOA
KqRZY0x59gE23wa3gd8FZOn5WtQoX4Cq0nc8SunMpD6h1cd9C8+pJX1R0xCCdthyK78daSu0dft9
2loLSmA6ZcRFw0rFSxmYQgHVfxecy93xQhYLVnO9Z4hgMEHhEZBp7gV0Wh335gPuoeE8BaGOFU1i
6a36ezHwJtMKULRW6/LrPQTAwS1F6EfW0oDn50bGir4j+rOT9lJRUQ8Xn/O5eF4YelBAewpdf9e/
SsOJuWnlE81s5SallAvGVh+c+C2LckqdJbCo1jxU0QSUzaCPMvTVChNgIfPW1A8wAPfSBSOXFKDO
atQnrT/Q9awX00VE7qWfgV1BmVH8MSzTFPE3tmQRB9dDSKj4nU7c/CRE1pXZjy6sEX8k9GPfdWOT
6SBX1lLyBweh1ktgcNwHS8eXzrXfTdUp8x+BQZFKG1GR/WlIEeEFmLELeVEAjgHkFISndMiNO+I9
007q9lybukLpwGmWsL56lhKkmPVVZvUFPBpgcJoKn5FUpoOXKlvBmvrzOD/5yIs+/3hjAs+sqo4U
e81523/1T/PQ9RGrDLTyXnnSRWoqlvjXFPhhEhMIK4dhvcccKSnKI0ubNFC0HqXWkf1VN4rFzFsd
fondImd+OO8VVLnt4oVkyRAenztbhJV0T3OC7sTB03gnBHZxyonEeQX5QItewzObp/DyTvimCavR
5nb3oBooSWNm7VauzqL7Zzjj2hth7dVNbSEmbmU5HeNrRZlmV42HudyWahl4OfGhVcj1MRBdYLuG
M1tFPCu5dQRtOLOUP33JSMXT2OmY5tiPAd5F+4Q3xMmoDiRwk4L8Ln89XcHHiXdDlLHuu915bSuo
D5xfnix4+icftVKOuxaOU7pY3oQmgkHJ4ZtkZfslh2vR+65TCHIHK57yo6imd6ku7oC5hPajfYeO
bjKPhy0SiLCVTbqqKnGGoEYPdu4XorG/RaIp55Wljol95VTsST1qZguL3600k7mW7JQIIvVlVbry
HViulSN8TU9R6MZ6BN90fdKznkgjdmelsGl2zXioajULwdZ/G1LdI/EySRYqpkP+slVeqDZHcHvI
VQNATx0kyizKeQmPetnNrsDEWpogStY5oneKxwTb/8C2+nVFmFsuFvSp9RThyVEZwPCxsOeOXKSV
Aranaz92EXoKKfhHR3Smfh2g6zVuykW9QX6GjdmfV9PMYFSbKlOD992Kuqq3143C/Tn+rcoWnmoC
ziF6Xu3vve8iG9ofuA/Ly5FUCTP042vYcXJs/132yAtyGh5fjF+QueKDrYUjR7sjKgDVGpkvLwBa
W9WWl+Aflf8j2+h88Z2mt3z4WSslwdJeAhhlzJ8IWDGGYNUk3rIX645YsAopstS+p01mHPdLmtIn
2H+7uJxRDNr1+bmZagpOFGAOMkMcvLs5OPQ43ljuYUoVovfyNu5al0i6OZxIb4Nc01SfbKmh4Zio
PcXN+fEJUVmPfqQ20p/oIvcSWOV479fW9p5Aihdl5SzH82zjMTM2nJ2S1QTEhfINNMgAE9Tbb5nG
3mR5mYDAHEO2plqlucjZCkYfKpAQPAsHpeSq0QmMRSDTYVTbAAOZ4MGQDxSBj6lrBROyMTdWbFvy
nz+4vbOskm22S6x31uk2g+jCjNPRxGAqsXVKNg9OB6uOCdnvqoIQpRxu578kOkCi4I+CwZoQt0In
Hj6DjjVRe0ZoJA2IWW6o0vIQId+Zym7LTnykmVeq+GT89KUVMTSbDWqevjA/jATq//Bov0y9kOxd
8KQfq//ZmNgqSC1/RXBYatAohGV8RWE+B5VDcU+GorQOxTCpXETErPDNF274s12/EYMaLFcPDbNx
7ysnj0Kw1PoAPaWpmvDi1IH5HlR0VcaXO/Y7Ys/wU30XhkAPmUGKwYuNv7AqCytz2z9iVI7qJHgT
yJMeXVkZKFQkI33vk8K+IpwmgrvjVJcnyBHjCQcAyBWPFV+kAjykalUCe8vFdyBEPRnFKE5Tfe6/
XyAWHe6HOxLYCYppizBpIWYbpDgLT35uUfCdgQqIL/rmXBa00a4wFm9wOeIVrdc/9HVaCwckiGeW
C5SsKIooIcsrOq+Kk/4jb3dSGeNlChDeienN64tWS3/cBe3n2VwW/ydUas8wU7cpZSLrAZxh8+5z
9xs/Y4OcbxKJVqu2ZTu2Gh6O7VRJVrucyaYeJz8TGRK5IxBSZdYCI6qCHa3Th70vpRE4Q7t0UF4+
mmC4ZDnab9Qb8xXSTQYaeMX2wDJ0E2uroih5DLW0ZmIcgVFJJivCgRLJ0jV++7VbUi1ZsSSLluiF
wvyefkcqkaWBkg2lDdD7Htul3fP/YCGcGf8+OZpd+DEMzSVukdNjc6RgVzV1IgiqEMX4Ebp0cS5C
k+z4ZfSh4QltdYr2nMFx2DaVIzdiZbk3EBdT2KtSPII2FcDDAUMA53BuCgNfRX8P6BVH2j/zzaEt
hBjaL4urW5IAAJ0KUXXk8SKB4WRSyrjHpt3Pasa9pi899XyGRssdHsfa0M6KuGEc1FN0K/k7DMtK
Xf/KtZ0pINCjL47JZpvfhONo3QXGF4GjfwFAR7Y+VW7F56vxK1tbWSCY3VDfyqq98yPPq8N3wIDK
/7VKC/aYLULHGAA+CDHDC5LcS250yi+7mz9LW7OAeeD3ZT2MwYFlDAitA9DXqYHvmIoWA2LvY5H4
Zp58l54WaWk+wycn4zPZiXarMuNeWnWCQl8XyrP15J6EhH6rBeV1jsG/+5u4eVlFVysk1WmHStYD
LwGqZJ2PCfPW42uK6fJhvGgfiOpm052seHR+h2xWOjMfqPxNREY0gDak08izB1yUTxEV8jOWh3Gn
5bUJBp8QyM+4hosDuk6iKsy/fm428osJHFR/NurCA70tNAg/x3JTVJr515IvsNY0qvnHXYhUGRaM
0Oz5FLg6WN19miQxm22ET4+R7Y4pLmDEOWAqeHL81M6RulyO+Fwgv9Dor2Fjcrh9PQWf1m3uNQvS
kwPeroab6hrpE6Fh128boRUoQYuRnSjWgm/2cTjlDLGopy/F06dk8gDVB2IwI4zTA7m+03xGSzfV
zp6RbojQIO/KOJX7euiEK3YZL61+rLMwCbyETwoj7s10lwENd/vIdEqS0x3/oPQI9xnr8bUePDSw
JLYY/4dl2NSjjdXU7J+keqxqS/NUbis3lTO53SxfsfhmKPdPhOj9Mi8+TfaSS+ogivCHrBUJfr8u
tCTrN+fQ2cIPeAhTOx7QgsSYpWJe7GVVvaHg85Bv1x+xELFYcwdzKHGiLkYmQlzjgqK1BYOpQzO7
wJ2wDpvZsrxoKnZi+rjR4FiRlsIg0lnlkpOAc8vQ5/Tw6SDz3uosO223IdA6sQabfE6ASnqMJye1
9HfsiH2m/IxPZQsWelqAKrSoZrZ9Av2E+JueZCGRs8PVDEwyXD/Ak/B1JiqSu26cWyKYehW75atq
2o7J6xpKzrjqiMSXz2gqANHAuxNbcsgy2B1p2t35GQP2YMuvLFAb4uZhJEuA8Hmi1KoI81c73dV5
KQIvyHEdgouUzz3GXwo5+lHBNxatlzBeifwnMszr0Pj52lIcQnBmZ+uJ5DLSbfPi123r1nJwL4fG
5R5tsPOBCUJcKrJpT//N92PP9pw5stQ4AZWdLcVzTkrTZot5MwFrlQD9xlktyFXEt4NFQai2+qRC
0McKVieNF3j8JBbQk3gVO/UCRxUJjiBDGj+sy+3nAby6Uh8oYih5M3Ly9scztsNmtCkS0bJdfGuJ
SUaF8bbhW4IymnhFLoKYbjKXVi2OHQwOoT/eOEK04UNzkjQlj9MZJZrkyS0wO+ZtbKkrzdzkdXsX
FjNMCXOyKfBuxZBxpRtuwGd05OFdhvklZBxBGglPtJHCklKlLB47dYuHmqsdSCxNc9ySD8Tl4ozR
tRGDnMarC/Ku3Wo5nC2y/ffjpOa1WCMSCeqsfBwpUQp5b3dUVRj1g1Xlodwst9PSNvPC0bZgKjid
qXfgNlnoDgsWw4FYPw5TD7OEJMV0dCxEil2T1I/L95HsRsaGslE3s+MSvfPK4ZlZurGrgnL5vfu/
NGhHLYKtBFvUZGN8mqAVyZw6RHePCZvX+UkPi60xEJX1ej1NbyuwHNg1PVZw8/Yq4cN/k0RAw7AH
oyUOKr0DoG/H8z9qmPe5lWLW3FhTPbAfaaQ3L9dopQLrH8JUtbFrcdtInWaCdQV/TBeSSStQuG6t
PEj9P6/heu7Ogaeh+UIUDebK1rOsus6+7QzRS9nBRgDdV18y4w4mC1bp3eHmQKq8JDS6UslBk72s
5FSJEs0okYADbTpXiQzbgDlua6H2js+2D1rJmWh5jlnGAxSWo1DCbwMeCNiHGl/NDylH3wPjuFGm
JfWtyJmIBYX3Mw6sLCar5n1dp+S06veCOhic/sn/8vWRSVdr32/r1pcExLM3dejdUcfr9Jma+fjs
nqFQNFbIPhYpL0y8RVlhdKCZb8hUI25hepMYu/ab0hvjRk/hDU9x5q3rnFOdexiriwwTVEy/zz3i
0wSwqEvHFhxYqLtKlKZopVKd2kVSzyNfR8LXTA0zUAtXZCrbx+z4Tb5EOqLih6dOSZ2BE9PDm8ux
B2NIkMgasrdou+04WUwywKPNWEqGnLqaTng7qI6YX3ifxpeKzIRBw90ycuZScZ+Qj/yVI856Js1t
foHi7CuApuAWu+a9jh4eXcg5tK1JS3r2FZH6vyMYeG17GraMK+DFoVGBlOGEI2jCTJW0F8E1Aeo1
TyApTndFhpHS259ElGfvwg6FP0Bmvt7tqjlJnce+UvSH9q4laVLOSLpSX0KH9TF4B589ygVcw1nK
rhuN+up8I44ZF+G9SsiPRwRtupsSrZGYh5G9EXKEzmTul+hStz/bY33MlWppWkJriElJoOzBCMAd
ovnfaXmGOGnTqE7Nar/uPLcVCQ6m/ayjfXhAkV/QWqvaYVrMZb49Cnb3gPQp/nm0Ptq5jaeGS1ts
K5BoPxKslHBfcRaOBx+JprhwL51EvwYC9ZMVIRvEM6vK7RNgwk7n+jkxpYqgarWAF9KwZGaZ36AB
ecQtuvo/cd80mxRO+UXc4B4yeAIZaxZU88snFT3UTfiSSzBYYRGZcdMPGvPS28zM1BMgKewGK7D7
qwHOl+66QX6gVzEpHEEXmHRcx4MQ6/p+PmAdzNBpB4EGjkd0RDlOYQ+myCebn5ryysgQIxRtAMqS
VPvjctfrWI2qktR8csLTbNvKUbctac9d08HBbwYP4wm2E8AYLDbUR/wo93+jZ4JFrr2kzTSFyP6H
pfgGTKHezEcjXhYGq6Hp+QrYg/YCHpcgCevsd7cjs6HwDWb6PPzStvecO+h4/XRL34ksdnxOFKHM
92Wd19cUtCJ/3GI1J4zQ8+rGTdZL4bibxGAJeiMeWSe+KZHh5eeHA15ws2DHmbxj1iQ4qtFNDURN
wvHd4CRFJlyqXJutL3B0+XQnSrq9ZMFMPRqMGyr0Kpuz/wxdbGlPStQvOhzXJJAlJZMYmteLCI9a
ASa9g2s029AQhAjOgAIZ0EVJwobrbCWDCehramr/hY7fy9y9JZpdv6YQhzPkn9zNo7e2dCE4pDAQ
ChS6MDBvkZcOgNq7nkP6bg8ovHc/9I3Ln7ZrNhFkNzLdHas4szN6HsleRJZ8GIUkhL++lTt1HKzd
6dhwfzokzMsrr3AD3NIj3ERdIzqeMi6L8niDbXk8ChWp1zFdyF73mSgLKRqoxBExRE2MQen0SIS1
ZN51d8o+90hMYZ0XMNUPMmo/21ytAK7n+S02CJZNnRyUp/HR+6MsAAz1KIX9GTHt8IO0TTNRHCUm
6lGwV1VPJxPnA7oIDQEdBDxb3zFuCa0DYYFDo9TqrZoWtKm2cltQCB01ELN2pGUztMAy8FzVHTHz
xd8j98c2mmtwpnd0+J24eQ9pPpYAKwDSFK9IlYulPbPxyYUpaG7pXdKzi3dHOBNPCBmTDIkVKPUC
KvTuFzwBhvl/t/eOoRD78+FK0lGPprXxVP/C2U1lho129g+jGCB30CnUHL26rhCNuYrEJTyRi6xf
7QHymvyceGap73np9XoxsH2U6xjgWaaZPVbgd753JdTotbDYn3KcK4edg6Zf63w6llJsnRQnkv6Z
IfdSk1sHZrot2nAQsAMGl0DTj6TzZD/vvvSR7WGzf+/sRk1Xh8QwnAepBkrP+HpEWN8bgBBHrmrJ
lbT2upkSSAqT3s+FDQYErhpvrox5Bt9IC/Ua5Uid48DXhwN7X5pA4ZfnUHNsOzlQf5xDgyobkbB0
Q7Bfz2t7C/8p5cwL8lR/JDtXYrEQ2YLZ7BXljy7MfUw0GgBk5ZEGY4+XeuUwKLZWMg2W+T/WoLgD
Vsf/a84YXA/Xd3xH9CdmXGUAEl2E/RrSA4ZZsqDaeithHvUsXlJEIQepIUGAgiWN3iA9YhS7kRoj
jESLItxwdTCJfyoTrU8AhLqzybLpR4JQP4hSx62OyruS3KVRsbadb3KzO4BWT4n5RdrB33MQ3fm1
8L/SUiArT/KXQD9GKNB/frpByJxWe2HbMjvxZ4TVhrV/dPqjwptGueZlduwrkGwr6Gz3P5ezCv6X
tkYkhyJhgk6c5chMZqz+Su3N+NzL6DaZWTb2R9Fz+u5Bszvc60HrkQxLQbuwimUyvkkRS/Swy3KL
6nsQcLUIqRwAJE98cjkBZu3I1mjwjlxWm60DPu+op0WOYzbq9XmUcqKNI3OTmD7Bam5geaQqdpTw
jtgrwI3porZj7g7wug6qnJYX+ib6iCuzFroqUxlRnVrvKEl97Uv3UGpO4j0ZyFKEfYo6+sDdWcD3
AHFlSiYVwMCnlYEKsu5IqOUc+KL2UgCMSx4cMn4cWDBOBEipQBgMbyotYLkOvfRGr44toPrkQiQg
Ryf700KxNM535uPqwkwhqGyOWLxMWMSzOTzmRviyxQAkNoN4m0INRRNTi2FqTOl+ykhnsZ5ujSHz
CP/0kbcIsY/e6MgchZV05NSV72gmmJxop64PP0vtBU+B/9icbFEgXAYGHKUkWL0ciuNcZIxp4H0K
CJMIpwIXFfHD3cITUeebCU3dLhXoYiCoWOu1agatJU7JjrRK5Xv9RdDs/WQOe4XNm7ZjkvlLOeA3
NEbJmHSE2ZEvry86aBRjF7BEvFy06tD4Id32QKrb4lts8+AK3Z2b5S7S5wbiVL1Kt52kMSBFz+fT
fS/qOffI6uU0X1lfHOd5i6NhrW5xlwu1x9NYBaY2y4QAw7WN3zlsDESQkZy4L9YCAjUPCQ0Fqi2e
SWHhUG3KhNRhyKLfdtTOqbeZlflOHqMXSJlFGf86uDBXs9FCc4kZgpSakN3IAOAMM4CW86BNdvNW
cmDKUdGd1DZX42/rVgEfh8pAQqo8+jQDB3O+iTm1pppzvvq/sh2+yma70Bo1U34ASbnPmBGw1vCa
K/nOQKB2eH83GOE1ENAAgZhevbtsiIBdMc7k4DkVQTBWAsv9WGpErNymFXxdmYGb/naAXXEELbGF
aR2s60yI0H9eaRtTjBF0S2S81TNbtBgB8Quwdr4jGmiLSLTYWD4CB7wFHFjpemXk8qrv6fGAldtO
cBrKTNVF8IuRPHBJXy138VHgWlnHV7gPDK8OTAhPgR6EucjIlBTrBz6uE68sUPg86rve4q/HqdqM
55Xur0oRaGXjSHz0zpB3PrzynjK8bx+n6E/Xk0Ha/XD+I484V65NKULqc6mzndX4gaI/zXZmdr1y
ikA1l2OR9zQ83wFLn2o/MFmNyqY24wAGqoizTOLctMfRqQyDLrWqeokkh8/wXsdVhC+X6Ix6WHJI
Uwy59EvG06RKx+9HDmyYUhGvr+vlOdKgYPcZtGP/qVFsnKlAFhR5Li4IbzBfG2G+u/HJFwEWOL6C
Dj6Qt3RZteC6q3zc50BVt5Bs4gP6fDElgdcbPiOoyiGX4oRnDB9ieQr+Nc3P/U0KbE3Kz38TTEp8
rSF2REDkK0GylpVwe1Fy0JOnJMeipQBl9EqWQFyG76YQMdQekvO2rJ/YL0V+T6Htm3x5V5VJewhF
2D3xh1jV9TxbxUp13oP9qaZtqw4KJEAVkUUB1fWnSPMQ0y9WlEJIj5TBNDY6/IsccoPg6IT8FTt/
2/CtTe6kJKrZpFxEQARs6uca5rzoMqq/EkZ1BVV4yfPwlfge0WWn72Qh2LC/VvYNXc/54aRHqQLD
J/zn5LngBjtIsVnBKWqykgqf0+PpnCRc5tdHWIz7iBKm3NAFiP9dxcOBT1DncI1CjMaiEyrtVFBT
iuV5RXoYwm/RlXGsX65sdhm7Texd9mfxRDRiTd44HZF7PmjONyL7YeTW6ZnJhH9WWiJFu6b6u0vi
hEgY7HWqGJ6wgG7SultNBCzCaJH6SREm4NhPOQGAc9U4lBpaMK664OF5PIwnING9iXvgex4gnEVv
4qmsf9DqKp86qx8ozxQ0EE+kiDICFL1JdUNiebtyLgXIKskhEG+g88EA9QQIuQ1Lhpce3bk8Sws3
oyBRPMWcLHj/e2/ehX0PBXk/V7aYUxrWkQkkefYpdBe5qbFrSbwmRvUr15k7VdGFXkNOQ5w7l/ft
zeSh3kr8kck3RpFXwQz0dgs8c9tpVw2LwRN2qsAdxNN256ddQuNmWBk6lNwZHZ59gC4ESzcMAniY
egChF080OjzYTuK5mqqT/N0NF+I0WvetLONb8AkTbp0GZbb7ftWOVqYEA0JaM1YQTZX0S/F/EXRy
DGfui7zS89BtGDMPI7aA0dbMuHCx5I1hcKlD7N4HqHKqR9BaGAOM8gF4L9WDwJZufFju4PLOjtPO
l1DHdWw9Q4kQFfkRdEbX1Hie2o+Zn8bB/QbgwCf/dic/uXeFAc+fL6AU6JlkSMjTHDowRdOjOlrd
xvxBEDK12VMDJumwWHLRgPDGoPLJComyHEzt2s+xdKLZzyBsCnNsIFQNdOyDKiMLVjAWX0VkgxmH
KcKX7L+4Tj49fwKKs4e11Yrkb1f2Sej5ns6XgQfnybhcpo3hXfN7ZukhNeN+P1JPYX/Io6lnhfTy
5a/kilijlM4yKrv39ykNbFtbUmp3pphH7AkCgt1BZBcntHAKrmEPpbrDVC9RXjQFpnyekWxNeWrJ
OCYfyfwkPAWp3/dC4zpHH3F36PBN+53VXe/Ii3UzaHEFqqKDv4MoUCVzGGTEuBSHYaZI0ORFlIe4
LABspzoV/VWvYNpw7SxjiY4l2SzwnLdulvEWYml4dFDunTVHjVv5pjHTmUv9ZKL006y5Btvpb/2S
S5H8HuE6VEiZ9eeT3aF6b790Treec1Zem9rRmUQnicLshE9hIvA+QaBBAK4GLj9XGIQvtWohgK9W
rTZ3sgRB7tsxRFiLDMHIp25RQ9OLmKkdysd4RhbRC8DoM+mZ6w1PFF2Js88koFelKxaDldc98j8e
kTUCEA3v9qm5KkB1W39fhZ7lPRP2lKG/x5l4+ddNzG26KOPAb4eJphJJvdzgSZth6g6/e6o01dkX
TYzuhgb/fPdCKQaz68oSJcKRHOJ94VOSpe3FicSJA2OMD5Z14+brv8Hx/oa+bGPszHwa8fiZj4qY
ehnJsPZSyOCZ/rsAfp/yY0WDEdWa/hrK6Zm56tP+XlET7SPnXvoDoovJ027aVCPkeb0tbnT0ojoX
+guaodIZbWEooHGyKlzjL9u/u2disxyFIcUkAxnWMecOPopJGN5+bGisstthsVc5B8GOdgbhsVrR
uU7RGubaHIidUxTQGhQ6S8SiLpnSALXQj2lEtCc/kBoyCqsAB1POGs3dFqTSMHLic8upPluBaV3E
lbevqQRQDwEiQK5f/4MsBy9m+fZo5UscgVlB4R0ZTH5/eq8ubM6L8VZZIfyFfLo404nWnqYBB5eM
W8fJZG8oDnwWYA6LTCH16/yszcqMuqjxxiIuR9mmxtCDr1nr9ckZDzzneDOrvODRE6nJCX4d0vzv
2eb0GJrTJvMq7sVQgWcOrpE1EOR/bjtc4ZksFGI2+Ni8MlFOh2cnTp+xdwGhrvWUhAb4wipMfnul
6JS6gmuNJmQng9RU/0hdSE+8YhButtG2oez3WpHn5p8b00cnV5NbbsuxSGmxDkNYfWu2W60lyxE9
UDPKVihU8SQjLJM7B6Eb5dQUKfwQ+GOSg4P1yXyrIKD+pzfR5etpfhR+VVA+/1I/IqdxiNFCzNMo
KkRsgxlN2V3Kym+QzF1iN2r05rB8czkmsOIPlCSRS79S1hSic4dNjgBXgW10DLPppMDhwdxQ65W/
9xKY+IPdQcbiCvuSvjlo8FZVcEjcb8cmsYkaXCEBJx5es/7D3mXIVJOifVQ1RBEPTRpeq2U9KnJx
D6b+xAoaEEAFf4h4SFnR8nx8TSFhHg3OT6cloRf6p8onGh+e8J5X0NEGSXSaPZkjqZ/oDzfiZgwt
/3aGzb9AJ5l4mHTGwaHSQl44hnoVybR8AGHXEZVxCqgNfuAw4FTmHfN5ZidTqQxwSrzAGRt62vfh
xusSekPKIlP/owU2zk626D1vZw7ZaPfskxcTqjwcNHmpmfRGgxbRE74bd8L7XUy622qZBdFmGve3
78Ape4Ohpzdlft0CIzRbXvy26oFxcBmgeuUU6iNebOGD8FNmSsLagFTBY98pVZXMjZz8UEd7KkuO
8QGFYee1tQnm7+RbMaDLTJxnpB7C27a4dv3XYMdBEQftPLdj8+yJwnuzAJNABBoHfhOzKSZh20JM
4LXDpoujGfIoS9f49LHVyp02nBjpLf+mhQUTSMSpULvC/4nTdw94HdxJJjmAGCjHUgs9Z/bb6BQi
OYVYJmSLdeVFh1DYRYXRcIHqxzNmIWJ0coLUFL2U6LZ+9+Lo3J09mXmjw90Z5S9yCvAGQsn/ulEp
iL0RXKTIXmY2r+jtpXIepYKTjcw4levRkcjt233h7snQmlgeD8JTKlpGNZ27zLbwrzKRFyWXhN6T
OuJmQVzp+TNsZa6zmgfuRAL5brKpjfD7cOs0YMoNnDaIUAE/ev7sQquT6vGJYHVatDpuLxXzFjbb
jiYYTdZ79Spoy61r9ilGj4IRRM/f3H6pyyCcw8n/n4nY8sgFD1tFXpgGEjxAlHLRHcxSGaqXENdp
VNLyvGoT3NhLZpC4L2QDfsQM8zx/GELOdolUz9hQHeWVKMwp+d9AvTXCQrhZ3twjHA3iDQo821Pc
6G4EtgxUDQKlSCwFyH4xRAILU2wFxS5ew4ndbfW2fkksJcqE2dFkAcdm5PsJBUuf0JlYMnwnr+Fb
X4eIc5KGW9CjPue3LlXsCeWd8nNrk0MCnDMsjQ6mhOb1j0R6ni4MoDq/eg1mXj3Gl/agGoh2xSSY
SrNFguzo2KwT4JfOVoms3pqTqLpmFrmKsnUSESid/36NOGWRxH/3W2fq3sucG7PYXRKE4YpmsqHR
csXYfEfDGBxDbV9bFf0s28QA+3e+I6Zq77K/xmPVrt0hhndBVH3yatrHgAe4PZbkRWmCD8G/ZvS5
sDkkm2dg9FclZhqS+RuWXKl2KQAOBLMwM5h6dJ0Y46AHFfhrXOD8P2iRGYIFpv6XqMedWoS2W51S
YbIMvERBiDMfroL5k2BELhDV5vmXGLBC9Y1hu26pVzAGCMPbgwqUVP7q3S3GICPYwyjP4dTzLmyE
8Yke+d1Dk75SqXRRS9OjjHp0ac2T3yP5WFXmOwJn1UNQXGZ08iN7Xos0AncfR2inFFiFJ90eIDzP
e36fY802ull1F6dq1A3q/y5u2Cfzb1dT94wAGIm5YY6Qw2b2LwRN95JlsABNrCRr56sTh7/k5mFm
yXtE6J3J+M8qHVKKxkOJhl5fwEvtnmbwR9zHNmLpbHv8mYfkxWsp5pwy2Ew06Lm2GOdPwvL/zAK3
bofWs+hZOHvyenUT0hAYDRUZ0XMKCdrdoIaLV26bxordKRkV6KFDhTpQxhGhNZUt2nhNfj3OfPjf
9UiwNOJEHSuzPp6Cb/cObwQ84jxtKq0Dg24XWcjYf55nLFPnyKWp/uiWRQnv/cpBCmsrHzuPkyEo
q3cy/FnKEaq+Gv9HF5zR29yT0h0baz7NNEvufiG/tdMZNDwimj+vTgGTupeZITBlsO1xCyf5CGMX
KRiA037HwpqMaa48BddRJDUu/pRs6f+DSNmDZ0pg0XAktm5/EQIFzPmTujBvchbGqnsbWY5AJm3P
WjSpYFkVAMgq7GAFlqTbw4OkpiCSVOrPSqhOnuV3mjnZ2+aaOOTMQ5yWGCQ/nPrbkTffrKNxMOlx
6TCya0xTeWud8zbxq1l/D4960z24LTCrlICSk0+h78oYJBwU0GM7LXyUyIsjk/RyDLnLWWqcw/Kp
PbNsokGgZ1yyDtelasgbjacCtdCOLDXQ5NaPBCLje1M2Z+vDTG5k3niDyQlLGRJJyw9i7Pkdj+6b
3BXZBBKZ82OzkY1t7BTuGLIZQ+D4sUTKbbk18EeRk6K3BkY5wrPibIbCf+j9lUoJKSoiCUCbKlMm
eXqquk/UsT79EMJBEkY9mmt1vc75kziTw2IGHIiyaTdacfrFSIRfktvRAg9sltya4cL1SaiD/g68
Y3CijW3OlfaurH//4zin1L7gOsYwwsQ7uKf+J4RoFNDcVVwHI2XVM0zvYSehkVqJhgDjR0NIVAzB
uCjCGYtJhKok2B1tXGr3VxwzlR4czsjJXEqok7dlqkAWfDXVjbS5qY3R37Ck+7nSe38aaqJbqi9u
LeaDuR30liMy0X3Z/YHY3aaIqwgXYwsrnscyIrYPjbVOaiGk4kEqf9Kz7cP7u+G7reTYildenqd2
PX+ZAuxnBGpqOUzFZ/YBMoAN1IyyF9kkotWixKBJ2AyQK798mA9Y/Apr0qAokkA5+f6FPhRcsYxA
fmfepfB590EwcH9NrnbUCmSZ8UxF++uF6VDtRFE2bHU9UPLTExPUmWoOSrsSSWmahuVJ5mCaIpWZ
6KKx3FhIOLKzA2fUXYwg5BgTlfBhkWNQGx0JS1ji7Rq7qylTu1d18MWtTGwOc7Ty13Jm3cPLyAhk
nJvj4yby1UI0Sj1QNtL02QVqKlUo+coieOCQKLho4c1bYvDYFyY64ILERtFJnvyL7l/UZd7EwbHX
GNfI3jGEIJL83mOC5K8RI2mN0lJswPopYkNZ3QEhREbhyt/VRfU8h64DArZpwmF+hs+dlbWfnqLC
9tZVgPNBPOklpI77nEMvYNy8rtYwnBuo7U+F71blVVB07RluKYc59REGdWzLnErjt3YPvPHbS50g
s9LoEjZFCdZ+sNtYc1vWfETSKGm509Sm81dymTfbaCZ/znKgVBXRl89TmE0R0kHNhPgq0olq1ya5
UG/Fo9OkLDQQP3akI7+8QZYOilLNs1a/PS0pEWCau/avWWFX6YH60epuPA8j5rDdwUFFBMyJCjeR
jTUl9mRDA8QdEhN0QOwyJfsVGmdv5Lm3njjhNWPlq60WF/IaXPkgRotnOjKRcqZNHyq1kF5IQBE6
MXshh5ilDkOi7mbIZ7E0wlctc3rslnvDtbG2+IaCdhYf047AZZvAz7zjSRUWAdWSZ4XXmBmhTm9G
SDn/vPm6ftDijbm2IMqXVChNsmAAhZbzBYWlRBi1qCTR/omz+Lh6yRvHzz0CjH5c72TWqK59aDpm
uY0a55zL2+AcRMSws46fZjmcMlfoh3gGf4TmmemTeKc5Y1cgG9pZ7m8KTDRpqosrFeForvTuFmiD
lv0GUDcYJLGdre33jZztSUDILloO8HfXuLLsaJCMq+yCUmGBc6Lb26f+vnd/lt4eTfefgfDL+upf
LkOnTRLPih2wwDOI0WShhOvQBLypMALNZJqLJhTVqoTeC/zJSMX04o2E1N+BWI1fkpySWyFutebm
9v6BkL64jU+ywHtwbobMXVMDNQeEmhDTMPzuwrATzVpJqeShR/BAcrYdruWrXRFfiL8EBNZTf/nS
MF/NX5CN09mB4gL/7qcEV9yIktQYuqc4trAqvgJbIcvxmCRAdAyYipW/3WIrY/HYw9BN5Jh88BCu
0cONjsx7phh99H0hZQ1kXwr9Ja7uIwIyiIDzkjqKUZTC6uaslQW8fQYilqCeSHPHbZtLogT7A24p
4eLujgIOjmlkyDc9Y0Z8PKmTDkC881VUD6dFS/GP07Nd3S/2a1affzsNnnfpwwb4g25fdNm30LPt
CWodWNxaBWnbwwUBuk2Y2D/2FZ10DKCZ/820Jur7hgPJ+SnyJucfCG2CYf9fP47hedQWX0c3/hb3
+O/+pv/so5Zx4waefyNEErpsvSUp6dy2TM1KU2ysYZKBNom9++I23C++tV3sRrdX5JO0WzAQpiUl
y7up8W9dAEejDV7Vc1S+0TYyU6NGLwJIOFvHUVOZKcV485PFgrL3l3le2hepBpdjKb1OfvIZaq4V
JIdbNeh+Tuqs1lCyQ1nwzUruf0G6QCltj7wmNeSGxEuu7TQdP//nOiOWNi5uNH5a7nMqHqz9vre5
02KDJBu67NHLO+ek2BRju4HF0gVzA3auXc4054Knl8wbFOubQ6q4lf5etIlxAbVDaRx0Y+HmhjJn
fLmgZtgrQ1EcnrEeyasOfwN0Kb1kb5k4vsQLffeiLcJJo2V0jSpe+Zyxsu/2My/VzoUA72USaAb0
l2xnaxdbKZJ7y+DbSgZp5RVO5WfL3sCSl6Vn5cwIgDtU+X1UuTRTO8LpFuixPkkv4BR2FD1uyCpv
bOfRIoZMUqm6lJZIf60Elqm4/8aMtLZt4K3YSTbzfiP70xInaAu9Rls6Yn3EVCEdMhlp6Hwuelk0
UuGt+44faPK7XZh8FJkj13eu+iR4+KL4Fl/N7ZQlPhYTkfXFr+PyfWn/OXwcXoqno2zrd8M/JnF+
w7WslY2maLwWBx4jRsy0y5ByI+dVC8T4x5yEhFogCijyf8/IrAjN2uuDrbTE3egpzTGphC0B1u10
AtuBUF6qoQWY6u+Mxsf9D31ZDVPLoyFG2G9MABF5YlmH+IEL0RuBe1vn4TeyzBZLF1Hfn1/2iR3X
Y5wxbLH+OVH3xY15zSEiEhnQfuqGH7enRWO41uI8IkkC1OI81qzLSzgNjMYtLZJRO5ulEG21SL9b
alJmEH9vKSK4YwUCoq2iWWFFD+/dendncpmSPF7N5Ovq5tcr9nIYPxFab9JM9Q65xmygDDlj9ZFJ
3VNaPWOZ/6dLxIRheMInuhfUHakDKYSw8+TcmPySuXgzZaz71i7/rCNkcE5Hy2MmAjC45HZbK7CW
YWB3yhFVH4+Ne14Hl7P7dGhCz5kF1OZ0rXZK9lTXp9x3wrKZkoj/HH+Ht1oA3iQbk2R197KigNaT
or+PA16SygCPjRLRL5bB4T4GFyrKijjhqLYKrwXgUZWVNWLVRE7FnXufTDIIecuFrHaofliYQunO
njjVfSp+ugYbB9gOl/Awm7JW4HSaUpud7LNxx8kBm6YXJ/ymonTiQtdVBCvrgrWHsYh1y+7bCPrb
foimKrrDtANHPhb5DVREIkf3D5QWkmxKN/eD72mMbPfPgu41+k+dHPWSJnwldfucIndkoO2eb6LM
exsvRHuzpmXs0PdLEYAN5vWOtqYR2ZpM3KOgTdhy4kg9eLyA2Sm5tG89NeVF9aU8xpLrCoOFiiVu
Lkecnxaqk2ead9wQAnoQ8R+sPl3lVlyv12DySaSbAMUJ6tWAhVN4eMoWJwiD/IYHmwoncSKTRLNK
2GO2Voax47ni9tZpXYR0FkooQjuTI6DpHM+q5nonZdHK9naqMUf3HxHa24Aryb+hdJw1F2A3CMVv
tBzOLvYfgBN0PI0CSHYbK9+jmbi+pJlJuwPMjzommoPHezCBVWso/p/utiw1Lo1I6tUJvJUlrqEh
U3q59pJNh19RjTnOw8/WgOQ4vVIGDERHf4V57tAUzYAlrBP18RtwzNC7aZkPzVVIxWockxqDgq5a
yA4om2RtIWnp1MOLYCpZrPtmHLdaimYH6sy5OWrZoYclfIu05HEiP7zZ6C2vjragCsTpPaShKY6h
2r4m2e4HZvqTOzwB11FVWSlpR88Kx0AfpsZCNDoxxmgvk1tn6cBc1soOWfelslQeOEeLUPpzNxec
+/dRYKebQ7xqUQEnlYStrwCYbFtB9DuL4xidUImmPbFETmDJTIl+/8wZHuVHs/QTEUjHrteS2e4G
0gM3HsNbDS8POsFcWZkT1eZFKLhg17YxQ1UTd/HEAHWL/Jndbp2eYEMJxIxd8LCtgvqy+CeNuNXC
FF0cysLgkk8P3ukzdPDAHp/s/Gfhvkf6L1f7bfImxsh2UW7D+Oru1VEBGlHjQd1IU25E4EkExela
ufCNUWuHyFIANQk64KR8nhzPf521q98L2Y4DZGmOwOiGRtKCYFgJ/1gGPo6F2lAqs4PnQo29uSCt
TbqhmiCINF7JWF1pNesx3Sf3WltWiXPnIk+fb3TD9FRLnDJYFkopbvWbEystgDd820gJheEcP3f1
Jm0FIouQmm65Vx7pEXEIBjN6zwDJRtUib6sj3ANgyngVcwoIKaGztpdydNHH+2DMRkCY9+kaHP/i
O0VIMag/DlmEgTEam3wJ9VQgHqLCy8hIiqO6yEAlFFgxjEhwSPAO2HwKUaGKtemjP1HloWCRgMvP
L665YX/MlKI/wZhctPvcsdavcChdMHz4ax0yebR5iMqYG+SyEsmlgak7QmriKRObygP4b4YizA6J
aSTrKz2b/RDA6zzNBFrGWNb4SNxriRoaEgiGEw7IrTgGZ/zUaFRwdOMIl5WW0yIjcmOFxhGe8nW5
sjM+ucZfrHYErHgYKHscfw2PMgLoj6WttEJ/qZQNO7U+F6z8hgDe9bYxEXP6LZPPZiqeOAeRRmBx
k8DvBh4wVR4Gv0hjwpgW9Z81sg7eytZIkIf+5RP5Zd07aaIYC7paSrbwnKHKdxKNIOzf5nCjTaRc
YdQWb0UG+j3ai/4iSXyOde7ZryHOvv2FBd/J4bUN6gk2WlWPBmoqkeR0hI7s3iWhL3C5r0gLvioO
G3ZNkHSUjGbizgqlTmFXD2+qPIT3I9MzuEI3jCfXi88qdVZLIyLs9qPG2nxOD8PI389WMrMgmNyF
86Sr+CLE54OArzmw1CrNH2cVy3OgiV35YMTrZoQF4+d1XUmhVggN/TOqibR07dlaRwZJdaSKmEl0
89kmC3LlsvAXeEOFm6VwcEJeuI2yDPAQz2wzZcMMS2OgeSXvjod6CI6zMGL7+/GQ97dieNpHqUOH
cqtk8Yr7WIA4psOxAm2S4by7qRajIl3vUC1eO6soXpFBN5g9I7ff37ut5OXSDMrlxrqkCX0vquy9
UUMEsk2LREUIQjKSXDRfSKHTFs3u3SQBULMVdWhpMn2PJGcJtbyFQUCambG4PXL0hgsUvQLj4j5K
jzKNlpxbQjaEzxcNduwcl8vWXV3ldoMLua+sgY3jlaI7dYtpOAsnZBrn/to5f+wG/d4b9uKYgiu3
fQXKKonMT8gBG2QRnSnQKAAZkPagB3bl4Lk9IUsev9Wyv74xqS7heBrRGPs4UzhwJEeFFGqNUsYJ
AKA9ojyHLiVOKtERveFRUUbc9bLxQvcdMusVKLv1L+nnBQXvUq65J+UyPwOScBiNTTXTEx93jQ97
eXaPwsZ2YRXf7Hz0oPtTuO05ea6atFM5XBgHGJgLReVeieOVK4DHzIGXdmTYy+ELODRd6DrjaHE6
2OQHiE7xFme+Is9+mB+SieP6apSpzW4O59Ghv3QL3BRPK0/f2FdS7KZdk63UqcscZTUV5vM4cRNe
ywkbSXFMGVOwM4xTuhMATD51FNs4jipJFXF01Wz9zCJWn9ypBEZ7junRnLUVWwvwyFzMUTnfVXl/
kcn+QFFKFoondytUIYsdshnaxJI1S4khKCv3p68BN/Sp3jmR8JColIo8QRBNJpxElcDEt2OV+P3O
WTFEFodFFJkQDuSjnnBACZ7ruU/8kqxaABrCPYD/H4SR4Sdc9/1YthuaIOEB9Ej4JGc8+meCjnlu
NTxPRR7Djv3kSvJwsPg3SyyHkC2U379Rrf3h/SsirXWtcU8lKAtYK2UbbvVODzNTBHDSEZsGeZB8
9SlF1+bmvLjNzT1s0z7FmlIhOy7i8kvYg24kSUskoePg8gmnesBGy8JeZvH3rbpMBPWD4iUg9ML5
CL/6LdZeYxamOw5flrZkOnEVXLr45Rx7H/q1OcHLwOZAontBZAPBQczzMi5bOb61b2rtfPiFd+ac
AgmIvTIfCR9cI9y3Wi5Igx3JYk9QDWKsN2CXGaJnFFKSd+iwLLE7WH7TivXR/Og/B/bGTIeQltnz
ZjAYnDlFp268jJjcgfqYemMyx1ZP2pYfTzJpcqImXyxeWK8FTQSKbMYHs6g8Pzln130XpO6pwSne
HvXYL1OwfPVBbIwuA0BQ1I+fpbFXG21iuaT7shYSahtDzSY3OrcQAUMSLD6KK9FWFX2F0bukVS20
ajuxYEr99NtWYP+AY58TwWo4Pgrk0d1ZhhcBWJSYje3l42z3nwK5zApozlQWMlL1vyaeFxmIIC1K
Ns8436LJH5Ob+BvPREN2mvhGq2dQcPTjCENO0wkQV0M5CEpmPxk6DyQs3C9qWIKlaLEzxPvtwc4k
UDhUqOwe9zI/QdYsDBhZiC+GAKOfgJQJWalLs7bfCGESCzVbHfwAUOlrcvNLmo5a9wzYQG0six5G
n2txy5OQDzmIg1blcTb82b2uyRrCxm9GMjurxaEFwr+GZzJMW/SWU474CvYu6S+N9TqZXKyGakMj
pbT//v6euESpjpaxVQTaXI52Nu0jXZ1OL+hAYlPpZwKgwqIOLipF1hoiGaSlU/sIg/qgf0TgTKnP
meAL31Ocm+Fjjwn6RC6E/JGa3iQSgUFTKOyG6tcNkUEpnbDST26eI8W75TqVZ6VJ+hp4lZvJBoWq
vrvW81toxLPO+TFfSDWNE7bm2zQjgnFhRh3EohPjTPGpgkkvh5Kg0f70OiJpR2QPjvYA44kF6jow
R34gx1/kOGq6R4z03ALa5ggxkxrBxE4fdY4232et4tPes7c5ct+DusHXNVjQzPrB+DNhKMtCcBmu
b2pLHQjLcpVroa+elDaSknuWXoieRLvWdK4Nm+GIErlCYbeyAxzdhmgA2PtyyDz1BzJAGpxuefbg
FBLcEQH2oaBnGeE3BQsrCgHqVbi0sG3EbDrqgxYR5N+nNaY62CeG9mYXRK4xh5lRU++Y24YX5ZP/
YxqtsXdZdWs1ShTWlB+uY/ly+1fnqcONT4XVNGEIioGM1sB5gLQXb9pdTWAgBlG8uTALd6kfpuuj
3r4LJK3Ib65JFLUBNlhpzRuQmMWN8x30TWVKpcVek09ZB7PyHYM9gtS4KFDlgZAH4OIUEVajqrCW
ZFvc89n8zRzJ+p3OqemwR2HXWT7GdWcpvk/cKaleQ8vR0TZKSGufMXfPORUjdpFORo2yJc9YYNKU
7mFnlWSPUHh+iYwwu/+kaI79/JLJvaI6VPi1WRm5NbKo9SfRCUfQkVJqUbmSV96s2segNAXP2Ohw
4xhpVKCoIB8kJmSoGJcaFRtWtdnTjkWLA3YerGZA8TI37bcDcO1izZWPOhsiXEE92rcHNcKLSCqr
VfM57Iug0x4+ekdFE43xXgmfxvrWts5jxn/YAKO9zuFzeHuCCBGkv1Afxn5T6OWdYAcdN3DUtljx
3+3tyxa/soFTHRzSO2F9mQNwYqHPGgO4NbWSdAaaMCbS1nCKF4//8po926wjBshFLWcc28ks1B4x
sg6foSfUISD4fhN1hjUIS19g0FYkQPY8EvZvu6qwCwWY632yOTgEaQu+yeetai4YI2m5DUQvJYOJ
T8Pt1KXZ5QXtvfgol6722w7mucJFjxJarlnDxp4otpkKb/vK+T8aQajyJoINAa2smymuJf8yZqJI
S3jugHWqYDBZurOoIRCs2YRI4V/1+RFDqlddvTVZBLxJhUlaVWtx1Tp/kzxbg1ienr9W5EMGieB6
AIc/jdjv0NFs9HtlU4OwHs4akzruLvr2poMYfv9lDH2xqCBcvrUgbIw089zczlqRplg3Lyonjnau
eRYAUTrjxD+5PQSayRg6KtHP3knGH6SdQRxltYfK8ZpU3+Ubd2EfqhpVpX9+keGeQhElVoRVJvbI
+yEo2lmi4BhwNfmEcATzeWV/cm18BE66suMWXdRLqFyesmh5ctuKVayQih+tCX4GwX3ZJB+mO4g0
QifSVScXTm4wEJ0TKfBJ4ldoPhO92VyoAfBPDX83XYYJbyjASM6bjloI8pyF20Kw8FOoJzeF4qx+
5VL2AntP20kY5lnN0p/4sm/maEXA0tIVt1S6uPwzZ4LMmXGZttknqmzH47cmm/17s2QAd/eqCG1J
IZ8XJzeIejWrtFMbRrsOVaqZ+LncffOABGKikVz0kC1Nj5FOypOsLwVMcD7uBsDlOBlUmZTYqIv9
4KFcK+S0bkG2EbzNkjYYGgBaL2znDcP86h7EcKyny0K6kwhyo0Xooz3oxRS9S1C98y2y/sr4jYdO
1c9ykmuIYJ1/WUXB8fbVOSjdnyaCzNNacuAMtfIvmpZOl+U4bp6qyfzkPhfJiwmro+4EULYugbeZ
dQp+IwPMlddCuVpg66iLf4e/MNdhoraq6oo4XvyifgOyJ3zlooNY2jzrbWNnnz3i4nPP21mVyaaS
SEI3pCWujHle+gtZrNAEYdQO3oX7VY6DS9zAm/Se1b/bHhMcDQ4AwPJ+QXe55O/ThkNycY45NO30
L77FMUw14ZPWOUqCFuY05XZo2uXrWfiy520UUPqeOCdHfxDyHDSYEDl6OUtiaAaa0JPLoob5iFya
dfDZDh688UWPVeh8VgOv8gppW8bDAEzPbjbe+kLphVPQdolMJIr7QTlWTKYJ2TBiLBiawWQ5rPhT
GM7GMKFrAM5xPPa+rtEHUwWQCqaeGZM7hFIkcS1wPr/D+2fHJ96ycsI/ib13nrPiwnbXepwrA9+r
vqD1D/HlWI08FzpZKR1bo6M4kYrh0GVT5+fi9I2T4lAoqLJXDYEBonG2lSRbGoR2J3jRopvw7myt
ZIirEZGeKk9OxC2YM7B0ggcFr7ZudJdXAMfXQAUHBSrXkQpXT9RTVAuUibua1UEO7wruyY18Lc1B
RcQMu+KBaMlUysc5C3YPGlcTnHdZmEOt9eFwP2pxQfdaAd+9M6KmXIl4/Fc9Yqszlum5MAJfSbIu
JxDmhahD3fdXUt7SnIeq/clZrISrzf4E9MqAHA02/7QuyAyaATVScRnY3zIpNt9wgDuPLJQ2O0FM
ZKfTHBFmsvQj2jUuzZ8papJ9POFNwtBPJ9QZskfPH8N3XuvsCY7Foo1uv1YEjRYlqj+nQhrv5muQ
Ng96hTDhRp/E95w0mNDWJjJZzOkKintWyYdReDgBSzS9BnosDsewsxw742i2Qr2uEa3XKimr+35P
nPrrlriBvMvB21LAX3DXNvlyHtijOFBPoRuW2qFOfObqD6gW0TGmDPqE7n75/Vu7MI8dKES7hwbm
N6U1xkrqMiMbHu6aKUZKUP9tt0t50AxBKcyyT8H0k3soXapnH4QRXjGEWKxhnJVd7Zy0eBDbfsMN
4ewg3XKRs/Sd7RS10gjAiEgTOXivqjX0MfTyI8fE7xn1K0NLWH8DzjNSHfbL+Mhr+kN5GdaD4/LM
DEc2135cudcfa30yZzRqAaM47PKDb2JwB58HRMBE5MG9R5CwSlk51jdonQ28KlySrSrsIkiOkM0l
+eJHENkke5Rf00xPygZ9wuriODSRY5b9RdQTBH6OiyTWMuehQWfiFogIwiWoGYhEqrUzYi2O4xYA
8XezJ2Kqh2amomzxntxW0VhvaORMBZ0Vq4vaTgh3X5WJzuoqnomxdfJJDoowbJ52g+TDtxFo94pe
M6MNoSBIzBFott7C63I52PVVyqt+AjWj0p/+aF2KeCME0KgNvqyszyuP/sLDn80+Z1qSxxGUFim3
+aEonnOHrSJY5hN9ENypPq+EkigMry0X3qyH7TbTvAlPVkkPPnVQikzychZSpqjzc6gE7Nqb1C4O
1Mu3WTZi2nbEi8SKq3f0DAgZw5qzklrYlnYD36Bs92CcFy/FYmizBYO1V/Z8CIZ1n1lXQ1B7SVXt
EgSzh3BxMrzP3WiliuIrpgpQHg7ewjof8UEWW3js9pYH2FADdoGEA62TRV4tOqO3zYrV881yHkrb
Yv3tpNMmSPxfjDDBV2xf+ArECr/k8eLiFKQO18mLaXrm/BVUfnCgqf+VIf1sbUvhDtWFHP2Dq4BK
rNijJtxWOt1GZPzIykkr9vtklmLdMITdiNRq5w/+yM0vqql7uokknDQ4Qzb5jGNhupsOzpru8qXG
1f8Df+if+9O8bjeGjYfdO+DeH3oA0MjSi2zYdbC90dGs7AMLN6jeqHhSQQHSFYy+WA79X4YQP8f8
uA79Kj2a3zY0oid9ln9ZozMLmqtUVlIPIy2HsorKHOxyxXw65DO9J8lKWU3s0UzGMwHS7cqU0Lqd
uZkAdMvfRceSqKMvxd45eRn86W6YS+mevbBWtRg+1GEAcot1mf3h5/Os1pzNgfyEHXqo+VxO4q4Z
qA3ieUcdEl5HFikHHtqcHHEFlhyD01TqeiByFLQjy+e6cHJ38xJmN7bSo3G/Kb21GdXI/Kh5dmX2
M/itoFemAF/lTNu8C/rpH3sE2TKACgK0+/jB6WjLSc/bS9St3fqYK6AafF6+BSl9XPjxQub5Ds+8
fZ1g8xPDOIPcJJrN96JKZV7ntzcQ4pR4C8L2A4iDOE6JMSOPcsNyseogb2Bk+qUTUYw/w9yShVPg
JxSVm8U9PocvR5bHu3uQPmGNo759AjKKMP1C0NE4hnqzl5vxedethPH6bHkHeeRWPCW7pE3XB/k7
HEU5mPfkKjNvJ+/uzNr7uF4plcnm1gzJSl3Y4Fx4+NSHpt9UTtlqxj6V1eJmPPkGiVaitP3gTmLF
JWuby/Hf0L1ryz9eEo692iT/SMBGlyfOSE72jwJIafWXepX51drkpgfnuZ13uWxsxJDrFdb/AaKK
X/uEL7IG2A3MEeCF5/nfYTR0sNm+5Ni+BM7sK+kjOy0qZmv8PqTFwTXInqnUsmYpAhW57+04CxCF
q3FtEXa+mS8J4d1BhW0ubmN7cUG7ljvXyYlYO+2ptoubTiWbO8OKBZWYBjR9czMSeD0PAUAdi5D9
UWCVJWMzp+rwl4daFvSRdAmpbjANPq4xqczWeE/ZZiJDViwQP9HqG30pVwV1L9UNs5jNHad+D5dC
4mckXSrZVBPcEwn4+6bYNtporSedUkv5Nww5AD5uVVGUORKP1tItjMUFJ430BFshcyKjEAi/1QGo
Tw4DKgzwaLDaOS4tRZ28wBKcwkOPK8RViLJw/2d1da+jhgqE3tCf/x5clFsM/1tjTvHemHw84kyh
lxaH00Tm40735y1U/WqDdy52w3heZOp8bo3+5jk33q5ZnZMbqHFM9tlkaAmNfqIyDw7ZqE/plHLD
Fc6vxwkzeJxpqw1EpYB0F80bsLOD3CZ87Y7Aao+O5aGs/9qggpJHOkm9iSASKSo5BuP1olqTXItL
/iBbycsAHnUhUEZfuPBLswsJX2xxr96xGwruWyfKZ8b7nKd6LIT8phQwQSTYMJavG47wy27nMpZV
obAVjptT96EM66g56W9dbJebM/Yi9CDUn1eoF26gAhWMnhPGwIy9Alq++maRbLMK03cfh76hpoSG
jGXh+HZcd042o+L5t0vfO5Xt7feVe9iWl9g8Rn29VQ6KBWGCju8cZ0/MtDYLgGKaXM4F58UgDgZe
We5sZHfQLDmAd1XNhxjnHsCPavVXj1QqSEP6OWqgA6WNupB6q3gIJS/UQqz2DikDFEM8tjhJYEt5
YiXtDuwPLdnpD20M5u6xeelB3lwWuC3HDTMKLaGWt6dupCvHiLrlhUj/9VeoECz7lHc7iiXtV9po
rrV3kY0ZO7RMzxegqXMMTthRhjjego070hQCjlECJw0XgrhvuWwSjfZ6NTrYwUu+XpBRru/YUoMN
3ynN5IWHvxVa+RuFA1bXNqaiJKLN5Rdd8vkOwzf790ru0EPoBEmvitQ1Mi65k7Yz09zn9+yAHmdN
5MLJpnHh80WZyKQkG7O4CdJrBiLJm/qigW3TPWBjLkiNGkin5T6NapoDzgidmW/XgMpk+3KyXUs4
G4K8zYM214PfwMmGS9Eeq0MyZyAlinlGJ89JeskHMHLPQH8cBF8ePpbfgu7zoXDWftmAc86atAZ/
N2emgZYw0DqIAWUJbBa9uQY9Jpl7F+FuOiZH2Ags15Tmhsc1HpmVXl00G9NCHKJKvkwqZDCVE9u9
YqYBAkCrbUCsz4uRdyEloBGl0t1/gxIgsXHNVR24izwAImub5yP59HaWwffo0gE/Dy8pZTzC9Xtp
duLC3SiiLLhTiaCB4B7dDHhfwHla45wQH4mhl8NfPVmmXIreBCdwKSvDKlgLYOTkw1EkcoNHK4lG
3RxFVTOnfKul9I07b0YJ9cOWrW9WYDZwC6X8PONkgqdTPP/akS6gvgneIMxPrPQbB8ZtBtBVDamv
5LkdCfESq5DPC5i9eWoJwaVKnCFdRKlIl2upIf1CYzn0bIIZaeK0HSjBJ2y66oCjLiw2ArSdMil7
jWgT46jnyWXi6cPMQsAnXFIkpb2L46NyCI0wgA+3oFpxJMf8EQO/yqsr5LsM78v1oENPHtwds9L4
tAW9KDUv+OE1DKnhh4kjtJwi08Ni8tF0ypTn2pll2lWFbNqU9rypWFxnek19o5aqCXNbqDNjQxkc
pgzMKLs7eUGsriK2j07kqnzOngAGIZsplNWYl25F2vZoaxJwNTDMdXTT2AhrG92tS+pb2Kdl4rcx
TphfZMzpMGAZzijhQTWjgfUEmplBFl2XBJJpHFY8fHx40uWlipLTl9ti8pSHkUc3APE/dFDZjxg6
vvzx523m57KnGbEMPulFZ+WQCMSLrvZ23i5JZ1iB+W3O6X14W4rWOdjccXLWmrvmv51QfN3zrdUB
p8pYfwf04uHwL4aPCset7qlyzOBxNDVENgKff76UcXQ9ch2CAc4bXyf0ugeup2QEy/wA71JYpc9M
xt7U2Bw8uwnHX/OBWwz499fRxrPC4ZVybCDSapFjr8GzKXumbd1k/HaQkeDaZ/XKwamHvn0wxYlR
VtsE2mKA9cADl7ALNtqLFQgJ2rowW13WYyEC6SFV9t+7IY9cipi5YrWLwWdXXkqGvIrhbXK0THQy
BVZSqL3xrPZVE2tDuKgfP+2fKYuc5U58SqDhdDooOgW0z9X5bg0mtSS3yavzsN520oyW/4LXINL5
+xNqgWvNdQ4oZMoHAcFhBXSUF3KI1bjn791ApTd8gL9shc+5JTaasWGMtzy8YKfNiwdzIqQ5jKqP
/GvuOKcUYgB/NatNtuTpLhYhFRA5IUnVQPpw0d9toI2sPIZo3uUcEsdebEA1gqF5LWX3qluUcNTe
trk2UmJCytCW8s1PEM9BSTCglZi4jdmKQ6EmX/pVnyiP249oBKL7cF36k2lybz69YO49+IxoKuYC
wOfPNYH3HYAI/8t0jtB5gB7C5s9fukWcuV8WQzHX8BGRfmcC6oHTAAm/iVWsOqeCP9TrXkc4B11N
c31cj/8K4vOQwDRzJvzcMcHlQDLlrCMV+nvBIfQGnhFkfkC7H40GUuztC1mAFnKq5rXgqwt3Tmwd
+aqWExXOZUMdWBREw4IpExQ4VIN2vYqw6Lyu6i7fVgITjpXQNQh7RsZ+cIVo7JiIREnbDMDaERlI
5EzUfN8S6AAVZ7AaNKbm+v+E1aQfu27khem1TVhDbiWW9KzGRGeVTvLnR3jFowbYgpC4VfUoSEea
tnIOCQ3K2IiEIw+j1ISpCfW5DSx7s9ruk0EuunsOs6NlQzXN2ynnkV0lpcVpDh3zeWaTVkYZHiXs
SqdkyyrH38KY5Ou4tbHf6HTQNN7kGiiY/YjSMOUbbJQyZoOsU3zCHuVAu7ixPyxecGPQxaEA6dUj
lrr6GBwgUQpTahB+luos/C1JELQMP1PxAtFlg/84arBpw7fIYubdEPWCANlmpB7lUdqo2301WbH6
PHYElnvZ5xG55OSj2ioEtR1/Rxd1pkQO1K2lU6Rv9+oitkR4CZInFI7JBeiYfRcx0NbggAA6a7Pg
ZgrOvU3mExBmQeNVfZniUEVIhNoERlvBuEWwPGwbOVucFhHZRdON8bxt/VPwDJwtr2yhYjrqqmPY
jJ6NCREosHCCKZpb7KVxLtqEIFLynmj0nVd/wVYC2bTNMDKye6wp7wvkclUQnyZ9UGq/Czl3PZkL
3o8KzFlY4dnQwTQK8Em8LevXcf7fNeVt0/ldcri/C2MkYtF/7We4A4GBF0EMBF9d1tVTDLEhoK0V
k2HBEjuQmw8x6BwlM1juw9QNVvlfYL+xphisgpcFbHBuuIjMvlWDW4oQ/02Uao5ZSw0Yt8Jkmyfh
JG+VQ+dWmBEy10n1Y2MMY9fRLlDSDQhdMxc29mS8HwStmyA7wJQx5FHJZlDPsPYyOLgPschDithY
EuIiigCXAV7oM6lYMGPBDH9+NM5bu9RrKKt31QaHGECUF0OWbScW9B5V5KM4SPFe+eeLuRqJBZVQ
YIq5FfhaqfaF7c8nllYupbsFIl3WhTMwb1Ghax6yWPWez8dXvCAl44vQIglgQ/jcuLVtyHCOjWAX
advD7LClqmANpAYZp7xxflpwkUySRUYqvNYkCbH3eInhMqOpN0hwYtWoV0Gfxt3vkVNkInyqvcv0
3BlTOOANjoxJHsD6Jm2CDzRs7tgAXNfNOMtagMRRRRnd4gKk3V6cwmBBG6GqASG8EJ9BgI4I3GdP
CB2B9i/9XKNftW8tbSBIzhjPSncpEPTRX6bCBrukmdKWl7n7O4q4y3iLSb+/Hwt2yXAcwGYT4BPQ
OEw2sMG/zzUvepjxCp6e3LxhKEHLqeWEN+bXslVldX0+iGHvcL+9S2mhu+xObIcHXqe69shjPX7D
u4rDG/Ub4dxmOmT4fCO6yrxXhNcZkeoZgrJt4mAsBInRL8XMpOmx7eecA70nrlMOek7agfqHO7xm
YGbzAyo9/EUpfN31dUYNZvoZTNaM7gTSbJ7xONmGsssn/zNImECU6GQBwzbmFlVTWdwu1Wf7GAdg
K60SXPJVcQuZQWNKljQ2DJb5jvsXSbAXR4Omq5MSmuW33bOd8V7sO2fq1lBKLLfR0wVPVcRSUHOc
9T41IjSA0Um7wtr8So8J9lOyyaiGHo8rx72btWk3tfnR4T0NhXM6Xd3RqkcLiTQDhsEK8c7JqLXv
ahPlxDjPdccGUTJrgT2R7n0M0YuJbQvSCTGl51yfW3H92eFaqtISZy/PAwdSUJtGRF81d/QWpgEz
LF9fJ4TgIeKRoak+/Z7o38oCsC8/HqHfGhrL+O86GrTvE5P9reFa37xM9rfF2wTQIAA6XszsWf/e
1hPPDr8YCTcvSud/mBwZevhrPabKoWZwzf1KctYGbt+38kniWnvf/uyqJMhLjK/Vl4ETtCB8R2RC
VzHIekq+fCxrgI/JdSBXf9dAFeYgpnkh08DJ/XVFEoUf8YosurOAczuNn1vQpQzp9CdDBSYpgAf/
uq0B6uzCgU04bOpktOZ0bqbIfP5oeN9JclEl4tadm4gWnIF29otMy/zgYB9RJQa6uFwODKSdb+cC
oud5HFlMt3Atn5xFRIVlMW9CSCCffbo6bQml0nY79kqbyHD4K+fg4zqa7Burouizn+N1u4jabJwv
kz5m5VvEBGJGeR09YpWXDMIU08miCEvj7eqRrD3uN0UryUzJmUNOvVrppzLN2OdrMgM5kGmdTt3X
Z5l6EmWXmK4ch3vSbKYaYkRBmeI115E5dYtJUAc3BC4El00fnvzLoCwwhEojjCIMmbW65srlrukk
txT9+geznJpvjokzGGGmuua/eO8qzllzg5x807NIxW0QNeho4XPre1etEux2xlHElTPhrtOR3maz
EyglIpn9lQQseAsLLKkILGvsYK+MxtQghw0lIEAbFu+LncoXqOxn3UFa58BaxfyHAx9cC9C2jlR9
FLp0/U4zmT4oLg+GUap6H33h+UleCnRijqhXNWO6F+PgTTZkenrRjqywKozJhzx/TZEnxVXkbHXS
VpS/kQA5uxW+uWAcCgStew9nWkIBIX2GxZ1O4U8lBDznjj4WzDUpirfYG2S4bqlGPcajBjE4lrqz
7HanvrR6pFvRTP+mkYEVgVez1j++we9rQtMCE+fzXsaaW4qhPE7AC3RTQvBgcNriQO3LpLM23hcT
Ujndkc+TMZSoNwAN9P4y6fQJiFS2QY1kcCVQcDHyCHn9VVaRy9eDqJoVA4RthjZFiH6+Vvg2u5n7
eKypxEUndYn6P6jZQzyuwNc1mBYEdL1bAEZvz7FpI5vexy5QhVcZIhcoTvyeAlwGtsrJZW7cm4F3
olk5e2pRb1RV+yxF8btsZFyxabJJfpvv04VbgrB6fxzxbUtUPt5ULwdtXZLyTjqCeciWPUJEg+B9
z8ZQDhmzR6c+sXsCit+NFGXZitKSsF11nb3ztkEm03lV1nZpnuGDk6AMb5ZDz2L5R7rHPOpWrNXW
XZqIwgIeRc7YHRzlhJ9gDQuZUDCEbL9d1R0S0M/9xaNW+XRmFv72s6oC7UjHjgOA8BQmYxY5u/g+
1FKQWKQ4yTQ2CASH6QeIGzTQgkx285FFmT3jDiqJ3BS/XNCenrKZzzP9ve2etfI3XNe/4WV9ZsoM
cjCi+nhXwHybN1johlHLQCLA4ABoL5dKMOFDFrnb4t4QzHlWyXG/DtGRqsKbfNMMW7mi6FgDysM8
lQDw1IcsMsMRWuIKvqlgHZYIuvqun3Vbja3bEZvkSEskI9oyM2Z2nT94esxcVlmYBk0MVR9P4RMR
0oaCqYcLJGgLFO28BWCkpCMbbQdoYtpleRsZOfVVLa388Tn/wdgcbiOVVeGWD96/YhP6wRQy73n/
gQZdvzGHGJ9T5meov/T+fYjDE/wwdwfUEoido4YqZSHOe/0ummoQdhEv8CcTj0rNCwYKgNNZutDc
b+fwXZpAzqZiWRlPMCMcDq7cPxyS0E+U4WvSmCJ5zNo3ztustRxFMBvrttgdDvQQJBZO5pjtkHCN
2sY6uzUnhWwRKjQCnh+L7F8RGwNAynAs6Elmv7C6TGQ9VYhkJW6LFM8zS7CWQq1i60PZMxgGFSpM
1J3pgWWMf8vWPdkERgRTYNLtAjAJXJVqktUdm+V5DweW3UYjaqq6P18nsGW5ocR0w217HT2sxCz2
syYBW3+7SjCGdZUmE/G5hBonj9eRDnICeLk9uCImCfkf9DM5q3pH6m8ePADhbCw6ZCtmZrgvigPn
W1R8alhUHbiNXJo0U4TAy7T+CjtRUctVD/oH8B+yxPVhjypnR/1nkII9uPKbZ84TTm62n8tuLWRM
5xpu5IfLJ8+YXK/uW+YaJJfoEL1GVuYyEidHu07wxYsB1DH5BHN7Wq8XeKwTXuxoQKAKEbYaWzUG
GXKmYL2WclFSuVNneZU7XC9xx9ywPG8zuAvNBDMM4OZXRWME0zZYwDpRr64dRyzed7iF97K/F6Lg
FjPgU2CXzCXp1CCz5IN0liVTE3MuoFf9p4NvJF5QwH1EWBWVJHPOtPUBILlu7IVlQZRew3Ci8y+f
Cv4xGv9R9kzfebb54piUU65CJ79ia7olCGQa6ATmBch2DGwQeVErF1x9LEdFcU4RePXECW41PjFn
7sjrj/GvvjxUG3O5+ugk9kAt8znJLf2CECaN10GVGi+0JSIA3WylfXq7hgOfqZHlAQaqdMzKQ4wH
BW8AgydmbI8iyqEkKd0YeHvjJiLIt3J/ji17V8hYc41zuBgpNIudL78ESc+VHalxDR2soTInIyBE
yosB5LzwfhaKPfmeBAVddHOcIAEjAeuM1wC2jcAilt+p4xJSJQvL5/D60NM3T7/ssmgIzg/0Stte
JCzpi05xbEa2HjlpOdeYirCoAOIPoeTQQUQgqk4c8K8k/Z4a0J/fHASY649vMsdeRsa+gM/sGnd1
+7BBHO1/wKeOZCKq32IkiiIl6uu/REU4NH8rJUX+EK1iFT1Wfw4ppFTQNN5v41L1h2Dl0r86juDq
MuX1DAdUR0GDFkXwZHXOwmPghWZxww9Fk93wP5kIDeEaVwFLRhCga3UUOyDGjNwWGA+ul9/gVRvd
yB+R2eclyMy71zPeLGdmv10ZLhJkw2zNMg6/vPWNeUyD9MeOj17ZQnGDF9yZ+Ng33K0TBloSw4q3
MPcSx6URpNnt2ZWmY1c5zj/yp+4QVMPSSk8Ue9dhbCOsYHqVVuRnvMIqJFKHTaZHKXeiBgRvDgAi
dYfoQAxU45aPwLrrsqMXeIkGpwxdCf03sAEyCVZKPFVirU0lbpmBv4sLc8ky7tc1bi5FHQeqkVgm
XHU2a4BKMW0VJTbATYE2lQnmdfauc5Sdttp7574H6lLDHSNVSQ9oYzj23cbqM52ui8ACOWUITWSj
z1vamDm0gxl3d+5wkSQxOKQ4JUlRXRa4c1mp5zcFwmSBmrbfjnDwT5RkazBCN7mIBX0TnUlv7J5G
6t+g/ZB5x3gQOda/TY4WfxauiTFt+yZFP/WGwD/UFH5S3ydCAFK7kITvfzZUjke28XKJYpmqUKJy
VaAXXCchl9KRz7M29Pcoa0t0MdzOuHXaseMwMxSNognbTjH3wloPAdP08lMuQrJZQMObFPm3TSjU
68mQ6Qv7vt2toDa2L8pJFAKmXX6HUaE8N8bPLps55vU0lZz9ncn4AcFCyH0cRSz2aNOLcaCr5WlY
SSeZdlwNdvfmoP5rIaxxaZ0j7TSfsASe3N9q5ZoxcqKxWlsnXD1xFHt6gCUGTVloKC3XazpiMGaP
25Eg/jHVqoyfoElW06AqdhzlpjSMmTLAo5bcNo2u6yAJBm6+G0oF9GTVYVyryxoR5DlFl5lOnElj
ZEWhVpS/r61SidVx+NoTSdl5uy2qh2SHtzSz6PbxCbHb8Z2W02EHMzk6nOCfae0WrN6ALCeQQD0w
ZpfIdWC810Gx3mtQ11y5s2B9f8tAM5I0Rs1tTU0pOJX83PgMWj51FhqCGZZvtUNW/VcD8LBTBtV+
j8aZa0NbNJN0KXH2uW7QQqOFmATxzWGsJ8FX9pSi5mREE16IlX4dEsWZCqSdI0kekOiRfiepJmTy
2vgof+nBU1A97VMWZ1IQa0ljwdZCbSNq1fEtL1paY6NhJGjCuWUa0dmkeysp9LJqt0aH4gCDxjDB
df1VN7HjOpDUcV8hb94lJLkQEpDH2W74l9yemcUzu5IG+oKESC2Wkr6/EG7w1p4YBdIb8HtXybIK
5+uawNr5Tgo8onw4axdvxv3wem7tbCcG+YfbDAwcjKa1BwC6dDvHEFfRGW1CY5IJVDs3aaXrD0kz
PE9I9b/bYAouGRTU68G06vBTMvmq6z+J9W0Qbq0xYg5ncNBRLTJaygZPqcLcN5+HwSBxxM9OEAwR
pyKCZMGTSTrSoQB13rz09gPRPoSWuGdJw7/zC0d+aOtZyaSXO3J2SxDalS4rdqIRoTa3zWVUT+gH
Oxl4PKnBgGGK6BzVcPoHpnfuk20VH/b2WMM8PBCxp+FeA/azPX5H0F/fQ/E7PcclOdRr1XUeZO0b
bPD7JCsKM5Z8SBTP1dKyV5v0t/51701DvygHaDtPUra14SFFglxhcIgrjmggxbtTIKj9w9CERHKH
BAa+bK2kXn3cuvuwmJwWTIKOysAI5WID7VecDXkONvJYO7EuAVtjH205RnBw427klP72rD+2Ga8M
ktd32YVtujXGkP33DXVNRvj4FEdgR7WtGiJqk5DECvUQlGGU7jIni3K1B2zb2iSp5RGgf/B9sYqy
Jl4ZAlgUPhlV+5w/5mtLcSFSMpNgvOEwEEWr97xGAt9Hu+SPiGGd4vs0YQakRbcGyEmGSrOddM/r
U9aOWSR2Tq5FaenOUFDpUPiBn9Z2tT9KftMWe+vnATKq95d6jQ0fZP/O/5CjSp2fx51mkHuYfcY6
UKtZfw1IWnCahXfpCuYPqDmPmxxhgy3N6oh2PGAt1yrU7DROadBhOe9Lfde1tbrtxDpqDISpE3vZ
/q6gov2s9MAOYIHGDtd20LjwL5tz+Fn3DqXe5u8VuTgAJ6AFGw2Iz4sQwl/gye7rgwmtj86ZugLA
6rJOvJhsBhYMCRhLCCjH8wBtl6WxPgN/u2IMUE7+eK7Kr47XPpLGvcu3LIQmH747+cDwrlqEuy0v
dvlHoGiyueADZaNH+CdYGmKHqAr6a2auCYjQFaBEgyWuznvQ7/rOQ2OGaJzRw7iHp0h7PgoEQfHE
LvSI2TxSlr6oPYkeK/Xc+FO1oEZFx1Jn+onE9hVwocmXF/sacWPunIRT8HowBumUr5CATfTmiDln
QiY3KGDjgwDly0J5IgrMHE7b5OqfnksLbCwK5U2mVAZUlX84a1/d2XhYDMcXh3PAtchQPM80Rp/8
76TygL9JAV56BJ8RCmIX6YJSoHbrMey7hJv6P+5CXW889zE0KwzDRcQNI8eBZNG1j+ZspdK02SDM
I2JYQAZjsAHFyMucCUIDiZWgxD8g87Je3nO4l8vgMnyuGI36QzWTv5S7whrY8SE/CBuuirYEA/II
N31Khsc/Ib6WiuQGs2ByDmU4qhPF7tB5gAGek6JN6jRb8PNmtNTc3GWgdwC+vth4ttw36y/pYHcw
5rv/ZEWf4cFJCOMNfRN3Zy/iRx8r58qh7izWnouj/iTaUNxRShyqFrzAhoJPsu4VTdTDA6QlSCHf
eazq1HFxgT5YuEpTUY1eJ3H/WR029XWGqn5LSzbrgixmW/b6r2NYxzUTA9jA9KVeEFofmzm2diTV
bkqhOWEXsSNnDiB5NbRpP2OwqeNhRaCXDVxCQ6FLpFa5SA0oCgm/R/TyvTUCNQUt7jh4tQalm88S
xYQpoGvWv/1PnmZMqasNwgn7tLpatWz7NTwfXiu2iH7mHIt8gy/5HIl6aEFKWsWyB7Q0elYWbssY
55N1QjENIEcocJ1NfCULWDWILk17cc9nVjZ8O5JgQbATiBCgsYIFgz+vtzTya/w6w0VehL5fUC5k
rscsrayApAUAtYe0a7jJ6o6PvdjRLOgw/ca6jjROfEIUAf9V+KNQYkyAn/Ng/67ilJASukQvIphM
7HDHyGZOrEKjIwn8TFJiVZe6BxB6y3Pbq2epkjJgObLnOcztKmKpaD/NKERKpgWPRs1B1lIRAV0B
bO6V+SXorWB5KdKH1cUlW3rLtlFKDyOgb1yYG+oY4p+HHI/lK0Ca12OORaJPgiwi146rIwmDfwD7
mZJbNjrPce7q24dGPhUpcHr34m7cgqgIkNkQmI8j7pki3jhnnTgoL4asPiGx7g48IFEyAjbiTNlU
rRshMiXvu+3bF0QYvpcWj0gpouS5EhQzl3hiByvstkv1FQnRKr4knPPcaSwIZq+SJGP0kAWa+1md
+8Tb9t7VPBPoUtwjmR6j5/DH7PlZVUydREL9v9ByiKY01NSC6wp2cx8TUI//Uq3t3eseE+d1MSp6
baa9q7qCrE1bJIMR03Vo4mL/StJSMYb0gY7qXPkG4DlsJjObEXvHNdrhOiGNbEJuP8f6c27GnK3b
3fq8p1HxjbgbwkYF7bROmAziRx0pEG/4Lb81dZvXo+njFQogtZZVFSjnH2LEl98vM5bSGUN88+/2
YrUpCOftEFhkMnociTcdJuXpO6yXk1UA+QeH7sXxvyEa0qf0K/uEALAaaq6SMrKW8OH3We7Pkhhp
fEYa5FSW4afgRmsLr8V4KkpVTYnCxCRgx/WltkvJR50aLqBw197QSEH2T0MQkXzlPbkeKf4CkzUQ
t0AyMa198NsRo+8jokSzJ1raJYQaC03BdObo7Ea+eSojuYyWQmEZCdvA+zlVUZsr+E6QS3rvvtZN
fg96F/T/arJTjN/z985+EG14mR88sGKxhb1hCvC132JnTHSIMjah5/V2I3oMsBB7KgRYzQSMJ3CI
NiPClMcQqP2glVvZYUkm/HWn78moenJvX96o5fndKTXut61b848YK6u2BwmpD6p8gCTXHlrQnWUF
cHixyUxwOcEHgPxl1L7uMODKZYlzXsF31IOYR4O1Um3bwNsrUUxsJyO4aZw8PUmpm7U82YRyCHBi
bJUo+q/WWg5YyGaI3hLmWHmh51ENNWB+m/ah8MMWgY2HE4wJsdZ/P7CSe1ILbZ7kbjIEHENW1GFg
M2s88z1tL71zQI/pEBcJTNC6dVsvelSUjc/WBy+vVi8Yg7PEVUIB81d8Ra8Tv8OPXteSDnCtgZkK
H94lXFSW7Jvzgrs+yLS1NdLnOFMBymTuvJLpnt6kKTcGwCvrpDXrfqXltqZ6mBSQ1+PVKZ2jv4oK
egE7sregCRvFeSjFSNUzNrGVfKOXD3mtetorpEmnp89qAqBsbYqy4UBpYEdllx2NiX9fvmRf4d+D
ZPw+THZDLrZjOMJcS6oIFkiBmg29XufwBb2Tjzu8AvgzClYt/O3ic89kNV0GCWVlb7bl1v8jkQmd
UII9xmjEpOW4QpnK8Cuflp/jHogcsgo0DbxzQn2p6UgLk+E9B2ZTAg4lizJJTbczIlmK9ek/d/Dv
MF6JWjEm+H66GTsD6HHhbGda44DL5I9jophls1upNAIgDs0n6SbfcLOMUX5Ke2pAm3I+KRV0Pud4
Ymt9KDxKpB8koVZO9cx1MxUIyfvLJLH9RsvcC6kVsvpXiwm/CzDD5Jx8dwcMKl5ggVxiWRaGxBZ6
m5AdRpm9EP5dyTmLztQGvAbtoTb8W57uvtGN957D8opkma2E/oiIYu76AdTLkkSp3UNJ+CJEfNu5
HQBwndw+Cys/jZn8pGeM8vWwn3UejiJGK/jSSIIscjA/u4svdzGDZybXqy38cpd5vCRtYRPlypJq
tMw3xD0u5ZcKDnPOkSAZFFTM44VHo8Tybpt7eroFdlmLSQBurtl8PQw4XUgSCsevWFr5ttfL6agH
1Agnsq3iuK8TvFYhBiOMmLR83Pkudm1vEbBnBTzuM7ZxHQXSeXfWQEcsZCr+VB/hi/+NcOsGI8nR
FceFbbJVH292JEaHEKvD6/o5Eli+Z1cG/avfBnWezSFrdQllNoUz+kioCh4FxCIfM/7eEz2aMhb5
Qo9r/cCOau2HfVZgDscAHx6NLoS/tEfzZuzlpJeTwxcx1gtx+tiXd0oGuvQVBMFN8vk3S2taaAPZ
yc4oMxu8xQiVU9NHcjre1qY6qh+eBFhSxNd/zZOEwKq55VjsElf2vBztW5KBGcvLVSXSl3VUnM1A
Hut0u0cJdXCWFWjjNHhUh5T5knHyHHeoRi5x38KL5AXlNAkYEvqbyUl6LbI3NLPBezaxDL4Q1EUm
lUTRbPxranigEWgbbcJPFqyruhY/VSlFhQ6KHxcU4DrQLMukXHEctL5dvQUSUlAmLN/rkTv04nNW
qjpDvFS7LzPW86BIYSbwaQ2BUHZIsYNpoZcoGVs0zWLy1ATYRd2Q0bFeWeuEFoVu9/+ZHl1A09Oq
HY1GQFzrf62RYTqRyF+GD9pSPdfNuvO8Ycm2wxqwnfAwRFGjhX7ahcPbpH7aZ7wlvGpyerK+EOqD
AITZkrGjhu/77VndKezLexG3m9IGArB7w+dQBlMhwad9aVoQ4ne78b0HKM+9lidYDvYFMEOLCKhA
oiN3rU1Hb4EvIqV8MOs3q1G/LY+/vS9q/SK90mDELGrRnKmJhYOKYwALjPcB1QsfHyJfxnckzsVO
EFfE+AG2A8E8FYGGr8ill4hF2MTzMPMzIkAD5vO3XsaFTFQaecnVeiNG4xJnt+5FTxbPL7NGLfB4
VMinPvZC+FGXE3Rx8ly2/OLnA0YFOS0AkbBEAJBTDHOZ2Ribt/BOm78BxOQzwB3MiZNorqoco49b
FwWyPhssvc+Sfr9z7fVAYgYqctI8GrrzZdHb2smstKNPZjTAwz3VtH/Pkndo0Wrl4KCThCPYmBvJ
gla0Bo4T1kQGPTNeCyZpSx6yv+HsFRViAhvAG/C970XhdCJ6yNU3AzhFaZi2REFe41AoWddVoP7S
QxfYoTbd0TZfvmHqojJqIRKqAgnIvX9CoQ1jAEh9UQRRjB81N8fgne+Zf9XfupUJmkUZkLuL1Kiz
jMeK/AA+WTlYQQpRJA3oaEGHsmPmmN8xn2kraSXIUdjkgeKkGiSATHfAVLNskYgj3VT41OwZ6BsB
rdlgZ6qmTu5y+HEowBh4jjtA+RuRNFT7O/LBiRxehs7TOj2Xu6Itu/YUYrTkRvelpLU3fkt3pnvY
Xx9qzwxm092mlvtCPq9Egx3RbN3U6zqYn5iKU60/C0eC5i/lt38Yc4FWOfmuOJksyALng6sErZiS
cBHSZseVr4Yn1xQFXAV2a/uXMSA327nayjr6F5xJxNMSTxw1fznYdN/s3T4tZrn+wBFwM0fIFjUf
kBxg5lGrFxcozs3130OkL0RkuNRu9NBxmlwDBXvqscD4+2NYANpUhc/ILzx0YiJtSED4bL9EGYK8
eDL8xgHJyTPeSnTDs5ThrBo92VP+8bQtjRzawTnA1sdgWRXNlXhuxphiA5oR4wTbK27dzgo+gCSz
gAx1Decp0I0e8sDDdZ8+MJNit34fRR3roXRQtSRyhZFffpfSqx/KDzupT/CGVn7ymsUpgIch2Oqe
DxvC7MPkJ3ds9Ieyv9JIosPWLgcd4rIBWEUwfoAhDx0Jfq/J8EPw/ecfa/nIPH/z4FAGB9pKPpc4
bqw7cT6vIC6FDZR3TEOzVV+y7whkRX9qT50Zk7ohYHi8oUoke2zoIGzZSV5LmyRs2kZAkQLptT6O
W/0SNLFyZH50ylyve/8E62n5+TY6xnt0b2iO3Svy8fa+3euJvoSqziNYHxfYXi3fvLTiSAlNTk3n
wRB4IltwkXT15DFRrfHc/PHZAQi2v81YhubiCofSwCgFugq4ZhasrMZ+ZnStBJBeKdiMlWCzaauR
V5xaf4QsQql/3XthnN1E76cTyvYeH0G8w8PO8JLqoU9KpKSnBl5+H6DUm7uQuCGOAwtvw/SRbiBP
f03zlK1urU6t1tD513CtK7j2qr8wNMMIzcf/EFXGi8o2rUruqQtergb+YegVv321u9Zmhha0Bpg4
7W2ohJLEOC5E4LP/uOVSPHr4zp8IrnOieVyOEcCStF04jrjQtRfUfwthu+knUYwx4Nv+pGIVH6bb
7WQDojSb5A4a5qg/o7uMMccDcJ395qWrZgHPmTlLcn/INW8znc1PD8acDsh4GuOCsThgfohG2qag
OJ5z44aRLW3qna6UqfgCoTPWgSQ7BY9ExZmFLYo3f3pHsELe/+/I9mX8xfNPaFegDO6EtpWDPzX2
shAaPbSsbrJDRuIbFTAXHt8abY5RbbQnsONvPRlASxtkpfetut5obn/hVkU+c6YRB1IXdklxXx51
XNDi2PY3cqLrJ87akA95I2SH5kQ+torUfsCq8AlTx8+iNHJHRRcvFbHFsw5EZvN7ZZx+pRHwnrny
0Ecl3R5rD1DYME4gBwwAVb1YYv8NgEoDL4s2UZIUfxefCasuqu9HhjbsH8IHZYlrZiP11SXuvKKL
IdDduCPlW24ioUb2tQWd4MrMzqZ6fiVjGS4yIMuwP3pl19mYLRliGnwN6WseQVOFgA82z6HBzVPt
+wO4LIvsj06M555wgdf5e3+3y2czHA9P9rZuqkiNPdhy0KuC1zrk96rHxS6DQvfHoRBbA6u4B2S7
KId6fE0xsxo8RnRvk1PS1a4ywbLDHxjfWIcA+Q8USl99NL/dYDa0J9jw/C+Q1zDwlJZWUA0bqTZl
YB6Kl/3TpipeTaNkeHV3fnwSiJHtXYlZ+t5QIMj+21KUwoqnQib1MMWvIsZieoT7rgqj8sKEsqLQ
NF2ME7JYJIzrV6g5y+m9C3i/T9CkWPdxN8O18jZCF82pVSwqjRwzzOO0Xeo5WxESaCw/lEnHFLuQ
JEtBjxhHbiG+ukoDo8Q4WptpRQKOdx+pvnHB/IcqzFbATRqEsO0uLhVMPi7Lt4wspjOCmElquIgn
tj+Vxg/Tcn+De3KgecYRM6EW7qh7GB+GNUM06fQiQjfC+t9nm0qrpBt/XKT0pn/M26EGc7xTDqO5
lpzjctHwdyuGrKY7bveZUOOEjcwvrZFYyzT3nrA62fsjJDewrPgzO/GOSukeTR8DKTn+ziGal4jV
DuX+ZwggA5cSs5u698zk9OsPuU6Y0VOD/RNZJhf6T6ND4RlzVhVEmsJ9sMnSSTpeoG6E2jr8FId1
WX/sPF0qhTwVltA3F41LDeRt5VCrdiuMX4Hrzl+3HCtpHvWi9zMsgn+lJ1Y2q0MO0HLrO7kXB9xK
5SOVoB1SAteJadaS0wRMG7ZX7vxTB8ekwz9yH6nid7nu6tE8ta9XKXK4PzKABZwoXb9FbaFz2qZ3
kNH9tgd/18MPba8zNLmijNZCo8me8Yel/4LQWMkbsUt4arfTDbO7IQqLkZNUxWs8vBb/Ct1a5JzD
zpxb5KpFyOrUZ7aXsMEs+dcFsPniEEufNUwHDH1k8Q1Vt06HOyb3WdK7uYXtQpM/cbhrb/U4QxzR
blUeHB9VaO8OMw34JfLVyLTgV2Nxfl08W/mRi9/Q+UXC0kW1LzV6Y3xw8VtxVZpaVitbz+P7Cbic
ufc9BVnQgsZvK+velazOJGZ5vY6lrKeISWLgKtmDd97VcXt+URjpVyKE36oungJnuRJpwoL/mybL
LelanUxNFt2ZrD2b+dtWhpufcPazDpv+ZKpegZ5tO/cDf836mPeI/sIJt/ID7I1DXLSY+m1SLLQa
Y8q9ej0Xwn/3Tyv1OqmH2UXis3ZS187+t460cxvlwpnkbvlQbgxi7SwefHbdWXbnC3TyQIvsS7Xf
63JE5ZedZtal1MQFS5F4rJTrXHo3Ky/BUtJXi/3I8l64A8fqToyBCcU9lg0sbpJIeuCrIjBXCDds
4dHgFIJw93UsOW727XVA/+iDbGtDvP7hOjDRSpM/VtrEASxJqhMUxxZj5uydPl7c7tK5YZvvxR8m
YPzifbwjHpApqkZPKtcvEaJUlVBaY7Ze22zLHuc1C0yAgKdInofOqyNTRsvUR6hRccoDlFZeh3uh
QEJjAjQ52HsYwESfwYA2p08cjvBD3HDHIyt/O5AkeR/DthuXmB5IDIYi6mV46w1iiHXBl58ljcPh
zQzAKjLLVPZKn6kPlxEFLIg5TEvITRjj+9zekpai1M/QaZY1kKaVWJIRuvx1Ktqcr+ae3l9APdai
QEKYZaAHoav6BfmN9JElEJjDRyqGziwDNafweiDvZLKD+Xr3mrPrnxMUgMnP/V86urO8tUfx1Ik8
FMZ9tfS6o0KLL/WJwhnIKdjWd3TUoAtMraVu4QsWZ0l147V6PBh88xOOXN6c/ckuj9nrpO46kuRS
LpfbHZbwJAD0Qw14/A0MBzdZ8o9mxjKe/MdITzNY9mEYx0WJ++FxirINrBpSEGJqZx4BcBDpIZQo
vjCPcOAm83ZtKhvjUj5mdobUtdZNAoqRppu3bm6Ny/NQDC2FMMhz4y9LFGZdi2+JHdgRINT0gR6P
i00TrsyjZzAp4OQ+Q7vSA2rYv+pzRDnVgsRKDrzdrFnGhYKJvsqDWbq+4dKR5gJdh09q5VZfCHNk
vy0h6oJqKK1qCYPRWETpZ2DydNXiQvu8z3uVob8Mo4FY54ohfWuzh0Irdz9QVrQR8Ncv54nMFZ7N
6o8Hu//txskVHN5Pwm50nxhChxHxzeruCBOG4Qp0UUIKMdZg5bBbERV6LrSp8/eH34Jd4Q7xjfHd
W8c7VitJ+0jvfVb2NKiJkpWv2jXeQkKywiHi6WiZGWfcBLecHjQjsrCuU+ZftZGnMxtXce4pGDZr
T9TU1mGBJWKWWsizBscwLuVvZ3Kld3hjrQYOrVHAbDBEPOfFlblq0PIB73U9xzn5gBLieXEBAldH
81pZJCTv9uhHpsi2NipAleFrO0+BmgawolCQS/bnmQRZTgo66EAnjwUsqXlfGChcfNEcLC5hmmIX
Lm/iAGoXyUcMKkrYFjdptqj3+0uRxJyqQgkRGzNSyib1688+7wkruR1Pzk5pPMy+vCclA5yyxaW7
hKJZAvFY4f9z9mSVGomasNJOzqE8mZwJxJl72jAK6Nwlx95KO/z5tQWq4+7c9rILgYO4N2HqWkyc
LL9qmEiPmTxf0StNHFdFHU9GjXhPxmQ4mHyhT5Euill3yEP4AZUWm1okcfzOzGPWiu8XINwuf2Bt
4ur0QsenE7eRzClrzlWrHXwSVmYEQ2DdNO44VD0q8JP9plnXRAqtabbSb1BxFc+nWIpH2gkW/Z0x
f3EWW4zzl24hvQBhRTtZi6l17Ztn932l3ddPdLMptFRRgH593LTwlGLT+r0hZAk1g+zrXpqra6SB
vKEGIpZI9SDiczNY84vArbvv5EYHoMLMJCm59KVZJO/Mn0mynlkCDiv6fEJFQDQMQuRnRF2x8YhC
iuJX73hdclyY1R3NveqQYMgnJH1L7yrM2YNAjIJOQ8EImnu94UgYgkRJwsTavKVjbedWg5g1cYqN
Km7FgSEqCFxHxnY7y8Paj+1K++qNgyQlAowKJKScxsl8omuMjRPGRLE85hQygBBBpQhHCU5iV7Ur
lxY9wQJY5ugYIfpECtvCVLu489YwPpYExy5TwdtytoWYlsWaHSoxUK3D6SVuPebhjX17d/L/z2er
iUrcVi5PT0LPxa8E4kR0wX7ObMylG6c+NAeJGUMYy0ZV1VlbPSAIh4SlLh7GhmEE8PQ2kefIuzlc
osA4/DURwyefD4i2bKFYHvG8cQzqLzqiHRDhFROhLxgjofficBbYYVJfttRJYlSpYu/1jbm0fa0k
AMJT8O55JaZyJYJdRF4drwIeSQ3suctC8KmDi2M2do4gAUKpIsS7N/q7ijkPDRv+gz4W44cP6tXr
1aa5FtKaLrkPiGClO54ey01piNQ23sII+VbwXJrIlijTIG2L0wxcMfEeAV6NEvT05vw50sCfa9tn
0GXtMs3eYkoBJNZSIhZHBt7p+5q0pSq9W9026nQpSf0GZXSjvly6hNYcPvLY3063i+sCCGqUrV/7
mZDEWYJnFfHFkOnINl7r//4C4Sg4Z8ZCsehXyuCWgqudJhzHJoL5qWdqKmq3tgz0GBdhE/KxyHto
Li+xVUEVqUuBa8rSi6PchRRV0te8T+FA7U7yWkFNLKVUpZ3YvwGmhMUsaYcd8m7MbfctE7+OHUAr
NL9xRrykUmQQqP+TbYRZZNL4liyDK3qH4mYuCK2HYF6nDvLX+hyYt18fMeXQoeE51NWV7+C2BlW/
iDTazeoiJ3DTNJH+lkjtg4SSFTsMMV2u9UHwR+5+rydZne2xVrGpiFSSnJg8Kf4LmUvupmcVw1l/
U4zjut0HLkG3MkECdoHPLbni1j73gD7IXl1jMwGTreMnE6VwucFdahH6iNEhWVrSsFVWcyQdBuX+
tr7thK06hcXY+RKsi480gGFciDRG5bCsxVoblMGEb+dSBL4f+hesUqg+fo6FdXnm+YgcG9JHL0h6
S5jc0H/Cfp/rUoxWZqP2Bpvy6s1HmN0mUIAn8Sd8BwEXST9gGu2CCqErhSOQQCm2JgCLEUvy89GT
fb88ZRJ82mrh9x1hcChvk8ONfGRsraYzDcMqzyl2ql7HdLSaRsuQH2ytB4Se8LYaupk/Vjo3UvNY
1yFKY/KdkEfy+Y0Aiv6JfKjBn4YMqpwHFd1egsMEXfT0ylQ8+OmNI5dY0cuTCYkEBUFkGFCX4TKn
vg0SEW9ihaWIa8TzWj9Rg+Iz3jtQxXTdRcoqtzE244RMp9+QU724aaZSs1QZ949C3bGVqnS+Cqln
0+4fYeRovrucyfBhScKJ5pr9N1NqRfhMVbDI1y0vnzV286oSjDmO0nxoGorxQFB+PoYTq0QX//oB
ej0ZSHzIr0Z+N6FUQf46y1wK2drFZTkqCEUIWecZPbwswCTqT89sw1Hd5B7w+LoBiTISMy6v0VAe
Maf+ouHEyGGf5t3Bvqjp/kzYT4Qp/z0XDIGihz1vyhLONS61dRu6GYibs/X0EfG58gXEacECzpCb
BJHAFuqQ8h/TI+wIlQ61A7IpbU40vEiTEbVvcWGkpxhTdE+r1OPRm8q8Bi01zF4vfNSGhAMwwrjQ
UCimPaXJgAVtIHh9FMEkdHm2QutfVhgrSgvhvUFITQHtE3RSoO8LMsxlAR/+Y/VjuEdStwpOUxwL
y4a1tVPwBcdukwCBaQq8gXX3IxBO0lptnOHE+E6z5YU+s17HTnzOkQ7ZBBWI2Wzf/iX6KBt5YPLy
4A96zqQLjYCTsG7+8ltDsLhR0fB5n92P+tl2A91xgNxc+pMski9BGtJNapBzZ5Pe03zySyoRH06K
Le/b0N/W2dCbjty6i3KOCtYscywVMFAfLYZeHVUeELoNo5bEVFqfbskUMdVPLIUzqPMrrMh0ewN2
sYpoxRMe4OQbFshGx7EZuEnxCPI0lmTelL2jO7SNhwmNsGj3beNXcvbXSl/eOwWf9gUfUri+nFfd
dKuRaWjicVXan5LuNrb3GfSEfx1Nuk7e5sjDr86ij4z3s/fUK1KLAYyG89jCuR9zECaNuKcGs8+R
u4HgztAoY1+CpF2S1N038BUIk0kNLJ20kLy/9dCwl2j+G8Z4/V7ggt4K0NOWv2bzZOhcdxUntat1
MxS++Kduw1jRPmRXGsoClzyhBzZv48EjjnpgfoNC7o630nt2NmhBeptB3GpZMCPRu1OYkwX+BB8s
Xs1sbFJPDIhfQPdaqNbAVQfcploY9gfmWU28hI3uRkkMU5ioP/8L/onRNkm20JNh0ttg5tTVO77x
8LqGVN/X59rxTX1YfXqAC5BO0T1HX/teCKjQghlrskEBe8fyNmziRP20dO/PZzv7GkrfLznQXIo1
Oqtnb6rAM+o+l5/J0ASIQv3QznhGjecQf5vF/ECGpAPDpA70+QkUy69yeiSduT0az1XgEFgOWwPo
BYEr1NHx7LFuMiIDetUCns3Z5ESC7NM700eVULQCvHJT5bpB2vs1c8CI74MHXC/20f6bhtdloyHt
FvTSy7dRc7EWGyPu9mcMKuGlUYt07mRTLMyisNplXAY6f2KpyDDa9LnGUQ6jRxC6azuOghmXA0aA
1zU7NVJSzjwktzUIfKocnC/gH6kuuLMTbmWKlVlzqPfoWeEJiALdVOulKj7pEXVYO8ZdRJB7j3uj
xk26jnlX4YdLZEf9KEkMER43DySJ2SCXmD3iKpmI1BAJNIH5FgmRrnvmXOf/LfcGeAr8Wr4sP8mc
KOaiScbgXdNdJnz4GR5wttsjvTGQ7JRjcnGVyMw8Bu/QSyTI9bAGtYwndkdwTbkvWXtt1PRsCzOq
Gg1orp9nR8WCUn5n4CrkwycwWMn8mYtwV6KVaKSIMblq9mRDYBD1QnN/qhAmmtfESwGtMiDkE9LB
B5a+Auf0aSd/BTWGyyd+LylQ1kHaInJn24kAkEUzX3ypcXW+AqrUtiMZMG0XwxRjSz9r61abA2dm
uktAOUKz9244MTq8wennCkJTE1xrdaxNe0kfshpkDS01TEkQL/Ed8F0kV1tQ7O0KktvwPvBI2/y1
uXYbNg4bILqG9X511KAHq05yUKZ8j8dduXlwRzcsXYGT5w98UG1l0Ezu/WABx4/73vQU3gSd4HoZ
GcmrUEibJNc4daCZnestkOWK7hLrlN8dio9IZwU61hGRGd+zwWBc83q4BqhrUFtSQTTHZNqhufX7
rD2DFCbczSgO5B86RZIrtYpOBKtiIe+6O9AuwvD/Sn690a1G5XKLcGmpH9QCmIF+KkudtalJi/9A
Ktc8xSxBBAeXAaiL4Vt/ezIwdHfI9CstTsUtd2cB/clrfmPriSRctd7u1G6z/e033A2KLHysY6o9
iXzxb4bKd1kO0ZMcdaiMvCpKFozhZIllk6fnZf6HFksB0yVrdh/cbrI2k8Y9BuyqnZqsHu639VOk
WwA6yAPNvnHXwvXJoVgrvKeksttz64Eso4V/++s2IjjaLU7hgBnjEL2tLguHTZSTVV5Mf1HFGgOJ
bieF9ospgn7pgeg3Q+SgbKjPZiOcRfY4UpX6KYKkIk8kyX8tTVvaNCcg262pOmBXQg3bO5VkzBUn
A89Ko8B3B5xzmuOpR3Q7OTs0a0U+t9czrJnUmUW0PxCViWges1h0NnXCGw7zDfRrVALWIumx7EPL
eOfYyeeb8fiGsvkjcOalu9oUukwOWJePWAKGb8qTV4YkKDA+yJ+ZfFZi2CrB7VNqZmPA3JVHgPI0
xMq8DnLBh2YCiQ9urCsz0roAr7xsORP1S6rlTBNg09xrnXAW6qKZBE9WgIV13fjTGx1ry3v5v39z
KkJNiU33oklzC6u6UNGv1GLOSZ4HfHSbM7bSyVUpMgVVCCzKqC3M1IwzNctwvpxl294ViTo7AgF3
a0RMvXfHRDBV2MokryitRljVWbvAKf7LxuyTXSXcKYIkwEayMn1zQeW46/tOTG5wFITqr4KTw7PX
Hox4v/gKNhisjgE1dCW6tEKZzyDQZK72fD5zrLr/QPpyUmwaY5CaehSW2ARjAFK2F/E56lqOGg0F
iuhLpKdhdmcjyFPmOuRTW7ZFvLYl9zlJ5nAnlmB2Rs24FVzmLVfiPddjSxrh61bcEcRpQcO8vvoT
HCn4ywyCkP/4+xWyZMsF2Zh75nTIyoaaVsiwRKRSlPGrolBPjcbWg5kV2/LPDlL3rVNjpSgwo1ZS
6/TqHV9fbRV/8OX1k+IBTICDkvm4kMAVMIxWXRLDCjAkYoZ++SQDdXJXOVYnXjr/XQQ+n9YwKEsV
i5/p7RbaTgsGtNQlfKdrJPv9UeBRBv+2uqzqsEhK8NrfA8voqLDdlubzo/p/cFlWE+78vb2LYqef
9aZe/lSgBrRA0tlJB7iur90IoR6UVjJAV/hUYKSv6vtugMvQipBXTYiemn0h63zAfGV7DWJFwbmE
Czy4I8eTb4ed/ceYZCPKUWgM3l6yV5vlXR9bICGjpsYjUVMc6REMWOLmbNUaGp86k32l7LDvfz1C
Zl+nRfyZVAawpVv7wLu9s+De1d/8RrNKaBca6Em+V5LvteANZqjEsF56Z4/uUMKxDkYwqHsO53o2
G5KPc0WdySweU5LhrI7QPADWp3XF5wwWDF0XiBygIhPrq8YkR/UFwS6JY+CPBlBhvMHONxII2NdN
CYzaWuvB9LJXZ0m2hQIKSruF3WrohLRhIzSezq2xpsFxDhQHszFY9OQPIBipKI1PnnhN9h/+C+ld
suZiiIzl6Z/kkiSe56wq3loSy1T01zFLqVn13bZammMPRTC67AXq8LFp6JnnKznZpvu08ykCYZSP
W1h/9tSJk+4KGFnAbnZHoRtR7N9DvTMckFfDyHcwktC1ARc8BAkbZ0rjEScAVfUg5GNS+hVW8wFW
houFIJzWuXM3qQWum2ml8BO0RO+kwgNBONKN2X97YBE/bVld+EMtoC9IuZgHoTzl+ApqizqYwi79
bNWYuJ3CCgQF5JIEeP9FbEUexD2R+c1mCvi3JVrGP1G7R3p+D0ihY8kv35bVNCIqdAGNrC/udkc6
yMgxHmMx5dyOfgqeSh/CalmwrY3hOe2dOoIl6Uzr6tFX0c61HxpNwd2y2lkB58idOMuZbs8uKnAf
fgOjAQUG1SEaiACja1aiIvPA01dqIWJAsojf3UhgrTvJmIL+SEhFOTG8bvrEwBQn7vPAWU1RGayG
L+lOsuNHJ5HWegLqQ0pBlwjHXa3vuajQMo1GbXvFEVWBMNV34vgj21DATZeVIPT7QriNmwJDppb8
VG5y/ggjAU+w1xAPeV9WsexMsaErFcU2W2o3edaDuXchy33yIrWVJbWezBHXxg7O/PowXOLBQyts
qyEnDibhnXsn22eK55KGJ59ThjUcy0wZWWctKR8L9EHNi/pG8zg4vGbwhbdDHcYf93dYTQu3r2H+
eYcUizA0CGKUk2VaT/On14vUODGTRpWWWJzXX9UXOj/dLtv72Bh8007lm+hmKwGWfIOU6snBvT/u
sjc2R64mRaRhA/Im+qrm/ptsHGwPPR8yTRXTyBnZj/1wewX7uBCjkmZSFOVynRzMdtytPfSMifU8
rIcV+FIjgQ2/aF5E88y9Y/7jPimHj47AQqzUO3qGbUL2F7Skc+NaPm+uKudZpQ3cLmFLZcvW6GTx
uwD99lD97cBxJ/4Di81mpJBUSZrkHT5kqLmJCXJo80mrxecOYgwihJXaX/3HF32NITyJ0P8rwpcq
Igkm0sNonbrgaHs1UkCppx6fYHcYVVNZXajzWzEaJ31G18uM8Qjvr28S2/H3a9pTAa9WDhCCk4hr
tE51WsewULDXfMD0tX/o9xetfADGn1LHNwPd1glJoUcwvUvQveLp52Xk+tJpDvLkLxx2ErRLMRcz
/iLPKC7cyJEim0vuZW9x/LKfGd8+FmVU3PFkumwnI0aYY3QrxPSpruPQ2BN75dFGAU1cRUeAPieB
BR5+g73AXCdxhFRjhq72WWuVMX8zq+TI1LXmnwRy8r8XJfnVEvceqT7qMfu1X2+0atAjEe5JX0Ae
c5zCDwVzyfKVGGCa3/C3CCIFAeBoSUPeu4JnB0DNI3XBJIPPqIEFbrpSd8zipXfAkQ5OXeYlsiNh
4Njn8NIixSz+WocRI7b2H77aISHDkUEseMvsqOxeRlBrXBshzkhjTaWYdMhLH5p/yVZqCHp2GBEg
/QfQUM+6iIOkupnjsD2yG2HJegKZ7L5tOSLlLToj94nr8OFnSQ5Xp4KSqkh15quJpomVQjoyfIy4
wgruBHkHF9EJjRbM+RXrwOfONazojagM55BIzMR1s16U0AiuoO74yNnpr4f2k85W6qRhMO4qhoXm
aRjXKBqVYIGN81FTmjQsFb+fg2bjUm2U+pyuBCqdGDS/wXh3BsRL8WeKMupRz9BX66XRkzOBI1Hd
AvhvFrORlH8XbSqbaQZAmXb18KzsmZJpRUhXcZbl/ubiWb8fznhpeqi9cl6kxRjdRXt4NQ/quQne
gLJuR+K0/fuuXji591Z5Cj5R1/y6HyusABz0aKCk8aToZTqVSOIIaJNCFK2LwX3pDFaxJ4FiF1Ko
ICdBryoGD7waMw+dZzogHdk3jDC5VeOSaQrxM4d0bNdda/NtqFW5ivmviSZ6j9pxJscJuts8Tk/0
7v0L4YeHkGiE3DLoLrHUsvyGTRIEbIJfmi7o6SiN7h1358Qxw36PX8aBB1nus87M3sygN+8hFDwT
R8YQJdwsgwrDVk3+fAYzLhQvW6A+Aj1eMZ3s/egHIBQs/eR48GiNSmVQFefKS/AlKeTmfcmjUEy6
2y6WK5n6L2M842gRwCBtv5TTmPpYgjf5t5fCHmEXQ2t0ndFjGIEfG2dJlVAF64s7aNRL6WpIJwk4
ZDP2WDexpO/jKcFJ455B4Pq9pDub3LUma2Ff0enfeR6H+5Ya0TEkHnpEFXhfm9ox5uI7AImFQo3Y
r+riaOGhgAbwp7bxtpbugidcnjCK3+Ay46LfxVB1LtDLarVOoUoNl26dTKQOtXFiCHPefBPGxV6j
D7ltTxI+5SnWv3V2lsM1LjSaLKjn/hq3uOu/JT0opUxG2c5f7lgl8oARn4EmaNjh8KoNPd1/VYoE
dUraesGynB38PxMCxCuqe/Gtbah4r36MKKLkqtLjn/eiqEXuSCmzUipUOpU6WUi+OvcbH+6qP3o/
+v8tIUoLm0Wi9Cb87y9eSTPuUxpBR4IJ9Heop/SQQ0gfgTZ9pS3m3vfGTME7sC+1EH3mEBNECYoV
jlUaYz+IcbC0vjqzezjLLkupNiuxp+mRGJAwU0wUqxqoqMgvDm9ygNTnt6wTBY+iZa9zCWhn+UW/
bsa08opOxwlrQt8p9294qG+dfl03KwAp0TWWw89GqdpULVjnvEWkBv2YAa8aXVKZOoLK3aL8E/gX
BV5Nc9ZBEXmMHrwSZWo1eG+VLGgECU+DvJNU99xeHBqnys4cKFg9cEbGW7Jm/befgGoozWiePHR/
D5TNL/sw3RFjFndG1yIJPnKxe4q0Et3u5Md86f5nqrrye3OavkLdhPJpCZRys9wC+BdUPTTswZcB
eaQXVEfwzRVhOxI6S5Vqcs4yBnRYD8LwXSu/EOgfGYtyovu8sTmL4Sh7AxOUc0eQQ4bItoqgRZWw
BH41Mlt4Y4Q38o7DjUgGdEfLpvzmIZDy5Ln6FSC2bO54aTp3Kg6qrfaRT6U0dtCqI6s4Omg74rJQ
6DGKdaISuWTvcCznISZYkop3Svp1IOC4ev3QU5aVd94D5y1d+ARd+fHST9iwAoaPsUYi+BkKAr0w
pyQirB3MWfdhhsf5rXFehrAp1Jx/8kxH0DZOHk9XPd/dXbxotDe8GGWYz6va24+0deh1NRySEI2Q
d3yvwoKPe1q/oA4JqNDocnjQcH7c+WKlxt/vpUTXEoj+kwgcUBSzzUCpskNMUAZFqCPHVlLUKe+h
bHtQNiy5iZZmb7Is0JKNHqgzGT/i1LYzCkgg2U82e4MzZt8Lw4kQmoBMYTfFBP6yE5LDVjA0fCXv
h0VZkXos8t7ZSEHh5DZ0oH1v1LxVjA1i1oLeuFtdcb3tpXYywziK2Gcx6/AgPgnmRJTcC0XKhem3
xpRUYq5SbpgcEBo9meCwV0HcYhaRUYGBJRC/eX45EvlT1GNkRe2q9Zc1ncF3E5cN1EDUigRz462x
vuwdx5vDDvfsbwM6zwrGqGphBKZotkCzrHLGcvM0yAJYLG44GjKYfSpg/ABnoh3Wora9UDk0kqri
LrfjBw/8R0zc+Pf38I9yPyGWVSxnpQUo891IvvxEHDvi0WO7HPc/z6iCWutTkl/ElKUJsLD4dWey
kx2ieVynNSmrZE9ATQoW85pEbUbtgFug0VltObwKFZ8vs7Iyc9TfMtsYbfavpuLCIDSUCIFCLCq7
31VMYUz61ewq5cnuKbSdLyANaccZsxQce2tGZw1/hw9W6+S1dAeHIfGxqmjJ34P4cw5C3fZBwzl/
jfSVpKRaRDMWv7CkeRXbQJz6cfHWl152o7kdh4if4U2sLf4zqN1UP3mPk3o8GfCRvpbViwCQRr2y
zr3HH2zxyE+O4VtXEoSqrZ7klC9aB2CNiatbsz6X0kFBgkjbD83BdzHgSDJOeaYbyibYFdSyYit1
yqmFpiGptN3OkNUD7+gZPotXH/I2Wi4mh11ij6cQcQ685C1oOjp+C8ExoiqOmc0jP6AnwrTyNUc6
78lEeIPtvQpS7mx8in63ITnvFPcQJnCHhX4uGJrxEWdd/IeTaf81ZF1NNXp1FpkFgimxirHZemka
klWGElxgnodz2FonBC3lpvq+Jy7wcnNKDBBE0qXCVke5gNtmUpPxVVcDAJK2Oqq/qx7ZCyyP9+jL
5Lp6dd92rNN9yA31JmKFTVexcZsgUKu9K+pf5PqQSsIyqZz9znhRLcN3QWqZqzyDsVFl/bWkDUoG
9hUT20R6cQotDOzh1fYYgqXmksjoVzLpbj9cGWAne/TMMtDADk8qF+x+IXMy628TMKb22S5jRQzB
s59PFPxV0lkeRnNzz6pfyoZZ9jzJ1dErEMGzJLf4PeVUPIUISqDkfO/eAJT+DBKNehn5rn3OWn0c
2YOTok48AwFFKMgvrLPjVHyZBLMZWs3jRKQx4VlzpzFiHe2iSFwalqIxk1pz/4b3O4y7YWX32HU/
9B+D6HBRDDHYhkISl57j/8OEo62JAE8euwDyE+4KiqW1FPbu8YfYRK0E2OlmOdbtE4JPvm5ysBBb
5mQY2JEJJ1ZcTgwSco9f5RGFIqRLom3eHSXYeGtdFsVi8S5cNAH/65Pa7FmHAAQESdFv1A14lSzY
sXk4+pXekQS9OR2gJ8AoPiu/G0TP8hs1s28pLFmXH1JRq1KynG1rR5pBrrmoVpZ2HifEVmgTSyO8
c58uwJvpJriX/ve6cnzEF3ueO6WOSH5UK6KEiwrdaMS2dVUB0UXNk2aDAPCGFnJ4LF7qceiQxue0
ifKchEpWHGIrlEeRK9g2sQQrknzcKzrd5URioTqlIZKt7XmYwx0jAe+yYV82ta77D4RQsdV3US/e
Peoy+Sa/8/ChW3suwArkgScIIkzR9P+RMEQwZoGL6oOGEwyrK2iC74V+dGE/pxgwOHVO209RFpQS
OoZ/FrRm9nLe+RF8ta+V8wesxDiWLfGb80PTuqSsO3b7LKaojNLqdZuH4aSng+S6HGnmLKo2nJ7M
yCRNwo8KF+2nyUwYsv89qLaT4a29rqGcF1J/1jcBrjsUBIjtuR6+irHj88+4QZ/cHUvO+8yBstGT
h+RYC+MaANWSnHqyx1HDj39v++Vq1IdrhUhzzYx5PsBrXG4EjYBqTjQ+FTtJLKxpw4lzeCEWbdss
7hbNMcbwI3Gyo43tjPkRlKs7JQBmMCkIer1Y7ThgFwCpVj+h4MybSf6Vxf7ZV5JBtgeM1K6TtfV/
7filMbmjoBIBLJkJTKG6ERWRxavGoulNSBy6YCmRmSsDMmfOztfpJXMV8RIJuC8sulF0PQasRjFm
aB2JPgpeBHZOF39v+Mbonu+MXQztePNrw9+oba9jdHZvr/8rIGPFfO7UO9VRbUwbPQrso7R/gqOa
T9np9gqfZJLKSgpRNSxCR2Npm/2ZapCRpevrTYXGTC5KeL2fbJUiQk5ZNTh/CufLZhrG6KZrr/Ok
yfMF210ukpkdM6ql+VI27T48vtDO96cFTC4KJDqyWSRdz3rPPIiqKEO8M+lnMx9Sbmxg8IWV6AP0
ca4n+5Mjek1a5PpetkmPEU+hqn9z2f8+yF6hdFKmh5YCHSYZpV7JuvyyMw6Rb32TaBflvaQMwSa8
LveIBtjFGIOg3IRrDF0uJBMeskf7KHGMnzmx5RqqEAMqBjPUQGrRiQhiVGuY3I3mktIJqfawgQpy
yVAZTBzL0EtKo3Cs0OimU5Xl1hQp9aN1JfwOVP0nSrdA+v52+s4M4HafmBVBNwoT0WvYm0tmSXgT
vIGF8JDOUGItvWOpyYt045WbOR85fwJguuHf/BoLtwX8+9c7XwP1rr7UPNjciZDN97TRUDnbH3B1
1C/aIEEF9CBsJYUXhFoVp37ugeN5OV1LJD64h2aDt+pEKQ7VLI4EkgjQwnhC+AMKvc9lu/QTwWdS
UZCyXUNSAeyAJld0uhG5D3LDqh8eEuragXpD92qbD6jx1sbkc1R84TFmQOTTLCwujBpqUF6v5fDL
00GmBm3yhgB4ozLhmhLodIbjeKm3lUV6iZ6VaXsxoKH1HD2M7dKed+NmvyHU6JzNUNynm8FludCy
dSPJ77sXKBYh4p9uVUZNHoBvBPv+RRANi/77WPgyNpEionwf8geOA/Dg1gD/ZUbMC9N/3CfEqdf2
zCF53cAEU9+S0JCq/KmUqr6n6WUoVlDl13bkQ+AqHgneyh1fdzE5QjocSeCiYNKEyCgrNpziiQyo
zHa+9lj7Yxpeo/2UwMETlp+MUY1tQaGlf4G1b57jdRdR4dAIsGzk+G5ocr+wQAQlIcxbo2Iji8ne
2QwLbOXhpbHVborlomw5dD8RFBg2CBUNy3mZjKvpZ6t932O1S3g+kVKysV8okw6qubU/65qRWoM+
aqI+SqLylBzu9RWEQgEOFHg9DQIMcLBCnQtDwt/5NL8p5MeGP2aMfEWu+Ewdv3iD6Hnuhsc4Gjvm
eLSJVlUMlYSrpq0nci7n+BUNOs3hBDioguX8z9riFnTRiXtMZc9CcET6cCFG7/pqVRPy8viVqS1q
il7O2HT9mobHbIoIUq0v1gyFdPAlTwK2TVFqjQwesx0xz14qktk1yzJ+UDLrObSDMMJMr/gwTHD2
OBiKZVd6Or+gZrWTR5j6mco2kAm+zOzlPZD1NJHQ5qfpm6yOS5wso6wbr7e/He7uU4WT5wnofET4
hOzDVTWAcZ7aF+exRY8dnb6WGnap1dRvA4JfpCMOkC1AzaektP8B9FQ3ygm5XBU22mYrXIa4p3nn
k5hiIev9kRRZYaBEznt6dvbPOhj19ttOdZzq9Hb74YPRGyrxkrVSHPE2LGroi0W33eGsiYcfm/6A
rmJH3gmYBxKAzzl2ytx/alpwTCREeJknQWtoaFVClm9Rpmmi2O7mg5AFRps2ntzXnYfAfP7aq0rN
cgdIo2hn1FanVWrJ7EL7+k/jrFIZrfdlEVQtCFelgcuOZZt6K218ndTqkDYIX1JgxCuPb/KKB0DQ
Dng0vwcgRQDrVHfuKFiHMEomWN5gNw581cU5EcXFIQyjviujW5SNadcyC4su54/+UVNrNuEbbtCS
e6iD2VJ+VgevcVF4GEEw8UOu/dVKEcmqu5RQoOfROnyKkMMlLionVcaE3QGxAYMRvLd4ywart1Er
9zjyjF7WFdOoAj0b08O25wsnEV5Q33+c+kIFQXby37f5DfiQL5teOQq7OKqjJbL5QmsMHz0rxvTp
a8PHtFAgl7eZkMOnmeMj0fctf+6NGPfNriVMbtpznKl9osWvJVt+4CS7dN4IqCsZgd6p/uOJUpiI
hZTwzyXzykGBmXljHVRROtcFMWjuCiflwit600reY7SdDU33wwzRKJCBkVGuf5gDLkf+UPYkY3CX
c6zhzCG7QptQPlH5bJkfY+ZGxbIzVrjvZpfixpiHiEXHkiJ0zPGePExCWe/h6W4tcPRTUz3KzZQW
B/1vloBrV5TjoXXTB9PshGBnlVuuLLZAphknZR3B2VrQrXRbr6PmQkOKDjaALQpuQV6YMHOvyCe/
4xYVOtjEMQJnKwmuXsXLfUVI1gqRi8HIZNgd5n0NxIc/TNyWvRM+1eVRi0e4AShpfLgLUZ4pJLMs
MZoKEOD8uXDMKnGCmFzDcN7d11XdJNWYj5sqW79QMyCotd2DoDIR/dXQQLNvdZHYKwMlo/h5VYX4
ycspBTFoY7tm5+gLxXKVwoNXNDaSDT7lrcLaU/Whl0L4ppfL45faVAA/1JRWL4wN/EZvHGVUhBeG
Ug14qrBUp0TRC1sr8K7W4OR70u1jYM3Q3XQv8y3C7H6Dj1urgbflag707r/RTJCrxtZ8kdAUfjo/
SPSYhiYSW7zUxfE6lhI8OgfjPmRMPGHDTjFDTh70ERjIHUpnqch8zny8z5mv6wP/WOnJIdufAYwg
gq3sGId9CX0lgxH52VVwUeK9JNskJb1e0FQAYlB/IXbH5fMsE1LtI6ywon9SGDqheTuasn5cmgPG
DYD092cEhwe5CL1G06X4IfPGISKqQKea4m0frHQRcfKZ8PKjOgherIMAFLXG1ydVUgkDD8U+dwAi
wziU/JGnU/35KBzZRQhgc5utE3dAZqDJgAaxIWur0MPpMR8wG6kzOGPU0y4t4N2/ivFOAiwKO4v8
pn4X7ijnpSekrGKch/4O7l04zdcDaWNwVx74dQIY9912j0YiiaS+ohBaHTAAuz/jloIQxHw6EOpP
WCPnC9+or/UnNk0FLAa3uQz11FDBaVZ0Jr/ctpP4JwiWi4AHvfgzvqgNhx6b2yYqMckSaHuzPiNr
ExqHRbpXb8yAadmjRuk/jO9Hq0HuBGA/JnMwOmPA2TSJfFhDLK61ic0QCW638HbOjMnk/qHgb5wK
QlSKK1xLuAngfKU5yRw1XGVFUJ4/ZGA7RJjxAnJPmj4WdsxWaSs0qCJY+HLcVsjICgL1KM4sZySR
1iLMsoogDdDDOVeFnUFguehFlQ26bbDWwVBAEK+zhA3SCuzClIdymsHGjdQBPu9rOF9655IrDfjG
pgwHr/E01LDgyw+yQp9FS0zgLVT0RES3GMArZ8XmZlhq2qPTwiCjq6DA86HqUCHIsrtydyY3yUjc
0XdLDEC9gwNIDktigM+oRvHqtjrmjJ19fCI4mA2S7erbJeeZ76X+fj00t0v2h2gcM07GS5wZU1Um
DZ3TPk8bcxuPHPQazCwEi+zsfGBAw3LBvujp5vH5IzvkO004QbR0dbia4n0HRLjFRqPF3z0YV89R
fQyW1L9luWPzMMCXObkFYhRgZBUGF/L5BZW4rfwyU6On0YZHaU6Q9cCIS9kvQgKL2nBKmdwBXiPG
TTV4heoSnT3MQ6DzJ8gJoYdxgbFqOOvYVKFmOTf4tgw7ERdmVQg/+50anIaAo6jGmGNZODpB3S6d
ulX79Y4UYnl1oPhzE1s+mSrBSmyvRvQyisRHg777EwgSLRadDGUMqiC4iz4qVfX2xzdbix+a7P2+
4E3F0cWjAKQLHZagOhh3z6y1z052kVWLjIX7B1TwKo2xog9br1F9Px3IK7r4gXdyyA+m8UcQU9wl
GLpz5pqhwfsBnuVsusAj/oUFCi2ma/mvSDszcwTRxXV4kDtfV2oSpnlm6TtE0ZSbj2sFc98aOhdz
NSa60jedVIG1+E6H0zp0zxuzpUcVYSmquw0Lhfo8XAOupR9pN02GENXC757XtEvuzn38YWRne327
BeOui0U9CNPCnFtAT+nQi63CHYKdo9BgcA3S8atvwFSZ2FGkOVIdr+Szej3GjVMK8ezP8C7F2mwB
YGO+RAdCKlgBwzROJ5lR7YUNdP0yoecxGSFVFsAVYatoDJrYP9R0F2fFAafdgIVrhrO9TxynIR6W
IUtcumcUO/BcRgH6jYjG0psSomlEeN3pRMcOYgdI3a5QO51PUhQsXfCo8NOZ9FsHpNoLcb9iwaxp
FdD6e/Mv2qPx8rWxNSYAITV2/5ilXGacl/FGyP4tXnTQs4Vu00aB807xvQ5LxGXEby3QDZRBVOes
+BnBEBxqeFAs5IgUSgUaIOkAn9faez8zYmLGVOKuxv4QsNKN64owsqwoCvud4le1mkmE4/ooSvNr
HFhRB4Is7eeO4/LtZaRw7cFKg/uSwrKekXhUCWoPUd1ClkWL+0gbPr29jfPfGG/fl5UdjdeIMYbm
x2O5FxFDXwVHigyI1pZCmv05j72bZcxKBZIjGCkY1BLQjFO7ayGFRrxlWWo8sfEOUMNjDJ93BreK
7g/Pj//8kEWXcyoGl9yZ0tErbqBN+NJXpzOrJb3JoUW4ZDwLbkoXnMkD0uhT4hJQ9Wh1PQhpfSEp
aAWggmSw910ezGtVv2aKdvz8kIPp1ZW5gXRmfHKKcC2+U8NyC5iCBNWe51SWP3qhpBNyy+ZqIcBr
c74lDCJHHqYxrbJsihKpS/pbCgdKVEsnuGqmAP9fLcE8gRsFV1lhizRmOiDcJHHJ+64ohl6DrG15
jZOpg00wpLuUjEjgJHzy4nBigZGSrCKbY0YU1oxPDtxSVswIUrXzEjawobDpJ5wD7XxzKWgOx5Ol
JHhjqdCd6Qm22QeyUn4IkST4qE9EyzzfA+zpvHJ/KPd2Ynpg4gvXVkM9d/uv8e6jsMC6PJnd2DaN
pDMgEfu3Csx/wGoicmhOtnXj6sP2HAuQjH5nac48B4sLDIDuAZLYQQjkYtoUR29YPiUyNOE6Un04
Yo4aeZ/UdOhppP6jG7WLfs2P6SlrXuZkIEhHwux0N0ujM2YRZJ2rxzaQf72doAahv9/rYvSSUqwt
lYiw5MII+9pJncCYqw5gkRNCwV+8TCtRNDdd0tjDkT7SUyFK/LSdLnfsWdXDuLAfXt35w/CdD/64
X8CvZI9eYEaReBnnOW7arPZZs8PQmRtWSHfSiRUdNAjASiKjiBwCkDtgt/ws62hvRrLqzbIdnFTX
p6Bq4LOtggySjXHe4ckR29QOPSokzrNGWFDK/Y6gKeziE8FelCodU556Ys4m11t4cRZkIDQK/I+N
WJA7kXQVNZZRKvmkEiPB3KraLbbqWaHwD+aLRov1PaB5bPv2cK9P//zwRKw8I1aWMn4gi2jkVBfk
L6eOA+2mYYoZHMdPkddnUWXML2juzcnVe8ftpD2WwN6oy5B97lEdUiL7BkiiA2slqLVNabH9+3GU
d81naLptg7OtmVAjdrsk7rvf04qbOieVTPbjBaF459IhSN9/Lb+Z11XmOBbSktzWNPYf1C2a5d7/
eqf0KMvBYsAmAtYOAVDEkkceS38DJgnjS/GSSndF8B+3D+vZBfJyt/ZQNP2HxOWmHXV/mTkvIqWv
BKwLyOOVsItw6H9R8KYofNqaH4u1nxZHNzz5K75MESfIwQVSCE3RbhLzY0NAGVPxFWCsVid+T+K/
308wcHuPZ7k4AnBeJB2vUYQnjlfsdD4oBW3EhelWwjGEg1wNXLcwtuD8HTCuIylY62PtcQz0qkc4
3vL2TAypGM/Jh9W5PjaDkvf4n9JfuF4qGJmHtxWa925mjHUWsgX3MJ4FndNjmcLs6yMTxi89sSgo
S7wqt2GXtug1XovhvHyWRE497ZqRNqTps2rZ37jlWmDy4UdhE5D0FQrtQDbhhBtaJXGVT9H9sHEz
YXCKJ7B+PDG2xQvlm1//TdLBM0Lavt/QFc+AO9+1I0Td5hHw8hLXR3D73zCZ5a8K6Y/dgTkWQl+z
FXXxhOH3WZ+qLUNJbvrwvu+HcuWYUXd1DOkI0FlB6TwvhgeY6SoVwbejxeBoUaHN0uAhnqU05s61
xjcVrflODi933veArsH20ld6iqnqNzf/hN5QNZLxeWkMlXR2VZg1RPCgbOvEfUa6UZevPV+9bDOT
uytSDuXkEAfllYk6Y7P5GwOwL4wHxvTQAicaOsCznAMj6Q9bt377wfsXXH3Kgimrc5YPJZLo3J4W
xkIfM4FFVxbnetApKvH+t2nNEf4+O79rdEMUuDp/R0yuvOy3xlVhBAUxyQFV6amMMO9A0k8LSk9E
ZCTxmX8PgcEyMnie909ggo8UlKemKI0Iegl7CPlWkBSOJsHoFGkZ1O2Vv2dITjNgpdKitTejaymq
J2w2zHsAwZgkrN1iBUsAyyP3Sw8GKV6GvB7R68xD55D9HUvYN7+fZSnyJM9LzC8FaSgM2Qitu6Zq
tplgtsRYzyGrHE7Tqq+xpHOprEtrNtsh6b8GqD79F+a0Zcx5cN3bv9fE6baqT3n9yCfMVHawdNYk
t/JiTt9ybVM+UBiv6L7gCeFim+1YzlGl3hg8G/cGugmC2FknySygUAJSxTNMY4eNzN41J6if8GyD
8ek8ZhhBSuZk43SMVtRCz3E7qcFsTklxl3CFzln1M9elLKkS8bDqWCGsZMX/7NZhpupnnQauuGkb
e359VTC1h0p1WhpMhhheKyUC1g2UpqSNvzd6lG4bZlmqEHYzFB1qwDi5YW7DVQ1uL5ZNAiej+V8E
nOxO97/wGQGsRATKf/El+NxeOqH1f0Udv4NNBa3/GxeXRmIoOz0nl/QikZY6NCui8f0wSf+/s0No
H8AKLfw/10sB9JG+P4rC1SjMUWe9icIph7ElAglQEPfI6goObI/Jybn+CuLX1BuWiDBTtj2SD6ah
iSrc6dOGAJ3uwwPejpECxPOMXEOoUROTR432CDLfrVf6In7pGESNeDfLTCScRWIQqsrIU9OuBUU/
jSCjNfyLqzjzSpekhBKXFbHTkmwVFjw4nk2kavsv4e3IxBd+1NzAxhInN3Ejtnu7oF16TKUuEm94
2N+gL1NOWWyV7goIfGdW8Pmojl9CpJUqasvWfIyGXn5gbPaZfjaypzHyrFtLiajj33rQzN1UxYk3
X2Dli//QgG0sukcxeFU3eYlGTWWlCDam5XH5+JGcZqEs+dCkNbANOHIunt9ShcMwTIJz0tjPBBsX
WfDDmcF5sUGEkUO3MsBOmJm7nXUtVD8iVqOvcCYFw1VSCvXanXam+lmdR23+AWgTwKjyy6QZlDMg
f4o30fLUJXp4uvyaYs9ssIBsuMXLD5UPYkBa8fF6Ix2EhQvlGtjYNVJPlV6EUzj0VM06HefooTM5
KcXftsl+QsJVWMiUvftPQ3QSN6rHrGX9P6/GJfi5xOEY7jHquhw6FoWE23AZpCiYBHJFRPnp5+E5
Xjfpw2f/o2yKiBeZ6nHBwkxtfgEd9b0mLiJzf3uoSyZBg5nizp7dSvPK7E32Z3npAqgLbo6w28dQ
tSB4YkIOQ5Ne464P17TOndiQNKFiZB0J+KXxwTcI3oJuru22lY5owD13AvNP5v6lZhlewL3dUGa+
Ebi5Wua+q/UZn2qBIwBoWVSAG3esJrUPBp3Vqnwm4E98pJK1S63QOIDAhmHnGTqHe8Ud97X7z+dO
EFrXUQLWaLfo4kKNcYB7riZqEPYzIlbLxQwthhTXDWcRNjn9MTtvAHmtDeUBYJn9oGPbcX0nskLu
JgX7N+v2TGGd8EPZN5UIg96fQOLL1/y6jA85bNH9J0OHz3iGRQuSeTZBXK/scCIjuxvKf9LESIrs
Pr+she62hnFHgvVBetgMj971d84JOC0VkHa6SHdFlXZMrVAzsDBazQ/qye6dXswOyfbvEqLlxrIy
GJRrfStiKRmYzJ8YTFVljyhgh32u3OW3MVt0b4uh8athnOPMF1iVUiiieijts7RrRIBmsiqsNB6w
dV1VssZlFm8+wjOL8RNcXILypRkee1ar+HK94/O6M4mPW/bKfiEaITQy2wpGTV8SOk8lZ41Um/7P
XQad68+nOSFarCGpdBt9tAarcxQcsA77AkoNlgOCvAmYo7AkxikeRrWw07ZxFD3MMcqlOW8jrLjo
ZXLJPJupk/RhPPFKNJN/3Au/RFqI9B0IiT6YhwIHTCXAiLH3ziVSjAFU2W1oJ/jYhIvhDUPSxa+e
JICbpLBLh1/hUVR6SIlnxWsLw8ATKo70MnKJg32VR29iymgmlte8JRjjCrxZA0XJo6733MoCEUaH
yXCtnESmLhvdx82JOOJXFP3n+YrnlFSkRnTNFMuvXkSjCYYpEC9sW2ePFys9TyLC35nOZrLOachZ
z7NHsKj42tQ9pN46JEUsr0fg+ElIJGngDuS/6YkERPWuWNt30QWBoFmlUZqBHkRFF3GQK0cCT/nK
t/n/binPCiRfhbMW80mhLzTxsykh4+BtWFKWzXaV/++lOPHN9sIv7YpSgix6KDrp5RCRTSXnLqbo
K5XjtFV2LveqTjoQp/M6SFPvvO0bDnFrs5GWL81xlqQ7lu42kNHNPT39LT66pLYMIjJdP8eG77sR
NTfuyxNfsBPptbYVqxLOABIZhhWykv2sM9E1MKHQRhsUAthmywpjY7DyFXml0jw2Yvd1GrXcMAal
U7EXwBcuxOf0DDI0EZWZT7Y0bpI80zRaDIXyZMQ2s34nSnzyUCHUk+RSt59EMMmDNTW8r1sibZo2
hcagEMU0kCqPENCqwvF1cpzlepDe5ZDlP7bAcW7+NYSvDEmLT1AZtymgKvx8rD+hrpaXIpqBIra3
kREEJZSiLNGA/k1mwgdLjPTfLknvVbrMVdWvISA/4cCJ+9g3dSlp51yvGVjSbdzZMB8OVazo4JOk
++yny0wmV+JyaEAcQzEF0LStl8H5Gv8kNLKNyLaDom+PQKCS/R/8KNrSiyLrUo8aPDwbGCt9+C78
6fKqg5tfpIIoG5ziMH4/VSdCSfMQsvEwTJoZInhfpmmKDXHs3U1Jr482L0b+kmygVplx4GKIaLAI
WJ5O3Pj7Und3aQiYgyZnQjHsgXpEv11QdIX3Q7C6IANpRxLKEdf3W02ctrHN7VYI4ANa+44cvBr6
ZgTddrmfEiCMw8nnFBkV+rp9s0kvk4FqWxAYJIp/5FoTEikAuxg3oy6j8HRosxourN1VwAIC52Yp
RN/rt3CCysEMMDZF/8fdUP5Z62+QDQUH08qcjtvYNHhZ4G3DvW6+pjPiZy2RaGA+JOdBr473KeE6
bQjtj+D3uWiQ50I+PlqAz6ZbQWXwKAOy5YAPBP2HdOiExA/UJ1wjwxadC/Rre38ENjQyok5Fs7ZK
UExrto3TG987GUwxi5BtFDe3Kw2XE/PueOtz/E/Fg/sq+6A6xe3Dz6bHQW8FGEu0teYpxFR5QIwc
ES3lfqGtGBLHyNBi5POfUmtGr2fzhVz6W+5o8Ma8mjmk9hg5Q04c7WBw7KRu73ogyfzMq77Dvvuy
ewS49kvFvLGCj4CiPvCdVmKr17OWweIUcspWRaR+ORaRUCH6zGFJ8B1j9AI9jMyS07tULDviQeSy
ZXIHZP6mSVHBuVXfB4LMONigrMBAsRnTSQJwjLQi8YRJ8bOzfJj6zqnm6j5FgVLrusdpneX48gZK
Fz8dVcwVC1BnMzxtInhKDmvKbcQpHpmUOKwjbu/BlGmNge6fpwIkLrEUV/+sLeHW4/MWrngbxI1P
u6BixQTKNjApwPAOjE0R54fMs2XIMkH2bQQY5hL6eZwuWNwRoYfmoRZARQS3+w08u8L+87B4+gMm
iGVVEbLu5pAUWFoKIdb6sJKSZI5MkjFhke+IiOoGrOMpAvw0WooxQ45T5fYn9aHtsvuGXpRHhkps
aPTITZC2G1302Jfoa5+ySfEgH+USdUZfHEht8q/j2wy/e2LWKXqvLErQtXR2LMNZyuTypT82X+bw
51rOEkcdR3x2iCZ/U19Wscvtr1Sbeb1JxihkTeM32RR+46chNjykumKqzT/e9EGOe0Mu1J3RNCMp
gpyeS5OsejpK6cvXyUG/NVYxmmeO7arLU+tT6p+lZB/5/LycuLaGhJ+F29PfeSOIVLomO6mVxpxa
SM4gpX8kTa9HSzv6naE3wMysPbG2MR0c3itPA/H7CaCpw+7sMaj7tYjCQtUEgEjRk3yMKJRyxNbY
+zH1+AO0BYcMp1NRcv1X5w8wcm79/Am9WHQ/KyvgEsQTGUVSmi2SksXSF7U2Qv+z0+uQCnyaI2BU
1lszEZk+yr/gymAjoIarpl14nmiQZOCFEIuqdOHQyI45tm2vWQhgczP7Rp1lrgSEwE764sT8nLkc
Ke3CSrwrvyfdKjyQu82r5Qzer7SiTTL9J/Xq92cXGKtYKBBN0FFabEwD1Vv902ch0/MWb28LpEq3
8kYSMKtQmVtw9JmDfHcGSe0saDYNO5WxM+IzkFayH3XWXVJBn7zG6uoglIggd7eXddgQPGr3az/d
wFnjkSVkuH8WJ7fE4Uz2ij3X+w9gSUANgjxuC+UhDsp8gRBfLK7srUhbCukktHydSaZSbCMXRYkA
yGKP3sOnOI4dSge9v/k2H8amiYZ0Y/KbvChflOo8JRroLxLLfMmGpZvX7FAIEHOzOCmbZeG852d4
VWGSmhwR+nDM+Sw/iNaS1vYHm8da0eLXIJfmTgEpxxPRZG8IXkq9Y/10uHJHhNEM3u9hAbElGfmu
TLJRTphqLWCXWuvcOwK7Z46gatIN67NHaa4jSLtf69/oHe0eWoO/d/MoyqqDxMWnICx52wUipn0m
59euSq3aiPNhwtnlK4Cy96CO3rpQR/d4D9YV1kk5el4LIy5jwQCCTsym32MvHpEGCE7phST3pysp
UtDv7H9Tpc4zYcqfNPapuzBR+muXiK1I7ibppoGpmCa2Jgl4/ZMI8jLQFsInTTWbbAXcqMSJCbbO
URQeufFrICawCzmlPJAtKoxlSJlcsAEmn1IrfCG16fWCeKpAIl8BXVRydnDlhPt4Q+bHlxqpCaUF
KUsjAQLB1pCVpfnxg5BE4qyFx2bWjGq67kW9kHTBD4wtm9KGPus7FmnLYp5I4a3ojk0dnif1KhAX
LrLYXZbMkgOk2/CINwsSBNcfTvG6Qiu98IY/fRVRxkdm/Mmn35e63RGdeKdzBUiQE2q/1qJ211As
dhll5KmfGH9ZGqjX5gQcJvqOPeCO7kTNNVjFQx6Z/tgaEPNtAWLoGUCH7veAqR9/eonBWEvgx04H
mBEi7qi0UGBdpgtkTSuEHcUR1vzeLgKVg540cbxJSkfzj5sH6OG7b6R8gz/LlcuZQLFBo9h+/ADL
b66PPgZL3zPkgG4cudJDZ1Bj8oqj2Ll8zmsuOyzN8xejli7zUdOcpWnJRAAAos6MieBf9LtZcGH4
GKz5vGCnDFjVOA6NvDOOFS3GyuzytSCPkUgTnzlCyLymlpomjO5j8SGLO6ik8i1QbRAu9yTlMfGj
KpIBRpYDurcOdGXLE2cP6uA0G2mEqMHnu2l/GrDa9hJvUmjbtUIcdexXWZcayaV7MsuwLCuBz/Ny
yLMOo33vPh2aiQFdbXgts0KzFKw/grVZUjZM4tShS6EsQgm7690megNGV2e5r4vumLMrznR+ZtrR
MxqZS/7o8qZg2/ucNWe5G5ICsrj5w56aGWSGnwX8v5vcWUf8y53UmT3+TAjhrltfcvKc1g8JBq36
Ui86HlCGrBSaraeHtvubkqtxrxXV+MYoMCLR9/x8gMufskFHyfTtaR9L1Y52qTLvoPAi4d0fVh3h
RhgGfZYmFMkl2oG5d9oUcvfSm+nC5d/qIA3ZgN5IuIOniRwzDPlg2Zvy8ODC97qqyxa+JdU35smA
j0mtWc3xKcJHB0T7ZaVz2S5MPwoIbSd8vkKhp4raQwMh25ucj7MieCD6l5YXw/YOKH0nTLaJTfNP
yXmGn+zk2igwOfNZXynCci0JfjdDqCLH6YRxotaNxd5at4rgeigDHxKbEOCsJFmBjXC6HT70X+sg
aAVhSV9c+q1d1IotgJs8Y7I4K4E7/FxBcDklObzSkeNuyA6vUDVxDbcCI6MsmKI3SSpLdaZMNFjZ
6BX1k2q2ncPw+p2mIPbUJMQ4udrBc066d4AsYxkhtxfmSW1xsK7MGpWS7V0wnQ8JpJ9381FDtHDh
Mqy0xNDJu1lhOJO1pyLKi0oZt9QZr3XiarBpHACaoNvGilISvPjKWsSeMRIEGLPMJZULnk/Bwzv/
cTqH4fEumoU1eNpgx5qNB+Inr1VH4WiXQZ0JCXe846DJY3GDvJIbRGArfOXy/ETzq8U/7U941Zt6
C9Kzz7KnmjmMyir/8Bw592QBf6WxHCGUK7BEu4Tz/im61VQ+6SWxnOweQAlbGl3wWQPBM9k0L5h7
Sj5q/T3/WiKx70LRkmyVzeSn3lYfgNWsj1XiT9+hXEtZjJscEB+TqJrL+PHxA96bo6qEVvPff0JT
PjDdxMZokpY5FL89GEERyjdSQNkilSzh4d2R049LRjwCRMqY8Sh+yF51F4NQuzvMgqgxtICgRKnN
6U1pcd0+B4DyQ7ftpHxeL0PDPanqzNKfO5AkFbLG3bUeVU0fWGQAvNjL4SggfAJm7mNpX6Dl1e+d
Lpa17zr4G6Ksv0dJWzjScxPG8H9UGTVSGP/AkO/w5h11xMMTa815xUq3OSErU+x4W0F0DqoZHvae
ZQZnoqZ1VtkXKPj3GeIckL3CGjZ6ENH5G4b7r45lj3LnjJgNG1zaPFWcvn10m+HKhGQwk0IVVAB6
rKLyOM+sVW8cgnLcgSqx/NbYw6dqsSwVFEi61qCAbRepZDWoTT8681cEFDTEzLPFILwegwVlPk/a
voUcLsh5py5LP+WWxxBTrN7MqDB0UUl2GovG8Y6J8I6l3MIonrZtuOsVdQeQKq4c3pNVz4aJLARc
Mi2C8Rimm/4DVZJOhnaADoHbMQrjrYj8gvsWbaE3i2vPVvmwWS0IZ6V5wCXwQHZ97SKwPXwZaskC
rCOEKpjpFu4HSNYiurP0t/djqGo48pdVz0/axAYPhJ8vvZw+ltwr14HrsCgDrqMnWzUBYlJ0/jTP
7o3FUPbRBA9aaLROivl90cdo6XNvJKc1nlIYcIKdOaYDEEcl1DG6WXX3GvorjKqnmfwd7WQzkOvd
ldu5aeGxrl52xKS71eUX44XsNMnCT/H/lwPvPJ0RcYCZsNNt/sgZWZ/W1asN02Qjpo3x60HimDSU
Nj4tNh4PwhCmdNE2XGxUVVmkVyMvZGKtBT7SKUEE42g+b0ZMSjPTGuNUnbufogloWIcCaOyMf+ni
RIkUj1B6OH+d34Omge1sNSbGHKID+vT5VxYFgNy7fQPaPYb0B+KPa3bZ+NPUX5dMSFJAQoRKcDTW
sx6OZSJM60XbqstO6J4sg84xFJGvfzp3wFCE3OecBU1R0Rf+eiup0/Fy65fISDGrG6JyaZw51Bcy
dQbWMCCXiWzaukoXrQhwrN1flKkbIRHNdSprG+Y42FEgQTPYFx8SPTKyeg3SPa5uvTamjcQ0nxyB
JTUv3XhWcgegcMUsqNDTfhajH94tjqDEpYBOCssE+FAOjg2qdxOZzt6bqWtwee+xLvMPTOZjyPHp
tG8tmk89nzDRs/Vf5W4abK0FzVRR+mgnjlAPgbucc/9oDJWCwp4To6jNnEaBLeS2Hni6bEC6f3nN
c9sK8f2uJceKcq70pCMlG5yBU3PURaqRwMQaniBTbi0ABN90e//JQDr/XSYmiy0P5BQpugxXwWpo
f0MGTgHzDomffnQ6d9U35S6m84E7PT/AqWJ/99EijtXAA2v+5MVNz6ZDwfVN7kxE2D5B7CBEnJl0
VlZLY+DpDvqxlUr5AzJphnDNB4PLU2L2JBQ7JpQJP03YmHCsKr/zy1Q80CZcIuaxHQfdFiGKmSrm
nJ1TZ2pd6eS7fiBi+7dXIPADmM6piN45CYHhwOo9+5bAlHkhTRSc+2Iz7sCFA3qaf4b6vqV8F6fj
PBZ1SyTC779Epk1uQNXMU03AZjp++dfVqUPMaIr+ptNCzpwoTuC4Gg8mPO7rWEFdPBMyNoekbSSH
em/NlwL5m4tYo/u3DwfLPsqyvzxoYHqI2tZKW929kGas3zi3e3x0twO4UKjCdSyNmjN2A7ClLCk7
MwucLLBpEGNBxAjjygj2o3ICJK5CibjHL2YXZnO40ZBNOIfZcJytHnzHjfctcn4I+T24tmqgED5a
mh5MdWrvqSnhqRqllwP1NYSSHXXyFam71cYteNdJKcVfk/3OhxyI2IBPUOxA4XGeGZmKHiBpsB2s
gq/5lgjEhpBDiUvedeSsRgGAr1WpsfqIKGGPWqV3yNcG5bgrc41WXKqjg+Zi+vgVhxi+JBw6si/W
vdMRwaRd190w+cdzJoMb/0X3U0oZxYAnHfRKI/boaZMP5G3Y0EBC2efDALT2itkAEszx4X8BfNgG
/pT+n3uo71meo30SCnT49/JFeeh5z3D8tzOmRv4UPlOGewwQy/fHYmJIS4krDB5szRe9vw6lPQet
nhN/K2L2zs2F4ivwktIaO7dF+X3/zPU6dEQu22yTzfigqCSnHhYS2JasmUHXo6ba151mZkXPtZT5
hEHv83elC0uLubGYtDVjgBU49DoCz1OU9cfxpmyDICaAi3nudUUDzGBfWJcoAgohVFpggNNRY84V
kAu327Lp+a5ZeZJzeo2Bu990y8JcbCwUxJ064mz0V8nKWpbJZY0kHkKHwnqmFAnkhczW5vAl9HfJ
MdZdMAePks/7ZLG26TSleDlSRYozWVx68Lp7HatAhCWbB7gGSzQJ9Wydq8Og9eRC6t/qrlJehQqx
/3cbN3aoNrsMU22EO5kr9myhaIiNkdUj95q5VO5ozrKaFIonC8RcAKT6tyW3OW6nJXkVLN7SMo35
n9k0SZEPEQxPnLDslD+8QkVoE+MG19JnFzdHEYDEhgJSooS9vjrg7PghE2Eim1HF4PtfnQL2QP5A
2hzeV2CGb2ecxOmVYXImJ/yZ7NCPtCmfnjeYN+bGN80SEAUzpu/7okIm0AcPfccT02wMxrTJio61
32e95l2pV+Zb8AwG2eM3be5LZXytcjMWU+aus1plHbPte/60TNS1eWZH6U80LmiWebC4NVG+6tbd
7nsb+xCOFwT1rcSUtsEV/0owJDXteCYNlmevP+G+2QjdNvh3lCnUUYGSVusQK82hDGlcOB9KSKev
rLLUgvIaeK/kfCDJ8LnA+vxcBmkrDziZYRmU5g6LHGQdxNq1YD87eQ8/uuFblb+YAvm4Kf1tRdrU
kF2b/t26+mRzlKVN9j1XylyL1LBLTiZwSJBbfxDDklNgCmIiiUpA/4bMvUDaeXzOhwwgfp1pyX93
mMLWaacFm2xWQaFYSDSY64jkggnleXQEkSnsjOI3i72m81oWEGOU5ZzbHh1ZKnbk82GqPBtmwRLx
DOvX5KSM6bdP5uA0KNx935uIw+yvwGEd11JpZyY5Kr/NbCFxTZMvBnnO7uu4uGgfxgHLyx2aXr3c
CA8IA/tRrMXUkCZ1RotfagTNqkAUogu4GehzSZv5Nf2FQYivrzeFW3KNlrvggOl4gIPP5qlJH/M+
54okd9Q+9TsE9eUztYlPyA5cgM5jrmJgfslgC70Gf2lsP+jR3ZUSAysbCz9nGaV3dTdtvW6nz3EZ
qH5DtnFV2xPR449tyDmU+D5N6snIH3ymRP+TvvOPHSbX5RNYpfIEZ/t5tDgy3mOwkSxy2pbJYEEY
LOT5fn89VWRnOc0vthJU3//WjuTO/oacCvOVg3VwEgvMUe6qEwU1/myB3Z++iC8riLUDkiI3eSHT
BOg2H0/DDIdwxhvPgqFT6xIKKanxd2QDpKv4yjrK5ab+zPflu8f7jT+l+3PUfmKL26FudtLpqadM
xF6Zp5Bp4bdXi5VcBLd83M9flC4lgjIGVCx3HmuUD7efF7l2jBLmrwmmzFR+dmz9RZG5w3bxPKkf
PawQzAPRGbaYuCUrOCV0ayI8hl1Sb5ac/g4JpV/ByvCXr/mVoAi90iQLz9aa7iqnVJcFYvYE/Ct8
cnIaCsxW6XZKSchWuBvhd/w6+qDhGsUtF0zeaO5c8A1q6YBeY/sc2ln0t23Az8kAB0mwgDE0PKCg
+uSBHK1yXpC12FSjyo2MfzpKNzwer9HFvz8m1wUgWYVtQvOqn5I05iRryeOEk4NIqpoPyRWEVKHC
UDZUYaXW1BUObcFaKEXea9lf4HrhYaYssLyfcJ8sNbu6ZIAAiFQw2stbUeTUWP48aoH4BsgzLBDo
KJeZyfV89G+GgP1T70mWrlpR8lGo1slJRcN08GTU68F19y91SlY1c0SJsAkP9rN9DPGdPLh6sf4Q
jpWkZxmvn/Esq3NdAg2uvWWS+UEh49XYm4Pt7482gxpTiBEwnVRt6RZhFJiRS8dIPvn+2uFgGZrZ
F3Vr57aZX4drONBhV6u8tgSM9ZTy7nsyWNGRtrRyhUIE3UbF4zS8VdWuzvdJwStOthU9IUyXbMZX
5WLC+RURKVTA6FLBIhTLfyh+nSJo48ItBzwIhDOvd17B6ETwBVdkx5oPVfBwxKmuy7RfkVp5mcgo
dOkIABzRgreT+d7sgZqxB7jzLS82J36eayerMpM+zz3fA5D9QrBwcPmVCS6hBXGoCYNqGkU1yR3Y
vDnlTYT0svxZkzpDsk0cmPvlm0LIMifxQGFXxMABCnUT+pgPPeKI+IMWG81DhAndctD7QN6UH2/n
rkzDlCd0YWS5h40VUyOPdww4yN9n4Mj9dB/F154cfWMPRB48wIDyBHCsbuy753CJQZDjqlPPU6ch
7VaJ9aEcwUkbfIfpnaFZFGQqRkjvpJvNc+HbZX0mvshunRhR+Tdygc3MUMri8kSbZ4KhK0E09Tk6
cI2okhSAbFjIwPowDpgRTYKyvhdsgmDg7vRCzRRIB5SHj1/Mc7DjG7G3JWlt0opaSeEhPEeJ1Oew
uvBoCfO9hMH+uL6CDC5piZcyHCFcHXYodVJOtWIii1LCZ+xqBijcQUW8EQmXV1A/uWgFkhKgQSA/
Irrn66rDGVvKDSAWhj/3TftVSDbnL77xYJKzh9gOJ3KNevu/SaV7n/2wLidn6ebQp3P7gO0dtR8I
WvjOobMZ9hvLWVmmMgEgfC98i+7141clDLORZYxTCa+xI/pMIXhlXWXhDLBc+3s90ChAO6lPmW2d
dVW+XVKQXNJRgAr9mATiMZkNZMjlMHpkk4GU4FDRZx+onzLO5lyeKfoo30CVlJjDIGhH4Z6nIQuW
cBquqq/MnIf4skkyHfxdCSEUWsfXeMSzQYu+wtv1P2cqtdD1dbsxuq3TfMK8ZvYxV5UUN+/ZwqRz
2LrYcSwtFxLaEILWP/nrtFT2UkcLd2U2g8mIpLbjxKWlPKH4Fo652xx/SqxM34U5AvCbpbLG7+yD
AdqzRmP/wXcNq5V31CdEakYDrpSUTttdJ3/iiHvgBh7ga0xrmsCHKbo7yTQtW8qrgi+dm9k5TBjJ
iKYorMM5c80VYtJmwDfjTvVx0epwCRYzuy7gq+g+2Msy9PLYTjrwQg6MIHB33HMtGCyp08Cscs71
i1K8j8xQV+ynedsh3YyekHYxMYN7zlaofJnugz4mNS/mto3rY9zQOJT9WSjGsVakVgJsE3OBIOTR
g5Ort59+A85F5WVDkUieenMvbDZT9vpMh34OuhB/5+aqKyRDd5q4UK6dZ0kZ+rT5HW/9HLstKCp0
OxKpLi74s0kvfEt/0O/OiCy5H03EpBYLrY7h//uBH7b7LsjNhM5b5I+SJTfJi+tFs90N+36QzSoS
od48OCE+DfdY+Kk/BIXm1Nz0Mae1UltSTk7+ZGswbB5Wyi84ulO37LPvaD8a+7a2qD1SfQi/3Eky
ZGweSgXJKIt3uTteSqgQOsmzRvQvJ2EWJcg5amocwXjR1ckRouZFMG7sU4kD4xNXnNT36dQykOFP
FF2Wsm037Vyugp6fpNvFTDWUyiVbNeNv5mirXDFtpTARinxt6xhzJ5+4KTYUjzsRRio9MhuQMT9s
9beLRpeLA1bFudcaZBYoI/P4HhUNy9QXLRxxUn89YLPJwWxERpi0x1rYo/aJZeyq1a+Eg48IUCwg
uYioCXtlja2w2S6yOsxja+ZTWyOe1O/2Yx4u9oBpri8NuwKWctuNETRdCan2egaDZN3Ji4K8t8s2
0ZnUJxvH0jnu0I1QnUhj6NBwx9nSrKrIXsb7K/pixU7UkA4blXJe1F7GaPhoK4Xt9y4mmRqV7X+m
c7ZLRmoQB+CO3M7T0dy5KjF9nSHprmGFgEnQG9JzJfmG7Z7p76EdhCIo5uV2H9twy+1eBVlz80Ib
A8ozA/MG4wzLuUny9s+t5Q7VunBRUUPHEYkPjYiaKo9nJcKLtS9OS9u+X0JrbTwLo7D9kiJIey3a
eFeHR9FQqJY+sU+rVye4aZCsXjwjoRF9A4BLorwhwHwu++NMJ2/hF2/py328cD6mqBVwcSdwry2L
sxsoLerGcPTCd+K9uVqaeJ25VrM72PGxfXZsFQXdoPM+cH26KBirKKG7pKBSxMmzy3vZ8XWiw7Cl
pFbCHz2xM/d0tGBrYtf2nVpF8lsTRxA+9BZStg4Hsj0B660qOVrVmyu5M3MqnsHi7UMPA6bPA48z
S6cZ55EtN76HjfTJWRpN0vGzt+wV0yVyfX11ijl6b/j9oAXNo3bYLBLIbPz99Tb0QWdGT7JeYPXD
igxbBhF6M18736RH70U732RWkeJ6DDvXpPOgegP9a/iOHg/FrBc71EhKkLsv1u43pRB3Y45Dezbg
NyF3o4UD2MUSgz/a8j4PIPbENCkhZgNebXEoiHkVkSkM4rHVyDYdxx2Iwsw5pKFT1XjwX2BOZAYb
DA9RoprxDFydRMV9TbGVvmX9i3/nlcWdt7G4UE4tKVDMcSZ4ZqLInEMAVLW8ZMeVv+vAad+1ZEZN
qD/36v+Vcoe9ZmqYFKFWqOrX1am7IOSvP1TZbFjsxzuW0J2VTgYRj74FDvxOTBaMfCySPai8UH8C
FBVHsKdZ3KTgFwzjabkttbdGhnf+Hp1/wPpaLGPRyJUdJl7qG/ZFoNI4nsaDm2XCelz7UeihNMRB
l6DHG6eRvh+MKKTBwWEMVyS6zEkr546dpvOuRVPmjeDC4ZeWPCKtNq1CgnGKhW+MffILsDmh8MTB
m5eyQm9Yoaoxb627XdmnjriPSzFwfK2DIQDXLeXLYxPQvAsoiQ1qdkJqdSeLVTk6YxRAjVrsov9k
VP5stbOjTUfLkoPXEgvqimvz3TLvR6t+FmN42UFTrNLB0yr4bxTW+TaZrO1DjMldxOm/3kiIxM1i
yD3UOyxxJNMAdbFt0XnDjFnwT9JbelVN5jrNAJXYTxekaJbj2apNRkUwMO0WM8BgL7M3bOZS7eF9
shSjBPhtD0ysVpJmo2G8TrJ6HoNviepJYdciCe+58ZXeSZVLn8bgSLuW2EVCpcwJ+CGW0AGjxbQU
oBATDIEvHVscpe8+3bvA2A1hlK11AZDuaSWtGTrV+b95vyePWU7IEr168+XYDfO+k6+NT7nyioiV
Yby7aFMw50xeJxogSErnNZ4w4aI4VPlPulIVk4FLtMMM4adpw/+eDO/P4V/tRskrF79y2XBU86bi
dH7uvEXx6ktMjcj0VHU4RySm8QEM8eJGMVgi8V7/7rBLqVziGt/tFDdUFZFBqDTDnd/kcRROrVqZ
flZmdtMR9U1zHAAw4ngo9CULDqFTrNCaxCJha28NjcyGrqIbS/QXrMhXUqAwZdql1RdwUoUmcZX8
6HTrg9QM9v53Ay4uaNnLKd73HWJRIG1ny8zr2LFQ1VNv+XgBIRseu9SzR6/Yh8oC2Kx0Oyynz0v3
qBOdvsMe3GgB82wLvqbqQeuWj+MoGbfPjZPU9Ymcu9TMkrfJPK5bPS7g7SOewPzjc6oPl33bTC0T
iPRUUj5MelI9aLc0ulkaJjKzqSMBO1tK2iYHIlejMTjYAmgGzYpJx6Auf10Oxo/JEzAHvQf4BRRB
U+LB00RfXfP+imdEVLq7d2wiGVXxvyHKtlRsyOUAlTR76lDjvk+f8tsEXXzw7FvbFtSWJOiIAali
5ztM49xdJKJztG1xaKR2XoGYYvXVbEPLQsOdcc5H/oO/+QtmIyaPpj2GRv+D8vkpUKbXG1yzWy+t
JFdBIQxYIseIu+xw7pqIYVG29llPXeiogHA5No0yJhY1roc5sv3uet508oiZxjGzjW+tkVjulqIB
BhNTYShqoSLhVv8x2SAdhScmDvZn1aKzgyLo6JupYaZRR3slzjLjCgk2RYUdSPcK6JCiwRcthEf7
/c+EhZRgHrT0HKBt+EqRfNI0twahrt1ke2sXZF1v5eG/rJP0En7g8RWdYxa4DpWa73feraKCVxgU
GtZdmVQqSxA2OPs2DlPPx5BGmSOxHEubuDtL3g6LV7tDtsmd7cPkh3BUecbpjUowJlBf1KiwnLZZ
mr0DjONFshgmLtkvQnInLtxB+ZdxQ1ThRf0loxJgKq4nOFyqhGnWbdrbdtWAXvYK2NaaEzmyrbVl
UQFJ2qo7nHQabwNiZBzV9zRI+MJJfbLFYNXdpEVKmsyH5bThRArZ8ZDDCiN/M2GKVw3gKP30gOGT
6yn01HJfJXQ1rc1wsLQQbszYvZxTFoD/KQvVJ6KsGZjKFA1LqOisKNA+JPbb0d8F7YzQdlP0zP6U
afqcFWTSKi3/XAxrc/p/US1MsfnBponrZBeX5TjlzN73ndTJWzsVTdrxJQ8GkwndEP9Xmj0OwVbw
rkpdnhb8cX/TDNzvQkYfOKfTuTsO0NFz6j0jFhibxvkCBRqGnWXOkNkdmnbcymxGKDZnN+1q6cXz
s19X49Ee8fBY3lnVQbxi9t7NDivHD8fDP7Tifl7lPLfX2H54mfTE8zK2TO4ZiRW4/osuRZDj4UZc
UpfJPIcj24p0CIx7YTIQVCKlynDlk52fgsRaz5kFVcLcVJBD6Juk70IuFFNTNf6HnR/zdGI+55s1
JCD+smQbnFeJd2hc4GJYc02qCnQf1eIkONZnbv10Fx8E+YrnLfggaYIkcvljgRqnPGJQUHp2ocjT
TCY+58dviVgrFqd9oj+hgmBVvj76cDnN1AfOswzkwSu1xICvkHZPUondXnZyNUz5I77y2gwO1Xop
Gy6ZXVKnpkaBYOsXVzzt8eSVzvJOdgRoV1XgVKb+QDiLlr5Ex1qEI6URREGhA2nSYR+d4akB3EXy
tlKGX7FnC1R0+kYZt/INncy5nl7keECGguCcfv6VButYqDzeXtpjSPdlw1fvKyg++r3n4p4Kq9sq
DrYsocn7Uxd2bfhQHfwvh2M7JHegX5JztLjWzq/zdxtMncofYaNSQfdmG2vsnsN+UEJnHQjuvSfA
tFdZdBo8DR5oMf7Kr/X7pa0uGPQLTLrt+wnwPAivelqOWgg/jl2oniYfYc8+EWTFhC0aSl8ByTwJ
Vw6GgZmPV/NxDI5zO0ipDky7zvUYGKLoYTRpPzKed58tBNu6qgqUfPRmEtEq/SZS+BiTXZaaPch6
PhWQMgRviVZiKU4tgo8g/3kolQ3tSCzyUJRBdhY0IuOn25mRF1Rlq0U5NuULIfPQhnjteZ2o6y0K
16e+n9JM7mrJAwQKUIbbmKN5RmwT0tMksUTXhJ5Uugc0rgjGC36PfgNUzyZf0vNaNsQcdwnnHAY1
QwOhIPTsALovLvuyRZQ6iIOMIWF09ALBPq+lXMs5gO9195JrKk2KDl51UQTEQfvandwskeATM06Q
ugtwNRhmWF6pG9NlMhk5TUGhZdEYgJLoe37fy5tBK6vMcbusIaNyrKeDLjb0X3LFnpVD7MSDixKw
Sjzo/9z6Z4p9eio4Cq3UmtqIYM7445yhafcHM7NXJVtRxAD5tPN0P6NzWtwjUJdelk72RCUIuuNi
VxjIMRsFmuwFIyspXeiPaHAqwtMVlGRqyBmuNIffbKjWC4lH0tIbJ6qePFEArLl+v/SIEnONrqYb
2mKyvREhPnWaJmjy/yGiMYIwI+23H7t9d15a3EJ6cJ5ut762+0RTCJ4WtMhLCeTgjV1H7ZaMNlOi
SSjis99/YZj4Z+63apUUaa9NlqqYP1YxgwWet5WAsfeoPL5st652zJlthn+Xo1jEekZwyd4ArBsT
OvExxOLqirCxqdB18KanKC7CJBA2w2NobSzKeTQc0y+rLry3Ytakg0awoPGTEZ84lRUXZRtHGeS/
X1TWTlSVMGIo8QdCt5IbnTMCFS6uIGwzYU8ezmos7WyN3DurnEu0omxjAG7mCrPJEkdDp55GzL9x
JpUzOMnqKazZAhDgQ3hpLPh7wIDMlZu1y1nKddacp0mGZNhGIsiac/tBIAzvPrN7LUJ4i3lImp9N
avcSRgpsqi1QLWFuPg8NFvf+PEIQq9OPzgK/y1gbAIKnAKIS+uHMPjEP8DoEn8pydcfa3i7BwlZz
p8e8WkzHYLxUdIj0zn9hmFBmnM9JZu2nLsSG6czeDEElgga4022GQEXzJuibuf5NGbFvzjw6V0ZL
UTiGM6w4R+EoI8NYXNX9Fycv1diNfZM++33HyJ/a2o+9RyHysdb6WTpDSfRRYr/NNHLcWV620fVF
pZ5z84Rfgo5UMD0DWz/GiqHmTGOr2TLf49n6E1N1tA+oNlTCxoxxTdk7H5uHyRH4Fx/MKN93yc5G
KCToxBqQ13BjVa6yphd5gavrqO3VqXMSCaDNxqtURLh4gsfMTdXKJ+Tm/1HWWx4Lbu68sGvIjv7j
F3Z+Jo9w/DjDfsW1T5ewFnsn4g+Row4wMna1RZE0yjAXCnWAp92kZD3zTKvUlGSCQvCOILf4NQD8
1wI3IiTN5+VcynZf21EgDBwF3g4eK0Cj2PIteUymItwZl8tKH++SNLn0Pgrr9VbDs4OHWelDkndq
+yQqdKehEcheHysdgIYmUMjXsa/78TG1VqVNIkU+SofHoT0qInCKiScw5bIYugwsGEdli2Egbmz6
5fWWqVbkFW1kyXj5eY9jAIEXm9VAc8xpNOZu2CuyHIbIhEen/ls3wyu04fuQDs6V+WttKqhiZn/D
saUJ71VOU969A72PJlM5yABDAXKYKq5GTCuqXcf0CnlUpoIH2RNRFAVAXTg2lq5dH2K7GvMMeuJU
NZlrKi+OSuMTF3WDAMW8AfDoXo+Wd80ShK7RFGreUBKvodb78C0euDXAsn+/pON7Hqt6mnIG85D4
ScP9FX2is9LNRpKy6lYqrvGLrmWGDQayPRHx5rUTP3MgQJxkSIdjs3ytWKzr04/vegFbF0d3LH9t
HGrmaz7Y9mBQgObJjwaFEFXxP0sPI/Ll7FJBva2hzQqpdA5Eh8rzC5lTvmMtSBRj96bfXBLr/SlC
saLLgXC6es1E7tPRUCvGZJqL8ECyhxTOfpcK7ayRUNxBrmZwCkHrDB9SgjeI2us1r53zy+GrZUAC
5RjWeWrCzau91Z9RjcUanUFkPkK+g6/JW6uE/0e5YTxD0DbIb6DLtZgHR5y8IJqrBNbO4NCvg7uN
OtyMXwFt7BIrLzpnEYzsa4oeKa7mVnNCUnmv423kmD9+aSLpIiDP4NXxYTsueUqTk8gNCVFi4Ycb
XZvmVk/MtktoFW+yOoTJOP0x95jy11fAK4gWLkuRcSvjJ0gPS8mgmg3oy6l9gJolGkrfte1e242s
cJ9G1E7c6xisaHkp5ZpVhilyQM4KD3qSJnY5wwfHmxrY/wxBxB+oIOn/lTaEOqXWF29pzMojYR8V
+FG567EkegV5Xh/ejwVVGkWoVNQUgNhht+UM7vFsSFL5t827LQgnSA8DROJR63Wpr8sFn5R8rwom
eHUi7A6OBSulPZMnvkdla2v2XZ+UkETbIgPovJ6fEN8mJLynvxRMTwQhbcl0UiM0Al1ZcdLS7+on
JlNaW3A95lMwxFMpRIaMyJ3Z3nSKf2mS/7Jq56ohxjghpIDx2nUjJtIsen0eADxPPk/5zRAWAHzh
QBzVWtVpOdE5QQZow2CWjxe2AOlRF35w0uzifi2ebvMKDG/Khr5TfNqC3MyhEcuI0CiNSI32p8Za
vuK5McxQS+AntDfa7SON3aZILmRgHotNl4CSbyD5Xwzbmw1j9xCWnje8GKq968FJfty03NWsZAc8
4C0wNcyc+Bkrctg3OOrxnwDyVFDGpW7XodNSvS9C9O8821SJaPCvczmm2MrsufkYHhOnVUruTOBm
PgyAcp3kkp3YQgNNXzv/Tf0w+/ol49aSRv+LBb9satqZOaWGIINH+xhcuz0KBtyPML1iFQ66y1+a
AWjWceNFpNRzi23wEN0snLI0pJYb6RvvyWn8BDtWfzdAKcAuG31VyFDQQit19NFbjkXWG1EF3Bz+
lW218vqb1lf6p6BVD9kIRXMkheNr1RFdvRqIK7kEFcclYZo37grTGUT9XViDFMlnLRkGWwqbIUtf
kxOUMmYniijTtN3j/EIf16c+SAzmmqwHFlj70cVrj/URjvKb5Ss4Ayx2hYQPfvz5OLHYac+BoSdh
eeGtqLI428f5Gztvbi6HFTyMM0n7BVbjkR5fEK5yKnkqhtS/PvnjCYtRLvBkeNwgq++KtHW2oWCA
LcE9z5eVoKxqPRSLqMzxZc04IPr4egLh4vCS4LDUWU/6u99RGIl31hqjx/9Pov0wtHN6blI3Q3hD
pbwd6b/MjPyblanKEr5gYLzt5MjsWkM2IowGKVcndIX/7gD2ztTBRy0kCMOo2xqediXYwCxjTP3I
Qxu4BqLToTqprlcL7vh6Bm/u2SdZG3CuymSP8tWufIuGj9PJSx3RxcwHEU+qRmdRAHwA6bM20TWZ
WQSDClbZrAWwDC5QEmsOZG/a+PG8wRflfHwCyP3XYhMbffx+e+0rvVN+wr91NuXWpsThdHPG3YEd
T7cXiY3jRegAgoHE2ZLURzbTPvAQvYeuyrUOH3NrBBjI98Rgb6PVaxwwsH9cz5J58yKGW1/vieTJ
UvvAFfF7jpUNwL87bzwyCJgEMDkDf765ZJxu+AhmrLcJ4ekXPzQAoXU4atTzngkupe1WKiurmp6d
a6Rx57ZruJYXOZ33Inypx1/cfb0yUeOE8I6+ZvA6RRtOE1ytuNWLBpKXztqkhPSI/wtjyHhmETUi
BtiLTJkuzCbND/bvUA0XXh/b8QmFHTJTQJ05kqMduedqFyc8U02Vu4Oe6JzAWQMzGdZBB4SCH/ah
0KPmkK2HsLPf4jRUEAecwzFXv2OyeUVlL8Yu4mMWqMZsnJ4jw19wPJamVxlja+7JneqVb75M+0kX
TKigbHcVSuYdESh0auyh2k9sIilmHhYOv6xMPG79GYaYJp+9JtNCkUEZmj/DIE7eDyhGGW1aLtU4
42dWniLNiEjDg89nAN2E+CcykcBKnGJ+iBJWkqT8D+toqbwL+LyCVxewviVwFrqxWNZ7Gtu26kTH
rFHPwoctU+zUKpQx0gj7jNqux5f7gNoatcz+F1Y2X86BFCcXib/y2aihKExkiVbs3Ejd0cxIdyD/
hC22V8IpCoTsrgbFjSdHyHgyoAjQADetlNGQcyX4p3tSUvJmqJnIoFK6OKI9CkIyMPa4fH/jKQk5
vsB1Seun6k8LJvsyNdBy+SG4ue2m4myIEtME1kGAB2i+JlAma9K+Rv6Z+hOoxiKP60Dcv0Yod1lQ
GIkzGPpkMxKSG7YunBetTcvVVy48Vn2a7Ssj5/0kIYuwSbU31bnhV0hKFXcpjclQ1JP36X3xt+E+
BWcM4BWjXeFTbaFzU1NTZUf3oLhqjr32YAo/0Vhe1KWOIXUM0nKXjiNKBprjdvUD3RKnKkTvfykQ
rJq6vf/sFtWLHpTU1ksfMocW7KeEI4Nrf5CCuV9mE4mk1DmtV0T8elMuUrkwcHQtE4mbwzRsUnEM
HpI77S7PpiqryBmYmNMGfmUSEArp18jAWu4pV+Lk2Pa6lWwXijqewB6oO4SoLs1LHejwe5Ni9jiM
f6Q7MIqaXBmyUsdHBAKqQexIyePYZdSAT4YjiU+y+9qOJOkKBIaanq4tPAgzRIcM+i26o3QJvMHX
l28WfHj6Zx1k6iXEEDR8KIWemuIRavJHbhBuJV4wLSC1u7aLn0WFddVBndqsCsnoy+8kO88gxvWy
RCoYlHYLDSIiARRkq3J4GwjxrQrzk4yoK4ZlYEaVr/Ilay3lOK5xMqx6NK9lWLJETbiJe2tsBVxi
7swpM/S+l3gY9397gqQV2TTmvo1XDV8iev7XzoIsdio9pL3QEOJOm1Qy17/IG23k2+/WvP/QT/cX
ZX6IrOEXk18MnnOkapbmLt2tfLeESSh21Kc2FNKX4zCHwp2T3daGUHdfYEz2suNd4L98j0IDIbku
UR5/iBlDNTDdMWj4lnbVGfKOatwj8BQshBYrGBjYQw+h/5tqHWC6bVZvbV4+m7V4YECXEcrS4F80
KBCE+ZykjxwzdMZ1RtkPkq3xeGw8F+TJSgg18Y+89cVdP7SBsy7MR/8FtVFhoz5nyWKZQQiapZmJ
TQFb4Ut/0hsheNyvLoKt6vEyrg4gHIlsgaG/qHDACQe19kgrVgWeJ+bxhKw+M827ACBjqwvdVylU
xPCFaaxbLMA0yia01BQEan0HB9ysgMO8WXSxJVuSHsCBdPOjIDTaHsoKRhgqZUSslat6Qtw8y3r4
EOb+xFWsvReXBSSreWxzaHUPZNzJDkKoaEA7ORzBkoofa82+WRePY/cZRufy/MKefcNlpMi8KnrN
3pl/b6PmmjzQxYW9pFCMTr0vbOh1bf+ikSXDOmA8K+dxVJ5xdyNkTuNQWQbn3vTCL2j8MRysbwd5
I6DKLQuoPcMpXucf5v7VEKGxUKLHVN0mqwUW9OhEGAiqca8r4LRp6vz8dxuUCEqoaw8Y36bVxDb2
3Of0zUiZ3dpzrQNvaaAZ4SvgjiN1uVWSwAS7CbXy1AI0ZVbQ5IVki15duob4boOdlMqvl6haflln
PIqlrQ8HU9UBLIy2qxP8fePRyv8AqyX3pc60mKkxZhgklaXOeT9uMU5zF9tNvy+2jRtznV8y2nZz
He3ZdIBvTbqlnckmcb1qLYfWNWR5jcOUH6Vys5zmxtHRhlgA3r24GiTg27WSZguqwScEw32sGMtU
UnSdLQyGc1Un4jUoHPrZancx6TZFnHW4UGdciOumMn42pHupyLkRpjOHBFhBWvt38UfARCyXsWq0
rptxCND76xr4wDiTvf1qozMZUOzobnaAUiMw7/vvk3pqI2n4nwsKyFsH3l/bflfVL1juqfuVSiXI
12VeHLQyOki1bdMfs1PzUbzny4BKMWzkOcaN/mbcjN35HLD9aMU1ZwdGYZCF8axkBq1RbudVwCSE
aRDLPVVS4/RebY2OyQZkJ363CkZW46/sy6cZxTlGTzlLmJ9KgW2IzU3SjBS/uh+4uD2C0zICsRgG
7IaatNxavQilKYGymo+5DXyuwirw5hhuUrLPe2HYh/+uYp5VdU99/jcyJgqxGM7bqDrbiIV62p+5
/UcAos9KwScKDAt+km68hEo4ruwCWDsct2YYvqWkMGQW758hc8jNT/WRuBI7KiAFgaTfMsMq6ONd
7fNIkOUItNkjuilqkhTcJtK9Nv4eIAv4aA2V0Hnzao7wg390gel26RltHw8vVAk17zzqZZ3NxJjl
Puvo1MUMkVk4J0v4ORwT0qRn7ajlbtH5WuYsXESgdHIA9asniRSL+RxB54CPTNl11a6foIKgxzt4
4YRVV4UEmJCMAHGLxN7VYdu+UwqxZ5FZ/I28HJcTuUyNNiRUOKQStmOGvZX7KZuWuZeS0eubTLJ+
VK5LuZ1rTVvK4lLItXcao8+iLk5eyag9iMeMVGtW+GcPl8stLRlK1dVOTmwwg4LAv49ec8SOcLNS
QgNINsXQtCopLJRZttrvpyYJ+f2ATbeG/224K0vCY8s+BX96Sd8DBPF7MCG6KwzxQOaWvH7kcAhI
Y/r57N4mVpEfm5MakIxeaq4L5iQ7Md5kFfXYAuaGZiPOJR/Sgt1wbDgMNSFQr8kkpXq3V6GEb518
2bgSd3VvwCNZ5gSGR8JiiyN7mupxUNwkXMNlq/MRsIfQPgtir0ArZfxrki0JbupFcJYXygJnLMCD
/y+dsRQ6kWZxgAu976gSJ0lhrR+p5w9IQiBFPMsKlCAMc2ztSiRewb95vswxKtFhWYhfuzW3beUt
CRJ9VRBZeK04uckIkIkoRZNwIZ8cytPo1+3iszfCcbIdbBisEPX52Q+MNvgjQJKMV7JBXZwtdug/
LYNNBfD8QOXovo7k+I7zEhzm8a3xRXFZIT6kmYeN4HNKLcC/s+cCdVPL7aA3Qp7MwIt/fLJK1FcW
ooIa0H5Kbls7jhFBOCBxAt5nHK4v/5lFOy9cqeQH/0MzcxUTkDH54D9aY0VOYtVKQ9RnYCe5S3s6
gvxTaZMWA/X/aOcPCdIa0i2fnAY4mM4Y/XYF94vn5SYJ4Q9ignD5zbUqaDmiGI3/ogR4QesESvpt
GfUHl5ocOUtOpBK/snhjjmZwEh5ZyxMzcLsMOqvU5sHUqgLBqttJIXA2gidOFIQdDhT60PKCw/c8
EfRTPZkentGdMW5bPbeKkV8XRoWLbpEe6iLondUctSx67jk8kHrbN5atRvj7Hg+hI4zL3ZFPRCxQ
lgWQ6q0K7z8l1/qJszVlgvsWfAhS/DW7wh5JupyiT9nbX8mTa/vGYC99Foqkop/8Aly8vshPIrzo
Om1k5ZQSeC24UYR47vhsrHTI2P0QXw1xydypa4na8xGqeENke8CygRYyeD3PFdoJpoYotEN2bQyt
v7l/2w7Ky6eSPQFMReTMElUe9a5sMyuGltUMfTBYuHkcvJMtKJov0bm28QOqMphHz2j7HdRES0/f
sTJCByjmZrNBC91yTozBStSU+pPS2uLfiVEnfMBUS5FyAt9MDAOCol/t9APPZiiajvTuCFFBprmn
S4TIe6EdWefzEWhktEOtoMYsZZ0kHeFL02FCyB2x/CB0rcw39uc4SHxp311AZhJBVxh3J7f0w4Xm
c9XHAK19VuU3/e+Q5kUGRhInmOVw2ADMgQSEMnXKIJdJsLGiu5TgfRifZjw0HjTlpLtaI+c2CuF+
gI+GVENwaH4tylE1JuiutRArOLZcm+PuVmCwJOR5ZLNkQREZpJJKE/PTsQoeeEfrBZGp0is9+eiP
di1qfeNOvJYWkPXvnhVSsZ5QKY9Me2N9QAp+1bG/NsPNgDfzowwLj7+u90AJS3j23YL/xbGH/MNp
x7DF+FTt5XjZB9izYroL0+gb+RgcAnCLK47cgEhwpDKTg4CqC70K4+AqaLHhXxzVH/bvOrq67+HX
TuJMGzvNkG85rh0pT51HszF1drog50W7lN0sBn8rNDj4EJ7sp0elkmdExejmGPm5qJ4eim0+O5tG
8k0K5GB49OBQsWQlp4NFTuHb6q59E5836cIwMXEs29t4G4YFkkqIsMn/MrlEgEUm2fb0sHPRRfTY
i5ICUoOZjtV6Np3gHxyyZmTuiDNDgvXk5BaeLU+Tjsvsyz9OT7qKPho5+pImX6URnb0bE6z7KDRT
irYMegFsEoq1m8jnHu/haz2bp6kRllmlcxp2KKt4RNyaqA8TQiVp8TmUXtAwppFQcQH7ZGGoxgmg
ebLDUH3Fl8btZANi4jFy4UmAzt/3btJ/IvBaHxOLEX8K+cZwCQWqzvJzwd6kJVcrsPxNuan83qpF
h50orC5l8EGizlw0w1lI3XhVlEOQeRIQOTErXdck30vBiKLaHZlSvaCG7W3q1B1K023v8BaFS74Y
LAzmzArUj+5bnSo7dPB8Sg5zFQYw7ZhD3TBfpGvrDM6Bp2B8kVMdcnsXv4WzPpsD5k0h58cnlIGS
sNA93f0LrXkL90Jk+SrU0bi1HFy5WUSYg6oL0KVE8W4qGvgHT32LSxBMrxmNhtiRalXFU8veuuj3
LhILdgYDQimJ12Bq8rGpPHIqvGzk0SdCboMrHBssdWqHDynloFt7l+TchtfJrSDcA6x84j4WVPaG
taW+5JGCNA1U/idvzXE9tqlAfGzpYnSSjlKMA1De3dXNjYbO0kCKHPr7oLygFkad9nnQSIsZCB2c
9+rqYfvVSneXZ4TDOQvqQnBYaWGXf5mejlIIwgmmipx94h7RFkR+TXfFt7PJ11CydkoU0y19QinV
gbO1gI1qlo6fxFdXa9/diZKKB4Q4C+CsBL4fjn28AIyzRsMPupAgpR3fyTqFGd7o59+eN4Jy6DrV
I4JMPtGG124+w4qO+qdDZLvWCQONKnzDRNq+nTG8vv3/8f92QFZ2mKqgMQLwx2sT8/ic22ewu+4W
Kfu340CB0gV6P+nEYV4KM/aIg9cOmszzV4p557N1sPqP6NVPiibXbj2PPhGHndfXkxbU4YleiqKx
ORmnQLXD+S5RVPsW+w0tnPxGLgUcFVPbxFmQZtij0IIHFT8UHB2ceQqBT6+fPZw31eOTq2pCSWGQ
yAF0TnEPtQV1uueJ93W9gxmQ7GC8yoboYbBPS1H3NAKle6MFsHkpF2p7trRzjzrIUh6Pc5jxTSGL
7Jj7L+5JN72i2qPPeUqr+eW6VUaZGweKITW186EQsT1Q3L9aqC30WeOlMTlriZraLaHNRryliWb9
aK3CIQ/8htfzZejJQipXNq0KSFYrgSvqQ/6Q3pRsudyDGPrnB36+R0QtRxQsSK6l1tYxiaH/jwzj
/8pQ+lmy+TgOW5veJx0HOsaKUy0r8RE8fhU2Lvbscg4Om/X7sxBG622taNo8eOdS+Q0OYCheTxfG
ZQV43j97mJznXjBoSeVKSRRHCJ7kRDDpI+ufaW5AEgD5SyS+YPjOq0BzaMj+jMBIGyNQWJ5ZieK/
ler3Jmhs7gyc/M3QJxrK22JeLS/CqlNjlpfHxvLHJVqbtsOadztE5N/oqAPuoo5tnE2F/06Ttsug
aRHqAT/QGC2U9BU+MUtKv6S2pIfJX34ytKWBWFAzkgWubwCR4IFFlFjNpWhmDcT0gSqzUs1ESryZ
y7gxEDNm1Sfo81OtBjcArnAN84nuMPF5GmCCojpR+cu9GU1ylBZy1mBl94tcW5J1Fr++HXXpDOqG
d/HxGven0635TQFb9GWwsN3KeshM/wo9wX7lrqsb7KZz0IWPa2sBA+jbG24X2hagUdRQi4nUdeXp
HRX+aGrN8rJKd0Ccv8kkSAFCLL/muDXfXu7uQuzyGQLN37w8GSvPCkrslxjUUtEU68jqs9ro1I3z
QtCerbm+9GHw3st4sH5BWGWn2LpZXPAb62sQJkurSUn2gT9HIDtELc7xMD7xeDHde6JyEjFoduHb
syUbGS5+evZWISEmwXJcW9MD7GB/oz4xtqBwgUjtJ5gevAjackA66HM6yrHnVdOyl0lzphVxj/7H
O5EI6L3JjCeIMfH2lI4V7vqK4Mp2cU57CsqmoANttAJT2OZD1zjqgWrkOvc9SLdKooKbWPFsWxRd
6pAaOEx5VTIgvc4I5zCdePH2IYQxt1zF/ZqQJeCAatiXHxeduVDSkd5NDLOZZHqEwcMvhrZCqfKM
Iq2YeFLk1q96/EM7sfkQePIStra/vLheFrVrDwXWX7CBY4b0o+LKsF/MK5UwaJLx2ywJvN35sEZo
xqSn4foJQknVYOI/sQ+8fQkALtMCXlwEgcVxOo68O3FiCbaLAFG8RWz6jdxp4AFFb12nypdREqvT
yoJBPcIlXd//qcV+GEJYdpd5QkmtPyIYnFc828ergLxKHZiCmgxc1zCpWZ07Ped7C/VJbCerSVCp
5JYQjuLHsPFXJrqZncMX1UFr7qwZoxpp0MAmy8mVdJKF9xIX+m6Z4hIlOeWLcTC41vPBcJr7XFa1
86Y3NPnl7jjwo6rYSMgv0rypXFGrYGSEzvn2Y7PBJzNiMdWV4EgE/biCme37Fzv+nN2UmNsL59ls
LMmGXp2tIxqSxIb3x7q11Ro6/FsqTEuHSCOXCrFeZWzEWjdtvlHMkrLIpcW4mevrHDtalEPsyXNl
DKK7huIdDS4WEW0N/ZavVB0g6x/DDdZfivA0OH5oJG91D4xS3xUzaae2ezu8Z6mD2GDN62DWMW7w
xrNFR7lnJSLnpb9r778m4xhxuv+4MpyOKHVHJKawxLEnybsDxfaOh6sY2QYs+623CpDHo8mGrW8i
UHeCQeU8SIsxPS1ZEFJOvsNkGHaIzyGE+IBhHFKlp2Sq6H3KVcUj/zAfDy+xkGW/S/f+FfaZRJIt
JugOG/HZ8ZI4G+8PcaU4MlOZkGU88F5Zi+s2YKLE0lD7GLGqaph8K+SLm7e+y5LWQomgoBaJ4JVP
1CpkJo4MvwGEpjc62yhkUmHQJ3xtv6KR8OIrtkNbPIe3EbiwfOdc62TnYf2s3vdeWWkQoLoPT+d8
Ju0/QvuX1d9YLZlf1F8dFC7pQEqTM752zTlpy4keaQfbGcaOcJ7IYc1tSwv9X6LkuScPkzlves7a
QybuaTCPLShCzp7dvT3T4Z+xTXJh0MXfGBMzxaqVBisn4HAhdxJKPBzcxR2JVO7a/ZBSTR36lgoe
D4Q3OQ4rQageI1BPyrB/99C74JqjplYzZSnE8AIsmMGUl05pppUkSNK8CvNS80vDwPCDXmK1I5Pe
f0bMZmPA1DEvIsT3o+OOxawsxI4nJnnRP8FBhlwjtQAwOZh6qV0pUs0znKspu7RpyxSFvN8bjJ1Q
YS4AZfu2mtsXbNm1V+oNP8m/Baa5ir7B+XnhRJ2xECUMp4UWzo0sJeq7sg3Lh7ocIGp5s16AeZOf
VlOPNay1i0P4I98CqrrUNqDl7yN8abHfc9GISvROK2qTQg9RB7nNVTM0RkmXo7YdaOZyJG86hl47
MxSu4gjy5v9KodQGMGNvqxiEyVrUEII20GFMWCC10xVsEeoVYHZSKBVjetOUPSW0I142ZDQj8Twd
j+UspnxI+cQaK/KEFp6YTOXewGBes4DjJuCLZL8WmNVfqHaJNvb92Utbp1oqss0jGgs+qjgkML0u
5oEWHLUCb3V2Bz+/7pTiq6ea4YynHthFdp/cZtFLFQs/RQb3W4Dfi080DTlH5Aya9+zs7LQY1oHY
M+e/lvuduti5lMZ+81kfLY8lRzMGVWsRWb/wqTfT2fUkDPfXR7TTmUpKmwXngWogBfmPUPNFphfj
KMCK0firJIK0Dl/IYy7n4pzcAbNlmJh6wu5irWs43ow9da675ozQ+V1bNHJar5Z4wg80ArmjBfJG
GtRrrrCv/ZwH9dnVBN5nIghY2kLMgg3GF0a2Jtv6J4O8+lB18l/QE3JIEMU1FjkaDD1pONLJLYZz
fyTBjTQSAf5UWcqr8R7tkmWJs2mIo8pxpe+UhHM9I9Bd794a9UCtVWope51G48HmEBMHDFTZuP4W
rpZiP0c4SePjyqBcT13A2flysilqnA6pwlLYtP3lPxSm+C58rcxWbH/Rxq/IdnSbqbXibGeBcbv4
l+hMI0iN+HBlR1+vAsAovrlZG6uhIRlMjSWRAFqfSIb5aVFlfmIDVga6/VDVjSRx0qn/4VJleBW4
O3mY7WY8d2KyvgoB72yTAmd0/Vay9t5FSqWstGUchZXQjtoOA2S3Yoc1h0baMjvgt2aqLL5TRBie
66WibYL0zsbguBFy7u2tsMmp31zfvtbzWuyuq4k2A4puKnbuR/k/YXb2T4kO3YLJapjRGo0rCkoi
+/VTMS9mUle9Qv1Ud6tSei0NfEXUgOjAU0S5XZ5IT+afKRCbgu1N1rsI7LdMQNvGkBCMlfaOJJA2
GJ2ueV/Z5W44fKiLexV3sKLWusxJiKoLWXirYXIT7QSHLKJZ9vpiwQKC7NhFRF2jtj9ZHqIBdQmf
UpHWndnubDITxK05iZpiK5oFeUncXXoHCNAnSqwmiYPGN6pwrmriStPMgvISrx3zX5cqXMuUEJUs
cJ/3PNDc6NHbg5oCwxomsTfGNQqCBs45upMZ7dzy5gn+G/pUuw0Pt8smgqvLz3+a7KjQrbo8Q0EJ
gn7alS13OuimEz9lqr8/uu+++rWOjKoUjr7/cTttOBdB4/wLEqqkD2yyLFy0PGSfA6Au4P1ED4jx
f2mmb5a5rsbzXuA0v+TEHsO8MH32mrBFrNyFUrl+KFCjz+hLV4jIFNaIR8DNb/COO1zXuKwScxB7
KLcJ6u2dENYKUWpi9wMxL7jUEW97/nUewysvnjOaaaQMD3oyDdgOzEkrp0h2+laPOPhGhCFLqpvK
Yiy3ur2WruepgaKlwtMp8iVop4/okwfCEP430/F6DZhihLi+zEfZLIZ2454QwrK653ZdR57Q5LVE
oQw9ESP6/+CcrjnifQ9Owp+HINDF3rpT/JjWp4jjEr71q/NPVcuCeREwm3ulaE7mZ15SYE/7kevF
9q11ZMqxKlnPgqlap7joOcZgfT1dFfvuNUBjxZ2EHgsFeTJ2W4pInH//Kom9HQJgsGlCRkKsdFei
bal4g+4F8F6ykGjR4N7Mqt774nH7tHPwwL5mPCB4bKH7MPwUHYSsrsFtPK/q1nYBEoErjtiiZ+N7
376PVShy0s5w5zzVTY0tEiIJ/7Q84UPK0z+OkPnFVBFqsvVuOluItDOb3Wp08l5PmLeFlDZafEGx
wO5D/5i86Ea8r4pE/AG3CEcAQB10pNxe3LUl5muRArkomlIHbmtkLt0CuETwJKk8sp3bKgkgQ612
Y4gshZjUhv/ZGRaldgOSsjcNDtIpuOoX0BSJ+pVXdKPUf+reY3883acKBO5/b+PxJc/wjzd+uxoq
fvI11QoBblDHLLeFxSZtVvvsNGTWCjPCPk7E5vKiBE/64QV6+4YZbXhr5N1/F3KonmJRTzl4M2nO
hZUQms+zt/h9E7YcJ5M7gpGNl0j7vwyC+81o/Bg5+C85GTXhbGTyFLtVEu/J5fdnlq0D0IECZooZ
LGGJlV3FCzmOZpyriChAuPCBrT0rW2PwEziPOLkUWOl7OKby9KGE0Xg52DjlOS8Ecbv8/eiRGbtu
YBspRd2qU1iA7WaBq+fcaYJtG05rsUIQGqqduDouCpFoA3r2OMoWJbORlkI9xSOCpt74dod6iDNM
vVtGtDWd0myVncg7hn4zWF+HgNoQELPbbS5Kwcn0azENYaKpA/xuqkfMkpyyxbtstEBGjYPx5uYY
gwxYC9+N3NPznbpmri6lYDWz6IAcXJCSs6TfE0+cePmA3uAqrLlQ1LjmHDcsz0dYGr8HtGPfsKAS
i5ibQfORvxpupP5VsAr6muSMQN8YQwR5UD8voa4FZ0dBDf7LOc85Af8af4Rl4dGtW4Cv5xV7+bvQ
uIoKTTP0OVYcfBvD2EBz/zppUrQHzoA2vGqN4ZqJl8z25S8+rwARKhQoc9r+DPGZ3AoSii2H3ebG
ywHZ40OvOs1X3t2XKlg88eHb4lw6vBkjHEgHAvZfBYMWTaqanDOld03yhzq+21I1XGaXNhfTJ3Zq
CmsyediZ/bVLeVR+NzBciDgY9ewzcVLtwEmLQL7iuLsHFrFOq2JjGvjphRlnB7OLASXOqCnCGvXA
fxVs/HF+vOu5mMTOmcaOdalUw4eoAvpPqwL+BhjLeBJwx5nwyUbotBsftCsXNTz8MFKg6cREYcWb
IibOx7YL9DDq73fkID7cYgCX4YPAAwEDlVSt5s4kd1HwyEzp8f80a1AD2hdd7GgeIx2YtEzyFlAZ
h7ME3mH+5KVn/z4IAkF9Me7BMFj5hQKcpXSXmmMSK+GGXJo6MFo1z/BqrzbDEFohaoaTKmefQrYL
YHdQFAmHhXrtX81Xcqx1w8E55W64RG+tOAN25MVkG12Jp3yMEeIGHn8jB6zruF7y/bZ9+nmV3FEz
ttuVaWh2uiDDE64ZRMgVtW8iEln6dbEQbapao/Bfr+WP81AajG07/xHE7lvSP/dvoHjXwSltZar5
LBQqwkWGjOurMqw9O7KoumBhIrfjw3yf0/fasg5iSSVFDVbn5MVuCDHw1zA1NCo4JRZRLJsLu0Dk
t76s4i4TunJGFoWw8SrpkdyfdK0vd03HaGAOrfZbOu575oNlCL371HSQBvD03eX6SgDu0fnIOp65
8ouFdsHFPbyFmHIgZpUYbjOS3jS8ofXap4v2gCa5L7fX66xBoM4KiR3+pejGZWJRjk2G2HfvX0At
CMsz8be9nP7FEyWTwStszAaFPIN7JaYCQFX1BhnVJeBc8Xye1+cnwUmF+eKppJHw1qns3HX0g5cT
GYmx3jZjaqns1Iu7L6zl8yaxciwrLp+GT6YQUs1NReFVqWgF3wuj/g/M3VM9Im2rt/wt3ccuTYQt
ACxMNdsSPXJH3WPxHUEzW396T0iyEDTwdQD7Z7UgzW2pPUbaIUEkvld3nzjqqzMldUg+AXAEWyQK
az7LduzHh8IGFm7XKkSkm6kwso7IxKGR1dPAqmNwmdn2TxZ053E9f0pieqiB1ZyX1dFhA31scTzs
tsQrOOs/wRMQZ9FwB64rrHgYs6YRhkrscv0+eFAWK7GwQ+wh7641FlaFWGpRASjuTrBujby6Wfaw
mYoydNlSaXya7V0OCPnvWKY+FJ9LwMLQrs2xJ2XLyztghlm4ouDBd+IfA/eOpCU+t6jPDDmW56LP
2C0iqHjFrZNuRehnavGIk+t8aBpfzw+/uTMLsqL7QqM4X2rLQIuNcS4HCTfpDANbnnNBFoh67+Af
RWcOqnkJ8EsckzfnuNQL0DB38iZBNPUDaYY7IwLNcV8//gP5VM/q0gZQxnbPpJJixbhoc2xCx6Aw
xNvaBFkKWkVAo+A/kHYhqmIQHcTb+kM5/HhHZYtKVHQOchS6R5fISMpVrR/fxmouKPatiGI32TdO
dSZOmCjphcAdeWcT9D33gX+6h0uH/8cWb3aN4RspOOkYEU3MoUr1dID9fITSm74dVPY5RKSLoFPY
BdvINrZJEKOWlUT/Q9DmbmTZEtXjeedfv4u2ruw+InbzT7TJJC9AtcdPFqKHuGICoCn9P8NCNWUB
LmVYCkG8i1TBXVciRdg2bg0ZP1BtYdA+fGMoSodVMJem0WtzwlCRVYiJp+tejKU7oejbCtLtWSlw
SXLy/2QxRGlUphECrc851h2mpQCt1X0rkwcE8wJY7sTK65dyAFgxQNXyKqtCyTqbsiRI5jL6EbD/
QMWwC58EPAaNS+1YvgvH2qpR3g9+LKIwRsH3U8hZOn7sFZ7u6e+3zgTd27EMSF/3NquSNLSL6mas
fLuZ2e47zgMHWeqtqWbQ1DxQw8tj4HhSFCGYHokGgmOljSJ4cSo1+yLjxXIWcJNUuxJRaPnXp1CF
B2m8nE7LfYZF9cVV2G4ZviYyRO6vP4nZQvtEGJG940PwXVNvuiKlsC326u8vpXOwZWrWW0GO88sh
tF6vzcdA+Zpa8no+jeeBlOJnPGWeRSj1RjSkCTdsq4XfFkkgLNpC2uWhrpdAsE+MR4FJmGGdiJ70
wUgxI3ndEGGSi1N7HdfoQ7k2zqoSiSCr/PfP0aKSP6IzueH03sXaX0JOer5KTLDsScqRA5l4zhSo
khpqJaLwsGtVktQW1CYYPT5rY+AJo8DKGdlShYv1kHP1Ikiwsw/PZ5f5/108Z7RH0/IYSnWmgJK5
+NTWE+2SU3mT7uwml1N6iMweNwWfjl0d3Ssq4DqfTDbE+E4HjWNPE9nond562/lCDJdY17UE+Kmf
IlPt5Fr1MqVOLD2q1+kDPHoQAwHiXGnuA/rYu9ct9eXMc/ZPuqckUNy4iN2dZ0Xok+9xigCWTIz7
yaHGQ868FSQoUFQCCSSpRwR7ZF7WwUb7AspTzVMg8EkgAxKxz2R3ovvU19Xiih3GuZyRt3oHxqZf
cElneiUabsraQhPjj8/Zw+Dsf1hTmhBQsofxyTBwuKQgF46rg/jpFxjQ5qMFPGaLHvHP+bl8HOcA
tXYTqCQNLgjpyZwtopbCygtkyYNQhDjwSHqAhg4q6VYhUc3NE0Q0MgQuAHcC83jQvx6/fxIJuw0x
FVM9YgxSvomEYDWydfmtYX1RnH/7MSfoBaUVVOmUK0fH3rHuLwNCg7+ZtnSz7HjljZ8QI0tXUsgf
YaVZ7sDVklF2yXT6JupsTb9KxIKWMvj8RRxh2rvjsI2niWSgbR74UKIF4msEPXv9X2H1la3l8N5G
KDf4qB0yaHifjzwUgSXvOWRiA/Acq1dlK7dLiJqukT0NzwK6vXz3CqHJ0Bqh5u3zJkaKfyiXAtxl
JdecAyJCUkA2PLWGcmXWCp7irbNrZBCddyx7+8hGpZPTRg57s3x0TOZG52HpUyqON/HaeBI2PMFI
ZJ1IuxHyCKsTYW2RkZbkl6+9ATmxPhUBUbvEbkRD17K5OIgJInvUoME2eMsZbjYzQyF9FRBz8nnT
pILHqCS6tqkLdDMcuBAw5IPD6AvPltgmAMJDyYT9VEb/F6MXS2ARHwDHrTduCDNVWb15ydyOb9nI
C2nlqPiWdFbrjy/xS+8+TCtTH4vGV9IMuQ1ycfwRZRajI13wANXx0+A7QqTH5G6IZXlSyC+9Ryc1
DbKm70bZ1IW9Y3YHfwWyxDnlmLpKfnB4oGOfPtvoUCQZ5aflunm0NbC/++B6VmcHNaftvHbo5L99
tGI9w3QWTNMj8RQ8sGmvrkAip72JZ/KZAjgdQCWZVLVmJ/mlUHw96YuGA+9h7cT3HbgGV1hb9Mcu
BTQCkAQsBsvgSMnTYcK7jGjyg6U+14SE7bUmWpwpXtw79zBdph0rTBv3rqrc82QHnFwtAtdtfcDp
Qr8eossXkPTu9iF4ujw5DL/ZtEKG+fQrsl3DFNL4CeL+Gq1gh3NGv0g71wEJvG/P6CXXzKezS2RF
f4HDgMq1cmgJQcbNcLEZsQneisXfnXONjaoNCXnV7vyVlnaJ2Dfx0D9D/yHfaESQ24uWl/o8Xa2/
gTVnUYYE0GGYMMdOBIbE0vkHhqC4zIVDzf6sfaDQBswGEAd1S9ZN9QscOT+z5HalZFfOdYXR0h8r
auAxGhzdNYFN/qp+BQcE4czjUcLvzdhUFSIs8799lzvtzS3Zz26MyN0RVtM1/Z5Z4p9NqNRWLvOT
g2X4OjTNyUWo6Voa3GE/Wwfd01/1OcV2IBOQWeda/jHMAvnRjWOJcHWZ0a0odGjM4fR5133AsU9J
qQtHZ8HOFhnz4ZZck0VQGn07ln7ElkYwqVAEmNsWET4LLwqPgOJzkv4Vs2sboyNqXRq8+NBDe/Kh
eB8c5BETcaJSnT+HWPaYCbrBu3SAM6qvKapGy28zSJJimCjGLXtY0dvo8zLGmSllpLoAfhSxZz3u
KO4zWlE+/yxFn4leFFxf6N6o6TkNkf36LCLhwMASu2BKr/Zj1v8HBOadIaP78O6W9unz/Lr6wXjM
gP2QmV3yP1NE16CafIfKrBwq4wv0ePqvrzqzadKCjXDRUh8THGE7UMEkAIFlSQv8mTacEQMP7224
Tla9Zav1AjXBvIa9ExRkE+skCg/RF9zCccMxUCcDLhno9sbiCimh1bXXhAZBGVl1JFMOJPQt4THf
vdI9IyBD1EKFr+/86R61QvjlgGUO36bVTDFOav08o/NlwK6H4UG5FELOLjuAWO4TWAoKvuDsYPNz
egolJ/JkzvLOEck6zj2AcWtU4SU1BLn47xveC2RGvotIEU8c45rqMxMs1m2AdIeXlFuf2Oe7eHWS
iHqOnO+ovsWXZ6Zl5i7WtczJbqrVkyr4CL2GzFuf1Nt0VPYRbeFdN8bfujhOFehVg3e8acLItT64
nvUPQEUqfbEWNFB+CFgi8VaOg5rPqPuNSbXmKWxSfm+tx5RSbfmlP8ANN06GDJTqh0V+CxHP6o31
oQyaAwLvHQotywT5Kh381hmHeSCyEu+69es6Rmou5oqY0Rs417ySoEL+1NYyXM7Qt8wG/wq1nZMF
BfK/dlaaVY4mkdMyy07C3XR4l5LpwPz0WT0PRS040sYyaMxF7J81hh1kLDLfuUYKWqKymjNpDcme
wDPZiUdqXKHSb+UAIU1EY60jnn22Tu05i8p9zRi9bAXrEwQEdLEU3RHpWl2WoaVp/A5Esr9R5bBN
A6lyr1PF3bb6o8SoaquL21uc9VIvfZe/a2WspX9572PNsSQzo3uGaJAKLV83UM/uyiO+dL4WPD4F
CoGdp0GKcWnMQszhRjg8vYwR8UTtjdAT7HG8AyES3ZjVxv3u8GYzOnMAyAnl6Zll+mPzYXzSIRlN
9XozfPrjTlGVW7v/8AcWLJTIN/9wAO2hnDKhTUDqzpwD2FHQ931f/L5zpOE1sSyqkgp8UTBxQJ8g
OdBLV4Ff9RqQ9o1pp9zf3aHX+i6lzEWVHrCdCEbBrl19DwhVYyEXEn9Plh2KPAqTLgMBnTjtCisE
jlXrLMrSlrbI1LXYWdt/4Lr1rMgRgZ09qH0iRogrzWETjaWjmGsb5OoXpb8K282QWRQezCB5SbDt
SEn2moadyCS8FDtrQ/jJTIXGeoRX9zAkhkX5s0P5Aq8dJgUmIfD5tBQQeOeJpV0unTFC/88Ancg0
oSAMOwvxnwqboaUA42Sru1sfAQ4u25ZCpJrF7V3/egfvfOInmviZ5KYXCzo9w1PNVYHslSJsr4PR
+xVWU/Q7m9PfER43mphILsrmifyp0osMD9Txdk5Y7DTkPsZ1nB2lLq3Ouo/8VE4Umzd2aeLlT6SU
TGP74G1hl4O3a2iIFARS++jRFdOPodwPcGKvtNtEWe33MKUeyp61LVFlORu+jPv5SyVSiKrCx4Wc
KBX7LczPrFcUlA0GIWZLcmSbdF5CGfxqWcdXTgm44Lnma510nTVl+/hYZd/PCyTKtb1mFyg99W62
9Qqi3yn5PQnwjKbk9bse2JRUOjh/x8pB2yghZxe4eCD91tD8ukNj818T8sagPrzJjRN8ZQ8VgZeb
Jlj8WT5T6mKP6Thmmx8ai9U6yUtNY+WSKL7+JGz72nbS7ZSHX/7CftvGwDxJNLQAZFUJkYsF/fKP
v30NUfCc34x5KNy13VBu8Q4s7B8uesaxFetxrm/2gbftVYY73qCQEUyDPlOao47OegpzTipzzlyV
NrfcgWWKOi49ZyRxhmFLUfWw7kXfU43XWSABPa2gn4voVS72KXPQCipDvP7avE9sfk5YTJk1uJXq
DSuO67u5H2+OGfyH3gweTux0MdCed3HlBddaJkH7kskA0zE1SdJ8ct4zvaP3BwldR7//y3DX1hjk
b3yggBB3RrzReycSYcKK/+1kuMdlGWyNAC+O0bqH/YKnqruw8RZFuTLWvQ9KpB8RXJVXvShwjbXU
XEuPqoZsqVYXlGslFTIqA/TGrxB6ERYHvoXGdumIAj5s3kARJ4yCBJn8TMXvaG7/qoKaMVezWNPf
MXY9pF8yke8FZ54usQlacfLl6nXbJnaku8HpQADAyRQkbWsjQTs4qUREbH0LqKjs61eswmIo+/p7
F/Umc4dTJKeCZeeLjJYrmcS5/bm5/A90oVmO6AZuXXNUXy7GPNxgTKuj2rHc/Fo5fUeRlTQA3a5g
2Ef7nB5tHO91q1tl63Swa2aIH0CpHyEKC3eaJU7eQmq2P103SB4G3XJy1KcwGCntINaBfpyXq3Du
jlinl0DzONk4kIN3eXrIxkCZAkOSXjNwb0mzEnBt9vzSV8ft+Oz0LtxxJ6J7bRUccC6Hjs3w9mfU
jMx0CYzGYwCb7bmRUhyshr+t6chOc9h8AX+qV73prwv1mTX4a6TZWB/9O845y0OpzPijEbOPoz9C
Nz+Uk/h5MXemqISxCfZeSdoHui51ldvnYqFOcNNg0KPSejKEpmpY0qi8TgfVTncLhKpyGkZ3bmAE
f4Vr5mzBCkveOLyR08tI/YZId0u82QWxzvy0NKE3Vn2hucMJTZCjQeu8ilGS5Jnh1A1eUloSy9Mm
eIdYWImpFBpChcIhv0329Rgmy3lYWb9c3NtbnqdmjhBodobVj9brJR3o+katLJU9bSCO1OIQYeWp
o9sQaA//ALFYsrZR5H9WciH9JwhZux8EAujJKUSP3PJij4rljFTkE2M5vkYt8EfK88GC0SH6469y
Zf4aqlrhJr2hm6b8nbGgJN3rQ/i5yex03OFPYhZALfXMsIi7suPQDyAMhujg8aKOz2BNKOnW53Gj
P9wtfctzT6rp91OD6xbO9m+cA1oVC+nQl9U4QlPdCLDtUTrdS2NFVmG6zGK52uuCrFnu3Vkxggk0
uqrvppFEYTc5spitOuR9JqTv9dvafw6GZ3Lr6hLOznFa3by2aNwfF4cMeJ2o4OduJQkH6usrlKfZ
TtWBo5WfzNqwKEY3KLYO2Nd6ifGkp7Yepa4T5Bt8jSl1v+1kg+quSza22TgjVGIC1Dfj/65q9XrY
pKMVUaYlcL79sSKKSHrIeMr2kJBdwnX2Ea3/NsgkQKLKmMiv2c/LsOciw8GxjNKhq2IidtgufKaZ
CIQ/pdi4PdDSwgflr6n856dq5q+ZRweWFLCZa64PpimJeSfunnOUvlyqODmfBhv8QHYqhEJ59Z0f
u0zVEcNGyisGYAj8N9VBbNeNwrPtmm8/ebehhy5Xah4eHrLeVoup+WTA3ZPtF5Wq4dtrmfbvNc7X
QRWqyGcYv8SFV0yOcyvyISIA/EgPehOvPkCZ8BH8d88Z9/4GQEziUnYgQ175HVwkBTJNNWHFA6ZW
1VTT2h7f1tiUIN451z3dRQeM/jPLPnFMOHrxqs/nUrSV4advrrXpYvqYu9JGLJNGgzQuO76picGn
/3SkhqQa9nXCrY2049UQ//P1jygqt9GHPW/EUfYeF/zlMKkwdmlKKrB8mriU26CczeTiFaQ6TMme
oQJ07OV2XLOhHcTSKXP377rR7nsAow1qrcjhMY87LrDmaZiGIgnsz/Sw8scnV5ZIrmdS8qkS43+B
WlKwExhFAHPz/OKSb5axWE73LrMw1pIJr8HeNjVKBoTTNtxokPy8hDC/7I3VgvQ6VJviXc7vS76z
sXo1iiYIcpD9FYjzfQXD7x6AVWwPnVOuNIZa1ab5ZHGa7z3UM7L8wVHfrU4n/SyJ17CD5HX6jjyo
bbqUtaExDveXgOhY2aKY+chaetlB86P4/kSRhiaV8e8j+sOK7GF+16D2Hu6Z+tnhrtKnaaDaS5MP
ULxsmhNwpur1h0nkiusvypIo5i0uFrOzhXtUDG6XrmLLE7bCoEF2DlOc2NYTJUXL8xXTZQObjltO
BgWSSQ7CXgj8qwWiAKneka2kxav4+ewKQy7R75BjVXACP3aXbweIJIirTQ4sqrFGflO7C4gY9FFy
2PI7Xqd/Cf4+R9AetZpaiGeymcByedd+WmBmHkedyJs+mOT/vV3ymRnxBmRRAqd2qDbfKdKMKbcG
fluB0mSGlfJYH9ZADuKKuvTaz7tf3fwUj11w9USk2mCjrz0TT3D2AzPX5YzazquxsAEtDRTkt3SC
LfhlS8Dxc2V4LkcdUV0X1MJn8CKNWCVunJSDJmOJd8L15kX9XblCslFqEo/tFNnXelEmM/Pse4Pm
DbMf70N0zZNZCquk8VUrOk9dvG9HswmW1S1mkJttqfc201gYhBboJf6+65FgOwhUuN77MbSRgGPW
G5TiiDwAJWnvbrxTMubAPTBu67bNRbHaFDZNje6iKrFqJCKZemEa4e0QF1DeuJIWnkW3uBJAR+bp
GhsCgNVcH6pJzfhC0YErmFpOaY6Lk2wsm7Jj2TIItCPpqjhQ89xRenbCkSHYiHDmCWBU2jwHxTn6
ic+yTlTUDQBbk8IAsSZvzr3yd7k0UPGnTnXzSDkJ3axSbwXNE5NEj2DHeTxlj/tOZFzYW7VBiy3/
YYPC+cpaDPkh7K5aSskLFa2FxaVUX51TTiOB6FAo2l9wADkVSRNZ4FWeqVV05J0Sp0BQoHxoeziy
x3zYXPNnC40iHcJh0NQs2+9bwC7Lmyj3vFfgIsDuwBzGcGRJjssjc1+axUH0Ns8Bu/zPHAAt5E+5
deS8snih+D0BsqP32wDxeTcuP9na8c/gbY7TEHCZVjOvc1LP8/vJdUlqMlf+nDnGT6k2WPyy0ckl
mCfb1gforVuob3KntnbFRi/E1YbCUxe50y+hTvca5nKSle/MnpMofvM9SLPe+08zJb5XjcZWuqKh
60Qc8nfvm0ZLHUJ/AtyP1Lh/SNPKWE1AGDghbN4mhBHi+m7sxbR1VGQe82uht7+GqaSsIs/lV4hV
0RoSo7Din1ITo7jQevzPN+V84wF/R7o9NdB1/rkwjg8J7hIlEWbymtcD8GPuMT8LqHVgHo/op3BP
6fayIwLyy6nqfvH3JPhBwzrxedTDWFV1yDuDqbdqeGfODvpN4ZVQ+MWmbhcrVnDV9GYTosGIjSCu
VzeuStG4PGA/MMzwvjEzcKVEqJAfKw+xc8mauLaW1pNpTBabjqqy3HlUBNu+jfKZ6FYR8RGgDuDf
HegeyVmQW820M7EMtEypYugYIVtkJHDyP6V9bPYXJuOxr4SLCQ6eyPN3Yk4eZ0uRXnxSf8Y0cNdE
s7ygrm8SWDexa81f/VzjXGhUE1N78QAC2b0n6C06XHH2u/O/kgJLWNSWAS+li1LdczkU+tCvMx+T
wa1Gt0nnD6GPvhWs83zPd9a3hUwERElzfhAYMadkhJR29FVgMWXKf2tiuZd5hphL5cvv1aDUpmZA
VPQpZPuwgveIlGCa36mMMt1B4P1Rc8z2nlBkTf104ezU7ohJKQjqEVQA9HAMnlHgvQlqhUXvL7y3
XP0TjRfV0BStCCz+rRE5YEJoVbV3+rFsP8NGR6oGdkX7mvvKCHQWIDo9TT7xTmf9F9I+Ga0l3Fmd
G5ZbYkDNio3xRVpdTjeLttrnFRAZg5hbLQo2E+RazBu42hSs2jxfDBBIGM4oLFtTqGwAHffYAtXV
5/Y877mKUaGGjWwR4Li033vzNx1X/WoyDYJy71ELodtwF5Tp5M4yIBGYu/a8FCwnj4Ycj3r/RN3C
jhm9fY5oJVzkZJTj7XvTE/yYZ9O0oIr2pSDJ/hYmjyLRvu23azBlfq/Zz5tUysbbntZq8e1+4hpY
yZRdndl04+UDI/gioR8j1dfbzw6Yfpn8zvoKb+Kz164BB4dlOt2F0rNDefNWPe3H2b3yU+4Iba+N
TX8oAaV6lsKs8p53pb+AByULBjF5daj/Hrsm9GLiIzmYoRv9uwbuNAZLGvN5NpX21efuqCsMEgSC
ksw9BQ5wEqbpFOKMHE7EdB8XOr7TCjObLRtZJEnLfYxxVyTbWaJJnO2t1/JYmWFSj4kcyF6dyW7i
zY88f5p/XEdo7N4IklUqLca46QzSLZd58zc2ddFX/mOTJSPcZVJxOmR5FE3b66D2mWKJ2B00IiJD
B3of59efpmcQGC+u0K5gBrABAjDhodDm9tnQUF8HeRuR33fl+6QFmc3oPzP1Itr+ZSQBRCN1Y6ZR
VtQExBuBExZsCShd15yR52cNGLSG8VkkerxTuA14W2JE7DBIlIZUaIpkgP3za9qdbXL5RDtULiuq
lZXKoC4hyJFFFs/KP6qvaDRmHZH+itbeFA477IENF57QP2lkd1g2dET1Ukhd2SSVqOWgziMYGOrx
E08nwJt11w2p3LNc3gzLOO6A+LV2XSbCHTaqxGDNJelNj5CV+5kp32uSmfrKkTXwbtdWC6T3zbDW
0xefRpyoOyYUNGBotGlu1iIpnWs1vw9jgM0fZLVUrRX4rzoYVmV2Usqga/V4XErvKDILOpSM3PXG
3Fd+Pjdffs4wGVXbEHdYMz0hkILOSzi8TWo1GdqJO7j1crq06gE2epAzyLzWkxdbSPHL6+WtFNe/
jG/w/SMtRtjyVUJms6CqHIKfbj7i0ukm6BwkcWfVa8jtNmKE+b84PribI4TKiM6ycXVerSWOYz2l
uZrRaRICekgCrn1ZuAzqLqoNpDqcrgaJCtrSIRyCivvGO7gxV0q1yYThtVTkzKiLhoL6KY2kd6tY
QqkTaU6vt25AxcKETsGK3cr1dPmrtHyWE5OvsuJsXGFpzOyANZ8wyLdZSqQ0oNz1ogEFBBh2Hh1w
vj92zJsITk8V7S6tGsjGiYRUeXuiC71Eq9avLGLC2PIj55VQB+5L74Goo3mvc3f2cR3Fbd+B5dW4
KtO63oojruPcwD5y0/kkCQQ3LqFV4WLaWLlq+wMxdy2pf3v+yhvUuqrkg4nEfJAzxBOeFWjfQQxD
4meUt+cvr4BB1RJyrz+MFemfFNCapqUxCEA//VeL3LE6tfpLeC8njJuTPaM+1uKh3nLobAY4owzX
NRR6v1d/J0Vd4dPsG78S4f21jRW48YNvvcK5iQ07hpIpX19ZyRDfe101m+syuk1uV/MThB/JhZTT
moLXBLN12Kol7ySJG+MUwnm/HGox/Itt3wAmjcXw+drmy+32q49MOW4VnsdHzkxeFNrA+E2c0vFZ
03jlxjqHICRwqwYWy6VbgTy6jmw93+MsWjw+xkhvVBZSGYF+rHLR3zl9krnxL+cgMZVtt16JqUK2
S6sx5k+5EFNUcY+a5tEr3aJrjbTakEEehNLFh0aTC7plnHycUypLZstBe5sjOMuCP2ZfMf2Oooqt
I0lgHSaPY2u/2a5Q5qQ0lvoZ6i4B1zlZU99QK1umpj5c8B88M2O0qfjZ2An5x47T3/nmL16Peblx
yFkbpK5OQm52ID+cja0IhmiMFD+bgnagHn7H93Uy3qudIolld1RpZsbmLfjJI2yXPdSEKZCiyDiL
Tc+sHlQLv2+/Wr8qZ5hktIITBRRw4HQ5FdTDMdWfhzcy/d9ZhDzdiWg1GR6yFKhuupQ4p1WITi53
f1SLbvw5LscI3TFUjcQpX3BaLYpxQeq2Otma6OWMQbzsTDvf4qk6dNDQJxm3Q/1JHkLRxVShXTbS
7WQMDXWU0/7YLe44yhYE6KPz6QZquf/MlkOetC8sZieeMNh45vVuJio3Gju17+n/S2bo4lBr7K3F
318Fb+lQwfscBvPBgq6j6ln88bCBLX9rXP88eFoEGVnTrCOftkm24JMvmCGRzxZj8DEGKSibVe7v
TsO+g4VepOuTynkbEG/xhwgr+nhq1gEbROsiAV+wG+83WFRrKR0YUYb6RLuDostslTk/Zo9EMm6Z
Ko+M6HwZdD9fK/8ObEEPqE+XprXIA0KoOTP3pKsa8vswLEbjVKpeSTDzC+WV3Fmh4JW662dmwo4M
Bo23oCHv0ygwzwRDYjEDxk9W8AXaSVE7G6omqrceKyUf3MeQ5szZgH0FYmOWdBW8IJ8tKVwkpYfj
IQTNg0BcUKvpF0x719MsSKi/ObCrFMc+e81FZGgsqHPbXIJPLURJaHh4korz78O/k5i/z9n01R2L
k8c7On77tbmUYnEmWQOnERCCDtAcZpQO1Jp77Z6WJE1JD55C3MycewJcRJJy6ghmx5gwGrHs6nxT
C4pQTCtnxJVtHf80vlcmsbbNz3LNJyXhNeD/EZ/EASVs4ZRIRu69n+ASNePxmBCpBHjqxugpfl9x
Jy0CY4v+3p0SvJPXZ9CTyxEjiDH02lAnMbfK9C63ABsgfAkHtWGdXN5D69Ez770dgGIVqOBxuvqd
6Uv2dDJ8HewyOVoRnEWRE3brf2DL03D9UKhbZ4agtuVMQMaCi6S7k3R9TJGA8teCL1k4jNjTPA94
XGu7chPeQBeL9QCM+jGyz/39/mPGphOpV8wuI7WYhYOIKHS+2IvUlzPhT/s+7zzEo7N+ZRBoOJ/Q
dAmWeLJxYXDOES81MXWwnRSm77d66j7NwlAMO/0jAtC8GNhoi+VfGHn39Un+Dr9wDX+fy0SJO+t9
orBJ8PqGezsI+G3jSQ2fyH/MP5TeNj5Kv1MXUed0wjvWnzvf0z4iP1vFg1C8R8/OoZRFJYmL9JLw
P4qKk2prh6NPEOtVR2fDJ60p032lHvGs2JD9N892sJpXQkrBMVXQqlAed3JOZQCxXg0ctR5SKiT5
k2PfYB9LXSGZmWv1Vj5q3BFc1DCfmYcgCB90xpMy1wXBBuowBqzBxWjC0bifVpYb7QWuOG6dFmGh
mXtkbl8rRmbqxh/dUhiCbWykF8+2PGlVsXjQ2bFzXrwLHf1PQD7BDy3JDd8P9848wYRQg+wVs28n
Lp4i7wNrSvEreCGWjjMGC632+udgpNe/qhP/i7dDehQyU3dIDO921JdzOa5EEFWiXrv5LfLMaNeg
gLE5aljjjZALoFagcw+bj0a/MciyHTY8CPBx1KB8ZKH3AeTypXW+02mkZjlbTt0LwdkK7bmv7tOF
6YQ+DeFQykOUhesYt1VMwKckzwwNwIG4g4EYD9H6vs8nA2ETOxPIvn0/6UL307P2S/hsKN3MfJ+J
uhM6YYKSjpz7dS7c99ZDqxGYscJRDSTomb6dZuWamJDkrpLvLeKz4wYlBSGdhL9lWdzmFcenVXMt
AJYfy+yKu8EGaHPlG2viThuJm5jGKVYCyIqSgd/7HHFkZfW+fNCozr7BJrNKnz7NJsAP/ZhfH4Je
vAxkbRkH5cKeusQKg7XcQ0ZbyuHKHBSxGE11oZ1fquK5Vjv9Pc/2edKY/njHlURWPGt49xiXxx30
gjaNuMYXy+yJriFJUyvhYx1PrUmPVWb/NV71aL8xM4nuOlhhC7zHrvElSHvpwI5mvBh9kw6uRkEt
jyXldL+VeFjQjLMVwvCJ5ig76KfY1VnthbIq/wIYG6g80BADuQnt4r9pIDXiOGc13ez0lrXGd68l
12IaMJnlp3GBIUZ7JCEOp2C8u0ap2ILLn3fl3UatQknAvyOIZH0YmxNJ/siSp0yYrKMzpZ4u8AAD
2I/ZosQm/wZ218xOqSZuAc9pvCz3XayN1bmoQi1HHi+ZMT+/wF/Mz00cWNgN4T8rhjh5XOOkLhZ6
w2MUp2TrM1z1itkpuB0gKGg1rNKRUO7Da8L2WvTPii7rlZ1OQfDXKsrKDpaTqAsBiVMr+r0i9kbA
RJGvwL1V6aeLzdLMclQHHecvPzeNaXiWr3Xo/VZPwoYuZjJkUDQ5PImUK5bP3braM+NyG+jWmfHf
LLWt9zwivfWbRvkmuaH4PTDZNZWf1l1LnKAftaVETi9+PXnDSJ5XP+kWgMcRI4/AdYmHZ++Xq0fw
eub2k34gNhtzOQu2PVCf9853Zpj3/vRd6KaFheykIHv1mC4CQRKVgiGyI1UqK5tgUH7EtEMM7AVq
jC7LQJsZzOoLgLNJ8/3YOrlNvFW94fPr1+h+p+i96RL9JSpF5QH1MNO9qzMZ6PmR79J1VcWkRVRw
H+QMki7hJDs5EYxgVoLmzEWjhS/0zfz32w34yQ7HhVqSaDE+JaXAEvQg7C5M3hq0M04DHVOIFtCz
a2HceeEIu+sP+dYAvnnkN6u9iQQuPElNpZYkl6wg6h0DZfQfL9lpU4LmHt+IaqnJYY5jTix7JpZn
exu/ZG0uvO6YnDlSSAsgEuZ6d79Lw0XD8MzqvqsrrYC+51Hevu8hhMzt+lXTyXrnlM0wKrcLZ3G1
WX9YFbfhtiNtnzv3l60+BCgLH9m6JHCDyyZ3uOA30DYFP55Z0q6UliHmgO+rsYLqST9h0fmp2Qo+
cJDwhEEPORGnFz4QgnGkznjwT+/ag4aXtQzpJIykX5jUH9KPRBTL0Ufxb5F7BRBBDvEPXCMekHWy
GvxVt74I7BPSF3UAxo+OXxpHoU0iLc2G6pmqJjyi0xzIoXtkXDWjaZoK0mq972Ji5IJRShwsRqM3
/rWm8J+VnerJCz2dWf5hOLPUVp8WfxwF7cCWCF2d/93HnzaqgyhfdRTFFc7NnCzoEar9JHjjpoQ+
hRV2LtdH74gLTYirsMRL+6OOOTfcc+lBkm2mQ4oLfBCGG3swHNrR4087TXpYLZqaEIU2Uefu5Uxf
32M+b0fxG3qSUO2kPXI11Fn9BqeKCybDYFLAzqKOxtdgTzpG8uvX86yYn2B2KteIcL2jYqQlt3Qd
127uLQpbu62nF7EXyOP8yFiRhYnDI//RKhjHfCdTEXgfCahn1pCOxUR/8d03EPiXvkex2bi8aosO
o4hhwPXWJSQ3GJxdo6FKn22bS5HTbZ3ypCuXmq7U3LTvIqwMZN4daL6GavjYmlg88hZ7Vu9y0aFK
+XCA4Bxct2PWg1hrIQC/YyjkAwwGjAWJNIir9pTQJ/IEqHb05wOopNbGjnLSQTPofUFMXhrXBwDC
9kh9MtIXreY1MVbtDf4ynAPLIQ1G8AP3lm4YE7C9NrQn+77OTXcoHRYblKvhjuCWCay3GOYoTYY4
0ME4NW5GItnL4JHjteNoO2wDs3RLcZiPTfMfH80xClxSsyLc+tRStEB9uYdEU54JiJHvyY1yLQ21
nvjgH9aRm/PfJ22Hbk4Hsk/Wau2IdeyyeEflkmk5cv8UNlQZT/VSoAcJvElfMmlb7bGNZH7N9mUh
lHGoEKwuQFEci7ltSvBrg1+LOvrA1fwierIS8oVNjEBpmg/QT/WPTcSkDHKcQFLLH+8Eu9dl9Tyb
PPvwGijxmJ5zXNChZlww1Wn9A3C27/ynoJ4ENFzCR6sUwycy8BVXqEbne5RUCLEZdUoSqsfRQY+z
DKGQL7+FK7KoRvNaV808IIOLooHRI+/t3bInu93436WdHXFQRkVZ+GqYHW0uqO+Kl5sfMjAM0j4F
OToGUfsu0koOjZzwMadZJ4I6Ga6W8rgQxL86G9s6SWotmHM4ZQIU4IIdDGc1C4nu0GdnbhC0Goff
8ebRWk2nE0FuIayGq59OK0m0IaMK7PToRGt7iYEWXXKwE70EEBeJa59f+Mb2St6kxhSMlSkJKuqf
PGmOif7xATc06+kIkApInR9YBY1oRIhsJp1bxgypLU8qkJbh6IaAGjTBofln4g4SR2U82r9jmZSL
60VNeIOMjULVS8+a2cuiQGd4lS17slNS683N40xXgv6csHYV+pHFNbY0IJWNswV21REJznBNUtm7
VzxT0vUYdow10pyfHlEcyRtPtfnoaeSJVAOnYWlK/rusKmRzRLH2Ntk/e5NXPT9HW0eDlffrsTot
SDLL4mY0BDPsFavX0C3M5JTS7pRz8A2wg35blfk5haVPydFgIk8hq87DniK5Yn76B56Ry1+gCPKj
4K4ST/FDcykWYvZAED/QGTQF0Ju1eRNYY5EOoTfimI+iKK9d7qsJxvJrljPiFwK2zc003JgsZNZK
eQkvSsI2Y7+VgCInbDWonUOKh4OVlduJFAnMDwytWHwG2aVqX1J2WNO25oucIsxCsV11o+LXP6LZ
AFZfWegzd1ZfL/5iVqu5LKUMeaGRlQ3R0IutPmThMt+fsRFQR0iT0KGZk224PiCgvMlvoxygMyce
9rzSXKwwDsE+UKh4T9In01G48VkJS21xBGF3ZrnO6mnNCK+iNdaBlAuPumYH4VhIPZl/kZkiJ3RL
7wzQlQJ+7jxrZf5iDE/39fGNcrHoRf9bLZ5zuHT4U5Ybpz3X/lfhzTCAEFTFNmapmK2Xt3J7glcc
6YugTMuZURPPCapg/o3qC1rxhIEPFHJeYR73nTCft3cYwVyp1V6YbkAETiiOcXfZBLYUGw3sNAmo
gwdEEpahk8akAEMC/6oDI2BLtyC+iH/Dg2pxcoQinkUtrU6ZZMFOtWYkSe+PYLM+sZ/73yZNy3en
DXi2LP8VpBG+GaY8xHaInZT2u3iNhtKozB2pSU+nfRajsrnNCRm6vVeHQxIN0MyvHrSxOWjw4yF9
MvNtC7qAiXfW40D12QLTlqueKIkD4LZYnEyVgIIVVzsjGg4Mbusf7OfyKL8dZNVrha8FJeRBP9Qq
5ErPXW7lxUkJF2M/jiBaDqhr9GCyrg3JyYWnm09U3+Su8TYBDWTj93gUq+3irPc5HYxhIlTgQLgG
wS3qhl6BgeytuBpwpoK9hSDVJdSCwqQ7OdKvUcwPKpp9kkXgQ/V026GmaGZUaCgSKtLU2kMdofuC
e+zUzRlynQst1rsowsxWg81fvO15RWlD1nINg0An12QXqBKm3QDtechJmGszSmqiFRNiT2jHVL9R
s/8GS/wq49nJpVzW8YdsQngf4CJ82WSX+nwcZlHbiLkI4QniMVjCpOvg0ekertsOMrcBJS8KQjLC
Yofl3fIoPPUcmG5uHgEH5Eo5IFOgs5YhOF1iF+AyLjjYdRR+LTInjifqk35E57In78FTWMDPuDEp
d40z8g4vUsz5RgmK+QXN85RsymsBUyewlHQSgblg6iueqFk8dzCBBE+SRlVJZSby+OaXVWSog8Aa
BXuEZOXe9T50+SpZYUx8gAwwlKyizLzVcyD4bxRe9Z6/RBdhrw5561u/Rh9AlFm/YN+lg+AhYc9a
26HHjNpx70TWuk8LR5BZmiNZ5gZ4IsQF9lTogHdE2w4RCFW860vg8eX/zworYeNll06yK+J/bOqA
kDR+o8D7XS5xWxfREExLgrXIws2oQeKLdOoEbymWA9pF3domm57Nw4XjCVgr0OLFhTFCrz6UU74L
NxsIutSJY6BXtpOg4v/TPyMrJSfAZCCMXWggboCqn3naTIfr/hXw//hmoqbEFrVRNoI/WXhylmix
zMmlhTAyhsnrks2o3SvT/EcgrXywQg4/51jY/rKgEptFkl+0I1FLMZZErm1oPI2sHSsWpvzM4VPM
KzHvEqhhffsYojksuz/i5uTrQf5D2NWIAkH0Z3S3ixcqSeWtYo8kiMOzYV4vu6xYn6kWjei6DeLH
xzNJ8/UWGFn7fdIiQdnJ2Wfbm78+1w6vc8wRPGdnRNqNFP1bSM/4nmVAnxzS8UVyHw78bPmN1zuq
NxLxr+mvGv6q5ULY1ncRHBjsdynAXyahTUIG7k4ITZ7eyG2qE3/T9fe2ATGg/htY15suXKCNJiDe
k/3x8h48FWewB8IgiDknFcG467E8dt2xULmFWXo4vhC+iVg71sm2EsPNMQ02J4l/Eihfx3aZTOI/
XyfmyKgVgcvcowMwKPrtZZUycpL/PWbHgN1oF98rR4W0Y/C3FG44HBAK95MuPClZu1e4KeB6fH8D
CPJNzd+r0IJFncLx1fRvo2lBvFmbK12vzQvf4497Ds2u+xl8QzAWcRVCkRq15z/fPIo7qpYiVQh2
S6fEmmiFbLG2D6fGGdOMTU0JNAo+kTGKz+gJh6QJk7tcfvScuOl2f16JOylqhTN0Dalott/jhRJD
qxLYSNPGG8Wp7pMEY/kKg9Bz4xvBrUA4MIwBCgrzew2AP2vqBHJYjmbQ5BbaIxtjirHzq2Mv/Nmn
ehoMC1I1pxhRU42qz0dqP0RT+i9DLdDphQIGXLrrrvNeczG6596BAvJPHGf8pCDo0PuAhVs43WbB
Ciy6yZS2RRLO9g+/PaizhKQxQ0tscc+u5zM+fOWwYYSd82DZVxgLJeM8FVtj7bPihk1PREfOLjes
0z7garoIgdQ7td95MyPJk+4BgPQuk4hQbnWNPHjQHJYcSEOucDPfMuICevoCvOxmxWHTNTVhgWwD
7sNZvLuBkcTCBywhwow5LBVdfynw+btt5El69Q8xlLZ7wLo5+X125CPctPIAUrNHkhYpLdu9NP39
c04LxhBtro9xdYRPFjDDPq1xpZRngUjgdKBYegq65p2UGvEwz4qo7bQpW2EfLK/prkS0QaX9U4kB
XuU82Vw+x2L6qZRftaKwTY+BmAJA0AzDRf0L0xHEDU75U6bJ1q9vpQwtlu1iI0BTyBXewG4/G35x
GoDQmL+e55py+nx8+PylPPEtj/cFGKtYZRnPhDiMLFfNO+lx5brC0e/UFsKR4sit1RpT9MDO+6Rp
leQoDTFUOtq8wCJ/wjcChNvoUFqrimAHJ1HHiJsbhd6Eb3acD0GSCGJDh341ClsqHLLV1zhBkUNs
E87lD9Y/kUYEjRSfDvsVZjOvo736bX9MyT6oo/OnnHG4Psezf1FV7kKnbIjwuG5FSuDANEbcuu8n
5JXM+0OVxJypDBZ6TIdGWgPUnGuKWJs1OU/lzUg1jNSdfoPPruLhOYoDRBArDsSk6jUTkLMdlt+b
JZJltFmnZyD8mLD/O79JBw2L3E7maHzL09szyXSSaSo9ZeDU4HmY71xEgy6wKj6rIY340HhYLm3j
JEYUovp/ht3Mk2EWkE+zmN1ZQzgCmYumfi0KlVjso+1DjPexaVzgbUK7NVOqtO6ueaORBawl8Dj7
nRBSxEixzBv9raMxiREYmbOZ53BBjgVq+xe0/JBasL+krjjsDr2jW9MONXAT6bTLYdtZlzlsygmH
OUVwGEsnEHrrJbWA6FZgjoO53Dp5EqgH+qWZymG5DqU7AiJ21T22mKCiyR2sdEURXSAPt5Dn8285
9uxLLD0Rcb/9D/xlbmSLA5OQDvqpWKnNVrX9+Uie5eSK/D+3polCpEkpGvjbk9AxCJYjwkdFcghX
QCW4/V1062YbN3eh9nCZnB8BtEj7tYmF0OY+fD96Vgex+5eivlUwSU4E2zMvyqp/Bhuu2PrBpgam
COiaPxPK8lzTfCSxsLHh8WC6riWaJLKcZwF0AoG9CCRwPkYiGIZcmnl/jrtNxMLNbvGR7wV40Egu
sOKdGkl2kxrs0af1iePNuEYVAZH730rZLo92sD2HOxPtSf/CC0mRXUnivugeCMqpwqmUCakEa0Wo
zv8Z/VIFMwKzZsm6MczATBwbdQqndzEDMdA0XDnT7Y/QWBPPWKALHvJtBZwjfzKeRnOwpsz2tRhc
obf26VeziW2LRYdTPyHiQIZ796HRZD+R0H6HyUyl1qAi5mSeEQ9VnEthl3MsFCH0Uo5trWjdGBN4
FzrO/CTYwOsPqSNTRHmmyF47DI23/8GUMVLAt+J78BB9Yg7U94ZgaWpe1DyCbdXlvVbC8sw9qKv+
F3PFwYGD8fWwt9PzcvsOE91V7UN937UN1pMqtNtH2QOXG3a+lam+L9iSIdk2ar9/jeeInXBO6X3N
EM2GCBb42sgdHelGdsLVnJkxFbjIgO7zkqe/zVfWt8NeTUD2gxXuQd8syhFTqsqAVCzJPBsEUS9b
WMTMvW1xjS0Nioqz8iiLzR2j5HsnrIxWMefyYRN/rcfOYbtmpeuxlA0sWu2gyTo9pgiugoZ9Wne0
UaE9jciGicXYVqdUEZ73FqHjIwNroQRK/OFTYVlrcBlF0/o4wX/NW4CvvQpsaEttnWRgeWd6UyKa
LLpSPCYGRmP1QtkFiqVUaY0597BktNkxPfcr2PltORRF7Y+JSDobRFVel+5i1cO4BTPmWIeJaFDX
3+mf0YIGUbWkiarsh12pDiZENqCfOOa7IO3Pnj25tZqjJUkZyiOjdTDIBs5QUG6uLmJacBymQVPP
msZzmq6ZQ8gk+bVX9krnxv+g54ZM8bOdKN+FgxfBlGqjdSNv5w79IQ7ukvvgPUrdAHBXcAv0S7Gu
GTI5jRsUcdNYyzO2LDaJnLV6JBPgnQKpiFTJE7UPGk/pOAIJ2Uu4mChOxnWZwLie45r3GYpmyRy4
S45gN8h+PVVMn9Qoul7KpdzI3j25vptGeN+zsSZLSpeWrHsCqC3DLySAwemZKu8yolhNx8Iyufuj
xI80rcEt8hqBobB/6WB3iffYQv4+9wcF8B95mNVTpr8QrpEtcWR/fI9Vfa0/lKhR6IlDpZ1dRcJJ
h87rroUxJVQr+E/SvYWszefMNCAa1hyZr0AueNrRBXGfyIJ2TFE2U71YxVcdBW2iFP19i5EPZdan
zaaAes2GSQsjqA7GVJe6YK3FiRipU9b1smGI3A44LzwVMng9iqTahsvs67x4qFaAx4+XzuAChVl6
OYkhQIQBGaDS5tjobLNwkVsedNpXQBoyPjtBQGsgYOMYPSur7b3msd8e5fippP75NFBJRUFCWzNq
Dv2vVT0iHoSwqOtAiMmnE02/iLkiojch+PsVePKqllYMqyTaeQnEQyQv9ORCbT/heWamw+dW5ZPq
pfDaj+qc1sGGsrIOH0byFw7v6oAr1LF8Bw02XYXlFni0P3C3maCmvcjo5Pzq6QAsSc1UlLbd94kF
Rw9iADVKwWS9t32RX6qeB1EIyiU9pglEKwrhGwoYr3KFucT0s+pmiuog9UeLeUdI9MBUIRxVZG9c
wBMWeTYSXIaDyiy2NLpAzQHvBlNzgBsbBFBPJSgUXBcAvdaR3xBCBsWNTCdYCNy+F7RU/DA417BT
AcBvYN5UqYSKq7M5fzyr0nZORNQ8EJBKUSRfof7wKzbIj+MppiM1kODJlvZ9EE/2v8REVNtK38MP
pBjSXx/twdkP09SaMbaOvLFLmPjngNAgYXmQIeOcAJ87KY4kfisEUxp4xNION+LnleO/G+gH7Dp/
FBZ6QWM0v8bgoj3Ok4NgZ0LUyZX6d3eX5oJey4NG2AgBa92OW3q44yEekxhJQHjAbSk3Q6mAU2t7
BEaIsjH9U/L9BcDgBuZ9rRDKXs1a+qqLMwfDCB8bkgV7j/mW//7mLkqPxiCIRNE76t/P/kleYWn6
02pQQD+N1yNxzJ47lyggubWA5nLyQuYMLUI3fk7oXnhHpEl8WrSkDsmNAJaE6H4vCxVeZvBOuktU
tawQRYf/bjHhAh8UT0UwY4ynTvA1QQYHg1GaPELJEAxSicM6WBhnEglDWEJpxvjbXgwKzL3zwqAZ
YCAR4yGqHOhyUrJFdoAuefVfHhR+s6elg2kDkC0tmbxXtRHfDeOk9gXIzzmfokpt/DIakakmwOEN
GAJhohD9kYqmmjMV2hPj9V4JgiLGzeUEljrW1ZBrEgKz+OrkzIpcL6OHpOOM82kWn+pehm63E2J5
EHqMNoM7/2ccjbHpzABMhjpwEwkpLUNIuUqmrny0uwYYUn5XxML0wr9WRp7hupQwdfDlmcBnAh0q
gspWxro+PNPmvEoQ3hVXprTuY9iDZkurtvg6v+M+oNmuGQs3DpF7Q9hR5Ft70UoTD112833+kgKg
uAyXtoX41skEzG0nlc1gWgI90XiP/6b8Ss4a4DQVb5YHEY4BWgaenOKhLf5k0+Xahd/HtO5jxcdW
7Xh3zMpVE+7AhsQechlZbslWuxe1gfeWqgKJ9KZ57OLecsO1JNIkKo9r6grynvmN9KGwgL4NNdap
eC7DmBfw8vEOwkEs+R+37SM5W00FdUoBiZaQbZgNm6ALNw5LzR8bz0NSGXxrTCpX8uo/gW2U9xiu
/FYuZ2hn6nC8oRg7l7sJLQisrIof8G91X703jUsBMBJiIHx6BUGWidFZxOZHSQzCrEfjydmkoyoE
TFs/2Ea5LUttEjC7WHu6F6jHchfas0HMwqSD/6e305sKW0/Fq1SfJNuIRtYBr6vHcgTJ2Xrmud8w
nqivqsLRHYmdqCyZ3aXfEShvLLIsB10BcKDQ7TtCnd8dtDFkck1MHGJOz7JHrncHW1LcqMqDp+Xj
XJTqKgolLFUdy9vklKZd94/6yMONwYMKB5H0P1Bd4Hzj8GJ1fJ4SkL/+WGFVAU4jX5VFIyVwT6cb
E7jZPL+EYMdp9hXCuN6MmruY1/CcWdxun32QwMXtnFpo13RRyKzIGbGLpXmJAYVDFum5HThEF4Fm
/uA1AzGFvHE/tU7lMCu8xg9AzMpVdkne7312b83K+j89IL3umMKHWYJOCvea2pGAyEzBO2SDYC5t
q0omECMvu2+JhSWd1A6wAo28QVH7XOAxEuA3wMpkJoAG4P4YJ3otutuAFLElo8o3WI/QiS6URKZb
cdBsUbw6/ECcTlvwHnIj5rQIO+zFI6oj3nLdS7LvUVRgb8ZlZYFOvPD6xXIXM2WlaU8B31mjkMmw
7SRz5XWtxloSd9r0PJDXwVKo9i7yYhFUuM5GiY7Qe3StRIIXggwKJKM9EMmzUrzBPR8qvzeuOskF
BTOnIh4LlV6ej2nVf5xsGJraADA+3an0IqvQlbvPbwrOb/2Ofm5FSKFyjsLpIet9Y2b/THZiwl3N
lBtixd7IZoStmrJN/Phmj+AoTs2yNGXPhT/XepehGyv4dPTgDHIkwhAbxEBo4ljIZBYKzqz9hV6P
uHPB3JEtx2nHnjn3eRqlnd+sb2IFQC4RA31VKvhkDw3Ft1v9NTL0W1yWm8NscSJ8j75nutSulonS
82UzeGGpb4fmpYxGKN9iCYrH3dWrZawvvqz40CW/DK6ynFwV+b/jxR18heOCeGbLgD9Y10K6Wm9t
YGzHSxAAbvcom5VajHM40iU/K6Vt4KmIPjnBVgvPM7z5tH0kdVcT8KNwUQgH/7Xk0I9gvFaatfOw
yMn4tUYjgyN/n0qOueDzHlF/3ItRDbMCRIEgPs0lfek4GMoWaLuznzTtX53wepMPp4EmthZlbDxF
cH8s2rTJ8zyiFQtoHZi3g0EmKLNEoM1tBpUk6Do5kfsbnnOGXtLzn+SEr7UGqpf8KvTEvV6yXBc3
R8beoQgoAXr6guoS+7KaRoGx9ILi4eQ9a4of7gtczgYDCnDSk9FnYQ6XW6z9oGTKw6OtZo/fjgMT
qDOk1U0KoSRxXxbyTO/dFFH02lQS09QXQQlgwtwuwKbPhkal1uWGFCfbazqI/j6y4CKDdVLMOVVi
ztWlI/G2edKj2ve+EyRPjOsgLSYurPRGNW4WEg8kDYUdQj5Y/tKP2dDIkN/bLdiKMLi/noptJg1E
fyw5V9iJPT1Dg8LttLMmYrT2SmPzjrhczoiyiuKo5qbRID1oIXrhBqU9GFKgV+8uXor17UHNuDIS
sKF8Wsekfe52UcLDgHkdbM+dh5NgDVTymSzcUqRFLuOE0ep15zlaOq8/tyUJMOy6XOFcj823bmR7
2ioJ9DOccRKdt4jIoNGEQWx8QKPCuGrQRlgkOezNFANMWA2Q3nXJuX4/rLsH9nrvf8CRUZw6/0sm
2emWsj9plYCmXCIi4F8d3taj+AngC4EdIXICZauFE//xpvQ7g+PB0Q+WiQL1KsoJooV/ZJIxWfG1
xrCq3yRIQTz3M9IiaqK00C20iQ7B79TmwId4KKZakZ2+scslSm5T5nVFvUDDLjA654STS3dnFNAh
TxGUhqVCfOhKGZhV7JSSVfij0hLRnD6/pHrH1x7uKIOs/Ok6q1mcdoUOTfVxkbZprE8nJlyd0L3A
uxqAS3EZHJvxHCvPH2fz4WJRtsStEsV/kgES+gJPVTq1Udmg2kKbDGHc4lB3RDFcvuO7CJwp/3Y0
i8qQC3+vK5FRJbjc1hWEBsgarVZOhGSf0vg4AdREV19gWdLjZ5ulslNJj7QiORqpjUe9pEgk74tv
VCx0Vrj68eUh8RouTHN6yw9KcPXU4/GdVhniV+9Zh9FIHw2FSeZ/MFwfSVOamAsOZunhl4l1ul8J
szbGBKee4NkkzARx5kzUAPTjRaO51ffrrG0E2+QRi155uDNQ0x1hw/qUelgYfL+KDjHj5kxpF7YC
2JWzXR7Zp8PKlOoDR3K7u9NpIpHSyh105I5vR9BegkFtx7XOw009D64R8AvzoA0rfFAQpHhr8mi4
FO6goQ0xzTXePv2laCmF6wfxRJZt8fIle58OVBZPoGa5m2O2FQgH1JbFQIFhW3e1w8kRBwJ93DIx
EucNOJlYyrha7ip7sdfgL2MeQvgqfQcmoUjd2/xZZN2HhA9Az4dyx/ZIEjuPkuUt4eB3mgBaYcP1
dZ9eq8wYIglZCjf58ibACCH/Rn8Jm8uhDfw/OerkOBQFmJ6lNcy+W6FckzXpjTR5Pypu3uPLkUUK
inyeMuzd249TnqO5lj6VPh2CDXLvFjbC9QyjsVY/7QFtZXojehdBcqFd/o40TJSWsQBK9Bnm1e0X
fTKrfmnuiYwQ4acCvX2kaZ/qoUvkXpvVQnyhZIpU6JVvpMLRwno8EFcQ58DTd3EOffiULACzkPZI
G+5/qjMYg9Ey/1F7pCKtzA59QsbgjdMdnZz4e/jcDVujySVFoZX6INTsWDpr4AHa7vZntEHr0ycP
dYh9CjPGgozQyrmWCUF/4lvG7MN7OX/8JHUbxIjbCh02D7qITpxYwCmrn95CZpAis92bIe9qP2zC
lY9uI9MlNwd/VoxgDVRoxJaeVMs+n99eLgbQMkuIyq0jjoDPnrDP005Zsc9bILk08UgMdArdiZ62
Y1c2C/KGcks3F8lNdwAdNdu7M4ayG+C4DRxMGSwMFef2nHRgtnX2Id25YYavMvEFatyue9edtU0q
aN6x5kjnuX61UO1gpWk0sMlbIoox1VT+yC9ryVLYy2llYEch4jKwadPN9v4MaOQ+NFL9eUV1GM/B
92DNf09XIZlbOiONRbErtaQB5r5A1dizJlJFRLadrcWSX+SgiMiVTWRVpCKAiWqsgcIIVHJPsi2O
ZnA2pP3hVWyu7mFjffcEvUx1V39ZZF22cLOUthbWuo9/9L/7XczVFov4HuWuBp62GAgmIOuXNDNX
jH4r0eCSm5dgtyMsd5WR0r3gSkqXph4UzWyhj3lHGvrLkVB8xs+wMtChE4w/sUvl6aaTfT0x1dR7
uuhhTzfCM7kIZNznqJXLYdi2Ua8ykF6eYcHGQq6fM+QBbWTHf9l3LKHnySeg4GaamMgmx1HFxVjD
wR9aOPX2nEXrZdhoQqXG7ywOozXtgUrZnYZZXN2celeJ3yry9jeHGPqE/emxHFUAFHPLs7q3wmW+
mGMdB0wXa9aQUI25eP7Kn5IMWGlWohInXRsu8osbrGtaeSw4XhnmQikHKHwykKwbPhjG9kfpOZKg
t5nv+nZErSp/YbBI5fov1sWFnghsy4RBhbq6rXD3NMLSfStd2KSZX5yUM69nmEi1m6Krg25YmQ/N
ea0bLdle8WiHFiD/v6LWfa5mDDinx0cpSyNWSosz8T3Dn/5uGfN2JCj+xS1u3GQx0s7yc0Yo5fx7
A/46hqvBkh9plysWyuxHakRnrHW43rDsp8uOemHJTU/D0M+IgwuM76oNhqqSt1KQ1xhcPyxuK07g
egYA/ar1IE9H8iqcueBVFIkIPqtLogHx09cyMuWJnB5SYGlQ6NkVRAboUNPUPe264zkPiQLoizhQ
rTfL/q+PeNEx6Pe4wHkkFw6GQB6rFS8yfgsdFyoBn93KO8QyAsK6Y1jM41kWlX+/R5tV/zVvvgax
urT3p+htZTJyy+zqtQ8P4z4ZKl751LEPHKFEBAlEYCVwk1M7HUWraVyZmbOfO8Cf2ZSI3UW/by9t
RSVeBeHzgfbfo7y4pN1rF3udKcl+m0ElDlhZ8PuOiDsUvoYjOCTO31FOvAJc/aiVDOsiEBCXK1vM
zA55D4ditRQCDn0SECTQJbJ5G4pcmCn6OCJGLFz6JpNKeFGL/ESNcp/E9f53E7zUXa15xK0SuSz2
PdRci+JoSIDI9W05sw4gPxZBPgBdT+fXF0JZ/InA+hRa9A/DcJ0NbJmeSvBy/P+mWAMVwDeAsdEt
p7feB3oeoVehHANvAC1r1lu3iw4bTrwOjveyFCP3r1CYM4RfRz1VUkyL1h7dxx1VGOy8FwxJXrCh
Lx5S7mGVWc8ORdKJt5XjXzknO8Pxdnkmr41U7fG99eMeH7WOGNpas1EqNCZVwN9bAoJVgBdcE6Sb
MGr7I/8Up1R6q7pYuylEG/Glb97jbAvp1xZfzT/vdUk0b/7T3w6KFnWYJbnmQgacHOc2omqan2si
FzSX8SIFiu44ijkBWeHpU1H7qASjvy+rR2UWwkDobyQrGEVdGLUU4KzCS3pi6MFbYG9yWvAWT01V
2ZKIuYLDx9nzYsaOgnVahuE48pTlhiGJB/pls8uaYjhPPZC7Dn5NDLcJDMQLyZ9oRbTtwNVmekF9
uqoI+eJVN0KJcG0f+6koPZs5F/WGHDHY7U8kDkUT0jCOZho7J9UOMt8LNQZNBhAH+1a5E2THzBTc
mqhS6JxCaJJ6oKNOI0xLl0+NdstKL8XWJZSkAVkseqA1kK+LtNR9vzBl1qoajcQ/ocTzzSdKJuab
IpNPjNnub9gJU8wipbYk7f7UIBhtWVWFl3yUrNEtWk7qpuwBwyf4krHZ877hz3foRR0xaOzatq1X
AKb6th+zewg6EPn3/BHPYIxYP2QhBf850SxhdJJAywe/D8zCq60ZDhVoHaomROdpZoskQa2HIR1G
YBNBqBV22hd/9KngMxDkhn0ic2+sMwOgJd2wvjAcp7/SqcQNVFLcdZ1b/epx9DmI182xGE+ERi/w
3Nb7ifaxra2RbKGTUXw9qxBhnbwt1TMOFD+ocfqNMDaDBdQFybDuhOzIGqINtlbxYrCYlyLYgWK3
szzumd+8yecbt/N4LT1D4BM/MKLegQmaCq6xkyYykNs7/t5ruoV4fZi6kldbvLhy0Gw/zwglpIZk
lj8cRHGvyPWcXHucJKS3s19FSPNRS6eTDtz/P/0Y4qU7+WMIoEGVWNmEOWD9hXeFy5XUERIIBwxE
62/WGWtccol6I9lYa5dbYjJbl1RERKylnfk2GWttTgIIbt/ttGm88luFRV14W1vKqZWuzeYkWCge
QccQpXSomPVK2EincKNfrhX7nXMfG8ycfAQC8xWsTJZRS0BvwBF0CbcfIT0Kf9+G119+AgbQo1hi
MUQaMwhdDooajI6P8TBnVDaKspqk7IqUHN0FSSGQZfK9FoclUBynU7x1OqB/XhUv7dPqWEbMAxKX
2mWeGkDvBpZ9R1UxA0hbjYVi7bgGiCKzeQ+HEV7rIdryBIyAr4tscWsAjUsgQXY0hxbQszqcr8eV
PIP9l5PuPjh09uhjzad0YVfeCvrZShL/eLTu4RDBdl1yiIIo2vP8MuXNymIg4LB2n71T+wyX8rk9
Px1AibOGryLY3eqmQ2pIguuRMNgexQJqZxkcFI4qgTeUwCi1n4yaFJIw4JSRA3QVELfNRfzJ1ABW
/HezaMocSUFbrOWtECF9F87DFe/pciAr9s+IW7pdd812sELAatyFt44+mMLXHzv0oLbmX709SAFY
2ylOzr7c0eHKCnAyAo4jk7XnkNvcT1KTTtZQDqUUjt42oq5Ahjc/2YXTXwqS2OJrwbL5+HF3TsyI
C3lsHNwLBEr/m+n0KaLyDsiwzRVPHYB5ww8V+TiBl7LN9swFfC+26UDh2CQUiOwFR7KqlIfH1DA6
6o9mWChymxesmq/HEyOT0VCm8+H9SyA6YGin9w6SUHkpA0e6WPysyUakab1/0hPIj8Il3rxszJ+p
pVkKi+uJG+7jlBd7yR90+yH0vboUgonEEpi0uBUGwH3PuwN7BhncWVYCqnBQ588wbdog86GytOJN
gU39PY2MtU8GkxKMTOSrfjcSwzeWIiv6Iq1fg+an0U9l4Ewg9TtbqG7GK6ztJTUb5Evy3618nPFd
JM5uFyO4nQG7+lNTPc//7Kzr7FUIjqo41MS0ZdoU85/odpC3FOc5qDE1k6L0sn8w1MDMbjeqkV7h
8zEQeRySn93OAXVckPuNY9TO7M0MgTa8nPw6Ca2xy8rhPmZajJZNGyodZN0e9mixuPerkwzO/bbe
yz9JNqF0s2ofM+P8MoKLg83AWO5KmvyVG0XHIkuhu5aO7O7YYjh6nUUNDLtnYfyQOn6zWQnZmiV4
FhlpFlvrf8/AjLjkr2JCZ325foLSrtBMZOMrz8B/1mzsO/JUFB/LhVcz6LCQ4UfDq9I7RZnS7W5r
nKMgQjDcmG0FSCq4KZ9O7AnBU8wRoDUJmxa4wv8prcGfep5KZ+0BOJ3/KlRHFf+8de+/gZjeE/Kz
chqhjzsSCaVTqMKRaDry5B9OSz+Rn1OQsdSpfi7Q9yDICxlojJ2hgH8yjI/eAlWZZ12a79qtL/LB
68WOz05Ro5Ox1htI1z700/n/OCkfyXZc4gIeV+3YQDpCbrkZgXg1bw7PDaeBOdMTYwj/odt1spVV
h7C1vbJ/8vVpy5lFWhQp2ajlAsfsmMtsT4pE09dHGq9alpCiObl5Dsp+W8QJigifMxKeMFwabiSa
rBvYkpmqwXIJYdI/biivpVb0xv6gAaletZSGlSvKLalF5Kx0+RzTuSzqm+7r8+XKitwuYEohZSre
lagd5aiuwOdI7ow3tAPXoWKEEdecz+iZWzJz4D3vEmgho2MzRtbDA7Rs29GBKoLzbCk270FwfabX
u1B9FVC/YqqIAfpf3eEBDGsy/4FU31uRj/ycBEh6HUNGyOnZ7MiREny3uZhHTBrKBn0fjRZQD2Mv
dv1VH57oWo3uKnUrOKoQ2vgFA3a5Nq0ASxfbgwykW5mb8NO/P1f1lcqA5+RLzJk32+tbYRBmnhNz
wtSetLCf6CvITfL1iNjz8PGOzH6QuKWnjYEKmljjCFCogcjX2WVKBh+FhRj2lT/eyMlNUVrcrg1n
T7QtFDfEdx6SGbOIdRR9R3Bi6VOWpT4o79x7C+4IVIsdOp+po4JC12yIecGo7Rz7DGpAMiOs8OTz
S8wh7vTEwgY1wpVOkAibHA5jQmFRBOUXjpsiH94EBUVt6WhOJQFCvW2WCbtldbXLZiA1OUU/gUqM
/OkQi5PceVdzyw2Psqk1Dy5OqI0Lp8W/rkeXYshgDKxH3oZv1zswOcndTZgKoeKyqv6u/gxyKbxO
vO3lxfsBe5Bv+nCubfdDSTc7RuhxKo1RPGPNRnuf6+Xzy2dCjro/8RkJhL9/5NOCt9aqqfH9KwNl
LTByPqQitk+Y7aSKagWwcbx5fskCueenGc/Ml9io8hkcEn4lHp3fstgcm5g6ZyEYwT1je12PJ9NT
56ZCcxfo6JAnSXpw27nO/UQLt1UxCCr+ngsRnFlbFPHtEvIx985Be22cOYPmWhjBrY5dNdMBKV3Y
5K824LJ96n0S5DyOqYyM7WtjTNIqrkk3bq2T2zZ+wzWJhDfkTK4xlj4Dbqe6/mqn+rr586HxTBVB
8zJHxzd0/EoVXnvvDSeyT0YWI7BPwWcVmH/uh3eCm9Veq0qjvenXjI4eFFACa9kPVgUXvN+tbJsj
E4+R4biE/KXgs1IemIjmaN14mmhdZ7V3i3sCP9TcW0QKcDabZAxpOsC1xcvpEsxG3JnWg2Vt4tR7
SBD+rxA6gO9Ci7vUwmP2ywHdGrdLjN5e3g3EC2hXU1V/xF0IhJpv36aID4R/Z2C2F3jN7IxMY6QY
y6O2PR02H679+GRuHKX0AK04JsUuv3EfaPFe6e8/+N2z7irQBPcxpEkTxLI0jgITEJgOqfezULcX
2cf7pjsQvJG/mqyBLgqag3rhY0oGcPJnKQLYHsy1c8xCiOR6fYqn60jafL3aLbZO6AFAzhmCpNW0
0Trg8IaOJZXjQQdRMtfcmapvNZ/+xXlLW2cHeF0cZ17ua3LeyIX5goA+Acp0ryKJio0ZlZCjBn6j
ut01oRBQXl3SnAqXzVWHW4evI9h6aR6bG78uY5OjEBunDqGdWTxKjRKH2pCqRy8rblEnq3QSHSq/
iG2EXKf+jfNoJtavpydAmjK5bGpKnsEnxVRWSQRhJPLXEGW9O7YJjVhTXQYTQxoQqv2XdLbFSy14
+EK20e91vbwuThengUa0Euq7FnnOE9tnIFsZiZcKpDLT0u7Qh26BZWtgTaE4SP7yqATEnwXRQREc
UovGm5yU2Eoay0DqDkdYe3313OdFjScZPRAJikPLpiWezhRfGn/RhnEYygcccT+BtaX/BbilNv4g
6Qjs8107nipz4ePnX7lJK9Pd3S1kAYtQW/xlxzTSCfCseMP2M9clR+q3acDX/T+Fd8Y+LEM4qmlr
RKT9o3hW8jFBhMkPRq5UHv3z6WiFEhIflusO1O6woFXJiI8ioAllsc0M+TxNxKjmsQosMo0+Qta2
f1az4iZrgyq0LT9PwYB5/m+CndtGbou5ll5Mnm5sPFaQtc2obE2oNmfsowkRHvFbBUE0N93RV+E7
byvrWWq3QuMA4l71vGBvc35CcZjDWIB0jXZIV/UoCICgXdmWDDU8LLNkrYi1XivUBfLkEf6Ml5nG
+NHy/wYXVY0bs2y7uq7b3ZcopRY+jukHOGMzLeu7r6XT83PvqYqEjBROC61LKxT+9byMJ3ydgz2N
S4+BJYe7Uw3NWQxKhKSTJ65fqd7NAmz5YlvpARJzp5tJkJ0EP1LAQH5rey2qrjzIu+KYmHkVbn0Q
my3BtLx52DrvdcpWsMlTD69Ksp4D4pLX2/96zextlLl+X5LgKh22VpF2KuVIYx8tJJbWleXc0SAH
hDbFOL5Byg0OUw/lJn1f+1SCQj4IBnHQEk/+7HLp+gJYo8XysT0U+31eNDYeVClbr1kq1i+lzheJ
zH7NgrX3gddsNw0WVqMk8rm6k4qOyl9F1BF5mlLYT+0yV94ISrfLeHWkc46XgEeEsM4QyYWTrgOJ
wABQyrwUeuAbJwhykUaWjJg/1p/TqeRDLXDxAh6yitgJ9xR8qJ/EyWWwof84Kafyi1rQvSgcGYG7
n/Tcaw0WfKeEJsRRdJtOo2jf8kfNXq18Wg/ZxKO5dX9q6MVlyh5mG0ovpAXfny9WI66RJFqzfuYl
G0twZUdUrKQdiNxEVvfch5547oZdDXk+QmvYxCwFLhkKrlNCAIBC2XhFkshtCKt6qhN+tHIVA+YW
+2Op8FNlJH25BkZ8o+5pBkgkuUufVATz6kNf3cKe2vyoEs0PRTuXq//nLxxHm6zNTf7rhOJAvF4Q
hPcMVoy4tJqrXQdGBWr0lG5pJ3nacGEbk8xnP+/41BzKaBW5qsp4kywlQEkbbn/A+ZKuYP5O7K8u
ZW91XMlVHMus37N3N3MRpnW7kbAfvPSu9h4/p07Knmr4FvK76VovmuK5wJsK2FEsI1hgOtBOequj
RKnMR1c4EeQ/Uz7M6D7OvPqXBqYjeXRQJFzMGEzpEWV2Y5phFX645V/2IPLxLorR/SFIn/B1KJjz
z6L2lMG9VVREYXszC/oGlJzYU9zD2/u5hp7HMSfsk8mGQHjPiEgXI8VZ2ucCkSuiovgZg7zWGtB9
gfmhWbREGe7GTZmVnaEhNZ1P9yrBu8fjBldgRhZZVCKguF8YMTfS2u8/Qfr1ooh9J5PcrwjN9W1R
xLqT+mjnPHbswf9IbLtUon+Qb10AQR0w2BCMQWgn4u5+uUSw8CAtzAep6x3Vx3QCsXKPx4QyFSt3
pmRx4dKbVnJWUSwLLmpqN7pSFkvv5i1eHURwMtpctqIsvRkO+gtF/njUyHKAPsGb7vJN/vcAJcLH
Lx/2N148HmQYvSJ9PGTnIerKrDHNdAEMPiGb+PU8TftEemrmhQCuyq+k0KA6/IEFhSqNgDI774Fe
ICJFXYoWW6bAFV573jeRqeyBXkktcePihnDtbjKx9K8oRCmj9WfazkQF0U3FXSToS4iMqPN7Rh0Z
FKhywFSeVUySNG2rqRBzKOykiAQD2A+W8D65BkGWjH6G9wdzqKuERV9Y6dohWyIqujbRiF2BWSRL
Q7WKAmfZXIq0njIn+1vv+II3OV3c5PXzTFVqKChJWZkGeTzTIfVLgAJvgT1GKvE3AAkYNoc9xPPT
RUGFSEyVE8nD73YC+LrANBibJEfE4H5HWSRNv5yqv06/aRXtHlGOI6XPNnr7Etq1SpvKC3WxYJ6m
m4nhxc41qbtv1wXZl7O2RZh5Co4qIlsUqM4rBXAtAsgn7gqiPcalIfKKVu95eMP6tJpx1JrLU0LM
eDlYAKJ+XCTJpwdENjDXsbUpTEz7hvfsCwTWXVEb5WWcBC2Ab72jPTnuWSc50Z8SMGPcM/GypIOD
mJfgTcPweu/nDKN15zTurV+wRK4Zixu0pgCcuS6QlXqFNhkngGsxtObzS7xDu2JEGiK8Cx5Rg7LD
L0rme+VBnkYCZWLJixjrC+/K9nhejl/0aKZwb7mnUbminU1QGhUijGSJvduU3xykt99SFyxzfL0O
K+0D9Wnam39YWKDsTZ1Y6n5M7EEM9uWrHjYPfqHyCQ1XYfDGXlS/TsJrAv1jSolm8KPn9vgNjYcg
ZMWtmjOK0e8VIR7grqoRgY+HgUPPqnj4Ge+Cb6+3mTd4ziCrUFAIRFKA5wWXiaxXameR7IR/EWFM
CMWLSDR+dPaAaFIzpq2y1NgFP7ctTBJxwdrnBVB03g6WW1xQuir+Hgrr8IiSV8SrdmrqqvWl051r
k1twVHkd8f8XOYpKC4YyPcJ9bS4rjRlGhBFIFjsy13/P547CiS5JO5lHWh5dNLQnpoNCxmuZHtGR
HNvPHSAzs5YH1QX2SYhDnYN4yWGfI81gae73ERoQGpyZDg0jFfoyGI5BKWqI7ojLTGa9uQtQunoF
o9hydAlLyA6wWFQqrLSoXnIXPQfB09/bBhhMO32ykTA+Q0FejCSVFoN/mVNbssCiUFqoXbbrhthT
/LnElX1bZX/OM3bWuAzXyFn8Sk8BRO1axMJAm4w0OcPTpnt3C3xkxTCoiswnVtGJ8BbTNcPB4vlU
OHLRxGrf2Mqz7Ev90gkF8cjTdfx7txbQO27eDqjp9JPnj3AmblJAI0aXQcGuDRJhMsIlyNH1J7zM
qYqTlPIT2xzktVwk20frvTSm38xvmYL6I9iMVEdmJ/mQSl+VS/q96bi2OnKUZQevm+p/DjoZZSMv
l4lVIgfEg3ji7Is+QFxKRDQAdUL0OIGg7EU3wJk2hNgr5ro/9Gs+6QV+5TRdmj9q6EKfxGTs14Yd
6YJqlJg0gszlWlVzHjAjzMus0oUK9WwtZ04eXETySN0DUgbHqLDCV0ki2siLibERgoiivgs9sWTs
FAGxuadGAwUQrOlqaoCjTcGqX/SnjrjUVWjqBC20xpuYO4qG2d71CaQfP6kCwjwBbBTaxp5bMnva
kUfzyAiPgVDjCvB/0AOZ4Z5fDb2E+w909Ed0NcvDGwGQHO/XEj8VGL9bp7Hhtx/r+TYufEzBe/L/
QmyDfSNslr5vkusaWHl3RJV0BI7bofdryc5UrHTBLDBR1LegcgwJWFETsodc63VjI/EgpiIwmuZl
hikktXJolITvMCpqvFeyS/wUzhA1XbzkY/ColSxH5l6vM5+bC0OagHtD7MpFWXRGVJspPDDqMnLQ
aiCl0sGMtiyuS60Tn7P9g5lt1ld81eukj2ol/Kth4O2kU/XW8Xsh8WwnHz2nLN++3dRrlH3hrzH1
0A+D3mdUpRITQbv5a25IIxxBaa21rXjD8iSBw4j69jbQ81KeuMK8xkArq1JwizMUJMroTx6iPhNY
cqYXw/bJ4ZLOReTnJk2i+rz9/D1O+Ty8Wp3FrqQJqzUaDBMeRAT3wK/fDmHlkKkHSGrqWq+AsAdX
hMvx3TYP6FHbQDgVugFhybjzvLnDTU+itbU1ovAQyfnuqKGoHLwuOHeEFx8GAe34qo6k2Qqy1Ml/
GwyZ1Kb1lTwk7p35aow6De4eIG7Zl6uDnwyVGV7JyMQAqRd1sQPZGmChy1Lj/Xguu6Fpesk336I+
P/JeIISCyXqDXHvV3RUh4eYwA7R64t4NLI/8KFOwJ6UXn1eq/tKO8K5IKe2Fh48XtIQhvPOipgI5
jtP5crkqJ1PIkuZMi+hOuPq7MDoy8KxLwnuJz71qZrrKZtigWxETcjsVzM8rXcA50d9WRNdleb+O
Egzdf8//gP4ClXrXVNJ+LQvt8TVavlY9u5yPsGloXj6bJVq6gdvHKSCb10MMzc1vDbNi2NDNPPce
PT7S2cMIlk5MtvF3w08iV1jNdnwWH7tqFYJZoP5Qv8BxvgREnmweySKbz19cstYamTWqCe4upCTr
/8IX/M3mfBRwYpYOvwgsFDNcQ+UG/+7ha35ePECWnvYDQMXyEk8H/qqG+KTqf/+uoqfL/VMGdE3Q
A4WQmay7BMaPPNGnDHd0SHMbmJlSYchqvBaEWH731LqB3QgjpU8GG+iBl7ZGO3DujQvcF0EfKDk6
EzqksJt/HlOlYUYmfiA5759yQEqK7y3rX7lXDcyyVl71JegNvyPcRqYqP1CXBF7u8GozjlhWlUcN
cbBdQpbyQJRAhiMWWmayZzSiw04A50w3iQ237PERZ4uoCxna4elrTSm1q7CLjpyUVXiq69KLNuPI
pPjaBN54ZiFnXI8cPromTEl85BPZ/VXXrPLaEURFEsWcOrrPHgN7gPcdvKm9mZ/Fi8dBOUOT3EeD
L8EcsfGbwWneR4xKT1XOuuGk37GEjIUAU0/glNBCmy7mkoHLQ8w0Yq+Qmh9YWAQqd7VAD+OUq2sa
aU6kjjw0WE7n8XIxNZvHPVJ+hTRkTamhfxrnbMfh0YsVVIDbUsF4a5ry3fDz648AsePO+7VC9th3
Om/BgntEnhjvKMOzkTg5CKytTjdiS3rMKwod9VlqNEl8LqmatNNUwdQ3kYKgbNEMEWEFZrED58Ed
/KFiciBWiBQMj5MrWHukDef8tEu6h7ubk2mQc3ypxoEBqpp847roqZmO90+WizDfShLsY8fIA8Vn
kS2Rq0KcRmymon0ppCoS+IQnsZDe985LdtyAAcF86/3sL8wQQVNhm00QaCqmW0daAI7idO/jONpz
rHCG9N3OUrJ8cuEVMCqHkmqcTWuJUUm+2bmULjGMwycyidosUg+UiXX/IvmdBNwm1hsdVPm3Wzwr
JW4g1YEJSMNBCJGKNKY871YeuBqmumHhD7GnI1ijLVU9pb1uyB84oTWBVXLC4MFZprxXEzdhlBuT
f5T0uz1NiiR1TgnA4XvgFxZFK4w/OBATMH9Wnrwm5I/7/HQx6fzGYex3pI0dfs1BL/5sa0HST3cn
DA4EHyzJFhM+3deQHZ/Cum+1+DAtaCZcQGA1DcYgmBn4NMfulyT+9/GWuXJTX76lY77NC+CruEED
Y5vqEcbiq+AdHtkiZfrbBwjWWrAe2RN+9vjLagBz0MUI90JBQYqFMk1iep4Y5oHK2Gz3/W0Mmcjt
RODnkZFr8RrVi7ZrO7IEuyzZFgHa3ueIzj1EkZXfxXssX1rWAwc7BlDYsyWuh2dY5AAOt9X4hd7K
pR69V8xmqx3dW+UVIAUc6ndt5Z3SF0YqVDitY/Lr2L1IbhT3SfMOQni2g+Hm8esfwgGX3sd5nxO5
AWrd+lCkkHoBAc+EzggI3++AFXphWw72pdV+yqJx0yKYEE/1be87S5p0tdYXD3E5ILxUv2vc/r8e
BXql5/ZweF+aXPCCg4Z9gXYXpp4DBvksTaYlP5y3a4PG3/hpBf9KCQcOw0AS8npz5q0EJbMxpbIc
H75ZnwKS5xQQntVWoog6Ts1ZOpeqgpdIb0tBbcD9igK1LmA4a+4SpCzs4HELTR1CvraSFWmy+W0X
NgigUi+3fA9/9rtqGPZGpYVO2cq0jGf2HF28E5S8hLXxK0WvYhhNhCOtvLE/BvXwRHDCx7ruLXQI
2kF5hqAUUj+CuqiZ7gmpYRcy5KN0LYxRcpXJBxVlWFywTsA79EEXN3nr5ATU0CFe08ulwIV7n3fV
GDW6xRppPqvjiJ2v3/jAczn5dRq4IhxvtucXVQIWVx52eHT/vRBo1uF+C0Gu6dEYSHg301sXZ8Hm
btTtKJ+XVuMDWp9vkhvdsEaMBTbZyZFwRgwbNMEfT6Dyhaszx632n2teUvcZpAcKjcF09u1eENBz
JKn3fL74O7qRwVrONHSnlUsiWKND2BT3MBptjCZcQykkslQRy9Umd6tkcBtPUpKiEVrYPlruvhBy
0OA2cLjNXnSAzWSowhrpE/PfDla5ZVcspEpWSJ2IRCXqylGLezEPg1ChRRFMgMTm8xZTQBbnj6G1
iQiLY3qZBgaCoB56BYMtrn7a4Fqt3f5WFX7nNDufjgIe/x6Is19DF377Pc60H0W11E7eq1Myfroc
4dpc57AZc7CjIn5/E0NNlIuHdfvTrRm2fAyC1g2ATIFNSqFMlG979o9IUTMI5+ehWkB36R7hPxe5
MFoJrmC2JjajmWAIjwEcHpFh3vMXCiFhpcnO9O2qES2WD7/0+P1e5fN/6MqSWtDLGB5B2NU90h/o
AHQ8RqhvZp3uzSQ8Kq8+ovd5cY0eEqshIg6F9pF4VznatD2tnkjqgyvLs63TcyMxuSK5nA13Ndr1
L0ih+cXWVF4nuWQQM6Qy/O1BqJQz/Q7x5e0YfGUGsUhBOIyX1w/UWtshHsX7k9Z9fGRBSYOS7Clx
453WAg43WdzY1rncjWyZAz9MbXrsvIiW9y9WQrQcvFG375+lqp/H5ookqige3nRxXI62+qdpSUd7
OYyd2QfVoNPJkxdBbkaR+xgXdZNsX0k+WvOQOT26OkYtDW2PM+5Fj3+AwQ4Y46SERSKeW+YgmytU
99d/wLQNnN5+A5oBdcSQAskUTZ60ZlTY08qQFh74p9kahmr6fzXnqMGMK0R7NhKVtGc9Mvwh1KrL
u7akghhlmItHJZnL6boMuWh66FY9k1fkJITrEOuytRgCcKjOdiMO8eWYvkYUgBU8S2soMlAP+QIv
AnbzVkR86A6DTnEL0eeQGYdr4NT9tVWnx2myfCBjPK5JAgSa+Ow8P4C9yC+JjnTZjAoqYQEI3Q5a
1WWp5I1jRziWFGohvEwPb0FBv37AKkyATBXLaguZcFB4XKJo0UA6J8WfY4m0xvwHiMa92SsIvV+k
hM9ShVvIqwk2nxymgh69AlgZifpn8n6c2lKtUb6KuYNy2XtFMnlJmcOkz5pNiAtr6IhzvBtLyy3K
TtEV/PcirgzppF1HV2MnAUDuruGVqicBV5Lc6OB+JIiQPviNaIc9mpfXfd4/5WPb9MU9+PVB3bia
Ef2NKuvqz314D7staHTtaLN3cwB/cPh91fqWBYcaUpL+sQYq+HbMTNLRfX5+OrRUlYWEAEbWqBPH
Sjuv7ZIv3Hgt5mE1p9JTA0a3zAhbiNj+JpNaYCu7n9gFmIHYwy8/RVHNVkNQMPcg4LBMuAdzhlbp
Bw0N80+dhA9ReJquYcVu3aNSWb0VRxzTiPSfeolKkpec3iqa68W/+Rp3W3oSvjP80IDjkEH6h3MF
S1Y6aOuLGXigIgZ2wM+G+NuFSF2+naEmNbUnXl4Ua2FUpCUWxcvkgwoVzMACDoPqlAO8CAVqcRuG
P8Y/rmW/Aj5ARaTYrc2lCkUlB7LRnnbyFRa3kRlapM+rbdXV8pxo9tYLtc3XkPWbBLJjG5iE595i
Gg30kOdM+z5r92nfe0rGTnQJBpK0Uf+654c08jDvMvFL8DvyJ4fIGi3R2oVtrVPHWkikE1Vd4n4J
7YY3VQ2NJzzxFasFmzG5SmibMVCzTiXUFKEKcQUjL3NpSGFvev2ETxEkP4hKUZBehVt/IWtz50PM
+efydvs2qJcjQ0MKXoEKTjmuENhbqikUncWw+7Jrr/UjXI+sCFkurafs6jgIKL5+MWZbFHsHJPct
eSgATIuOJGW3uK8DxaA/nTkWJJI4FJL2N2bfY7F/N2jh85hl+enkkYKTyd8Aj59JwKZH+pxA5cpz
v+aBq6wekDkKOsunRAkiy2kowWhA0zlr7f/1ISIpKDNxuwoMQkut6Qbtqs7XYl2QhEd/3gcOvxmQ
aYtqVMvoj7UM9JuEVNbMwVQLSvz155cEJeRXtrsrs7Ph0NCKu8w9CgiT3VNuk3bgOpAP4c8u2Ld8
aI8+PTinDP0lvnrsEENdTeHDc0qdN305AG7305ku7deXV3/6dI/PTPuVR9TODee41e+NMltweD0q
qDlqYTWU6IcTHAjhZZvX4LrKhZdXmr8U59uy4+lmE4EkbQj8V7hmYtOruh54v5wGGVDlPfBfVnlX
lSoql6X/uezOP2g7xc5frtLAYVCh6ArV/h6W9VH1KpSq69wlt9YKCe9KJSjPMGTQyg8OGTk3Q8r6
oDGeXeCaRKFyxtd8rP9LPvzrV7lJwGabGsW5yTpdOoBARb/2JtwXofapLl84dbZa+GkXGVypdJA3
hW2DiUkAyfrw58lUjJeL1ivNKTP/GB9gCpPtNkvId3+0SteMgdQT4vhjPAnK1EUUAHCYlFziRxjj
PeSseiG3mNUQtlBMqwr+DJ4uPahWKC6DBZwtoJdE28ChPPGSJmDTm8KC3fjza01Le9ZIB5p8WNjm
2G77XQJ0jISVP3a9t4M2qjuppB3ssuUixJuxHGFn0JNpmfhscjQlMqTu7tFgezPzS4P6jLuBQahz
ZxWVIVkQ9ltFjcbjxdfeEOb9X4SE1Wq+mpUJTV/VjF7qTSEYfNVceGBu5aiPtU2/dmXPrIN/4Zzf
sZCFbo4Th7Ts6qjHC62vTZ0DNoGUVQOrnxrf/PWy1ErDXCw3VfeTniqLOaDhVxZY5rDBQF2mB3HJ
X5j3Wru3dAxIcjSBlhu+fs85A023LrNGNRvws9gt6cLcgNWriPOr8isBap5m3eRg0L3JSoeRQYH1
MIcLuFjMjJNUWUL7QGBC1+QOdahnwaD3s3Qyi6lZ25CTqD7WNIuB/Ilu8KoOLyiiyWZ1KqUjwswB
aASjPdezEGR+zGhDt6ldMbdUmbuQEYLHzFUP3ELaJ5sCVGMPL5mcE+hPPEAvOq0VdBscrznoXAua
EzgfXerqmIM/iP/XfjIJS09vfQrGweOxdBcvset4LKy4Hk863PHHxYKNiDssRz8jt1C/sriaNbYX
klUcBo1Nhxu22xayaTKnQVcydlR38FrprM/cSgNdni6tJ4hYBDGJSmvOD0lX3ba4hwuZVhHqqlK8
qv58aNTAWZ7DcGtfjio8YFmM7OgDNWkMEJRglAZ+m087A+jqwujxUgOmodSA+bGS7ybzQBX47gnp
fabqMANOIrZER1LDrS3V/RFnnCagCOKQMC4VbwZNk2u7xyKv1Gbcechp42r03/w7zbEJIKnDIZZk
X3md4iNgCZs18oDUEqTcO8vUyA4UKcEgLyqvX8gN95Emq5Buk9HDK9l7beORHCS0RSYFn19R/Y09
YRHfheWCyX2/28+tm3de18uATqBIQonIQaWLHfIrqww3E6UExAhdcsoDmYZgesHt6FCpgWEkhcCo
4QbVEJeb9ZQW6/X1zw5Emz1MV7SxQ3hrJ5nDZpk/zJBgtryQZpGS3e56/xJR8+X2ZV8/usxssRLh
1t3mdbi44uLfci+Km24RTE4CLI9wOeMsliCU7nAE4PGE3y/AhHUJWVfdYezQQUa+iWX8LC6zMpij
+GaTpeWDHwlD82YcMZyN4E/B2KBiqVp5WWeKu8f15MK41+qHrTs48gfHgds1+iNI04CTHs1WXY1Q
rvGhOp2Qzdwlr9XL5zhkVg1M0UHcnGawoWh8B5aLonwCn6hfC4H+RpxaNQkRNKZYD9Cp3JhcksR5
6+wZaxOZAyuU55IbOSszuHJhRyBU19zZnBLRozPfQIbUfI0cg1mvUE+hv/7NevWJbsJ/oL3OfWT9
oMJJiFNQdyckqWVBLObR4jvTy1hSUu852XgWoojvyBPtaUVpIR1S5StGXQuQ7BEcgROvqygtXkAl
GBr6qnDj7xwS8TDmQfUm0Y1T555I9LwvxtHQlgw/X7FLXM8aEjjJMnKzuY/6wrtxwTx9aTvgrmXh
1zQGpa2QfeEn+Rr4bYCvLSuOVV/gDux+sel/gOTs2X73V2QWt8zXZq2VjKYbEHzTZ3Tccnc60Q41
H4CIe+2jAFC7N6C2PtjFS520RpVj2H8DoZAVQ7j/5gYDIfbgWhJxpeMPL+ULp9Iu/Wy6EhXbfzSO
7p/R8lT5SP4bbpA2uB+dY3rQsrbSHYax8YWfSKiPxtWrrfhyYJZ+VuPoUbKPjetzN7HTFsFUi/eZ
ECASE2MkOFy3pjdSp8JpfWCAuYcvKuQBLoCFu8F9WOoloh3eD2IHskt8A+feFWmYjCilwVXIGokb
qp41CxaLMgRD2wjoQS4wz3HEY+/Axt6aM4vuf9ri7B+KrUJtxAScpzPLHvFhZBTPa8U9QcDSmS7W
AkQzUZEkgmudCOz5RsRX9Tekx6s2LXGVnuqEKS+s1G3qIgF5hoT5jy5VOkeOMyT0wgzLcnvb6aZF
jFpwxC2rKebPZ4wcCgN2gaUW/Ynrug6eokag9HULdEzqpuVRmursQonFx//P5P8QeW3f/yhBAZSm
nLLcnZapfmPf8lxMwzSw3U8sILweW1kXnlzGs1jN0YEZlQaicULqDktXZrTbZgpPAflEOGH4nOpm
4UMF8snfi2ebwDd3FPxdlgGqFtcIqyHpev+0+hZ3zYs1OO5fHb/RkR79k4yRDkXVVjrpSoT+4wsr
rpEW8v5VSlF8NG/VwWE2sjb/6/IP3zablc0SfBiD1NFMXE1n2Jgc57YmN6YdYB68najXzshQYMeU
eA6tzy4gfsvHHy1RLtiXP4wEsyt1zcxgAH5ejrEp3Up4yF/QDL7l/0ktY2VmRcvQOa9nBgWasKwF
bCZ23o5jxlEWwbTmCRF7P24V8brkCzq3PsFk5+vdtv5xtr3qMA1+KUoNXr2Zv7z6xhkJy40jxTZX
Yxk5aT4UxefPG5u/lVLOmz4cppK9rbMJecFyZFv0HdXhcpaJDcKGPwY8Bd02Ps+mWaHn+bjWaaHU
xbjtpNsvg7UqrLgPHphKMCgDf+zTSsGA0EgbGgR7a11DlAy4jNEDVB7UHVkr4k7cduKIOACdQU+q
KiDhdnZeEQMCEzYuODBre6C7kuFkspacmn1nhgAXdk2zfi9FqfbGUTGLigsECkNFv89iS5BMYt7P
WrULyi0/UrSQNNuOBEypKkyWy4TXgg3CzcRwIq+46sdYJzi090HU5TvzZLs/dLfLl3mUmK+kQFkX
IWLIXYi/CS6iQmKCHWqwKB55L+QY5bEK7dqEJ09sJuHsyACTukJvZYiOKao+kjMonzhvhCP7rR90
RIsVNW0sszAxU0vxbnkywbZZ3JlZBHMqp2yi6TCqHggglE2IGcItIK4w2cDqy751cJUNtFtHTL8A
rN/6kEfyICvI7ETs+MkYv9qSYxpuq/6OetPTa9h8XdpWmZLSnUGqlbELTSBIBEyyS0sMNHHupJoO
wkt3oBZIBUrHgTdJE2LEnQ147ftRbUom6j/Pnb50WrT0dJIvJURCO/JGGIKvdKFvW686FMz9SVhw
u2yr1V+FImt3B0TATbgiFFMWJfsN/reOSvp861JIVxYdfrp6CMIcqa/ZB0J9W3EDCJDvcQejV3R2
3+3/xwzrjIbW1wAfP9RmTV31gpgslxnpzJ48uXQr9676bKGKgYHA3cxuiCVdQNvsf3vmbtYJjXiY
qrGOKNyPNejXtzHdOYL9bgGeqCxw9zbVMyPZjCkQPFUvltfDaB4z5Qp2YWvxXFUt431JqqgDwn+e
+0q7b8GfwlcZQavJlYhrGOpTbBkJPQVTmm29rx0kVr/lR097dSTqpgoEeyihoqnRlOHXb5c35rYJ
adf9tepqVoLafATS+fC/v66er+wIFnR0gqO/oqDRQw8UAKV42gYPyq7tesR+ei2Z7fAGT8U5GTFP
VGjOtQBKEsgfgbUVw3uqmjxkygF2+n6JQF6BvzS8LMk6jOJ4TKY5qPd/0rtsf1bp2/iHLelkBI8q
nO4sVDdh81RR38LOCnI9AbKYZcu2xHVUTywX0heAQvuQmzLtjZ7cfCuAZYN5edH3RJ7P3hZ6A2+x
Inw9KYV+yBcTPe6alY+P4+YuwQTZxkJNowAglKSFiY98HOyDMrIxnTlM/bNO9lg8bimNVtzcb1o9
QnHtp/1VK96IcIEx8m1o9ED8JfqRFdKevSY/7yYkMRlT3xuMVuJGKq8hLKaPXxlmBajxR6KGVpR1
EH5XtgjOI/lhGxmhiJFDfTOQMRQuPKRVJN1cYaHRelGdll+ZITBe/rj9WmaNxBJYgunjr+hzK2hf
9CcOqzxeRiS6I3mHyQlIiDDN47oizBfKhRaVNhtQF2WrTpxhm2zJ5lPfk3cFB/sQdMTpFAHswh1z
ufzuRZqVFntKtcENUta1dZiKf4weXT0ByeInuEpkD6CseaGeYAfALxu1kO5aVhJ1lY4UCrAJX9nH
SjkazDZhTSZtZvcjv9lWH9PQiTsDtYzYsIv4e+nGRM1KFYZARZPYaakv5n7ROJHMAWoEW/yACal6
/vyOYaBD5WxWd0MuzsFJpZk0SO6hisCxNNZWSZ8+ii6HkQil8ufHIrKadhW++evl6axG1dv08qAL
FCuaD6lEyP4CY3VHgmgHtnTyq4tYmBIMDMohTk08ZjniiawBtVn/3F2FJKsYwRBBUaZ6Wuh7rLFd
ff6oLqNVW5xVz4utSEdOGrc88NUN3nDZvbk26S4MlEG8NGRgYap0uw6gxnmpCrc0N4TBWS2Xl+Su
D8yOjcQv66HEDin6unH2xApMBc5i1AGUAybYujk+11D5ixBQLMg4dmagahHStmn8fgxincs7N70T
2O48jR6xH+Mqh4l/9n+dXDQjnLnSx564tExGptpW0OH/WsPV0LL83X+EM0zLqY2IznwSoUdGHnZh
6KOva9F+xfEVO0GebdorPxDWEeTpueg3XFQAEME/G9/wMAtxuFAxLJPfqXfJnyhYZeHAutKMKpfY
wCOZtmgO3wpyqZYAG/uxRL6cuwZCYEIb6CC4ZVFvkGb224tMjAnmJwMV/mzp3D3PT7VwEuNCWcME
YWEEIo1iae09fllPZO6yxU9wJtKoR1quzdFz5Q8lNB0ezgTFBScUtj2/oNM5Iyk6WCcGe+aVzNqJ
CCKJmgyGznxGhmZV7qHzrsVEtq2luWNdQ703gX70mqr1ENZ+gIXdsh5eg+zkmfxwU8wC4OmB0gPP
tv1zZ6rNwCtjr1gXsVTkhJwSjQPYEg7wivbYTHVdHtMi1MsOa9h59i+lBGnnBz+JC9aHdyriHw+x
Ls0saGjtFSZrM8hmP+/yf4sc0Z/0tVwXIQ5u8xhcIRb8jENjNIURVA8cwRMO2xxPyOvIi8lyc8eN
7kYBDU5ABU5EwfD/3ceCMfLmtmN0Im2azOS6AVHXbt/8T4p4wSgyvZsx2Q9dX0GOImazn0n0WO/M
yxrGDI461k1lXvXpgxlP5Dxj9AGfwIKwOXKDmTmdgIJ3uhTfmWE4N+N3XZuAjsL6+Q7KqSZm0Cto
J1XC7pg4M9lL9lkZCwkIKMR0l/nJSP+PLDduD5jnvljbY9RUVd7W7xif89PO36u9EtI1O4aWFUZy
ZJ5lSjCfwvAma6wfR4PY3iqDoRczg3M+G70VagDqR8tqfdl7dk7gdT8ZPSDx7ZSpMq99juuAM09g
1kOWwDWpnbz6Yfv1UNAwFFvZPA3m+V93Q41rIC5E4A/hD6tkUFpOCErFfgQnNU0Er6J1PKHHHp85
h/fEZRVIm411+82dUTYpCOzBwojUdkofo+TzWCepCPMnua25dX87hu11pSKs1+W9MCe4PyxX62rN
q9MdxWN3CaH8AMzalWNXj8LfUc0EJHd6BjMXwY3AOkaFQdHO4dt2h1iM7sgstr1uHgYP6AZiaLcN
tUeqWpfKVadDTZXrTbqdFjVPp8SVGUwqgIHz9EOrpaVwcCW28W4Yp3oqXqlkjll3lBX3zlpq9gUJ
NZmXrMeG1pRs82R0kx3+OCnVRYuo3Nw5XezN80ES0Llm8Wde/DA9FoQsh100hmNtGpabHDqV30pP
30NR4w6ODMkH8NaymsZm/tiGNhZleLiKnpDrSbvR0dUvS1Th02VaGTABjKEUdgaeMHnQqf0qyPTf
gca7EIxeiFi/euBZxvZw1KwTI3dgEPa6YehUymCESUU7BoOF+iQBGQxj7GkU7gODr6BjcdcSf5vY
NYOkvgcFCo9JGscjCq6E8EIc/pN9/ScLnBzwbqqNtj9+N9a/qEp9OgoEvhtt5x5rBGl9Zkcha/iZ
yT4M4l6/0AQPXmnphz8N2pt0wm0qhU/S0Gx1q4D378dWjthUywMEJoU4rTCmlapxgvu4tWedYWzF
sts05AzyF66YBlrTZqoaLWoRpAdL1hgbC0mJVp5TLLHOXVWq96onOoFYMAZrWomgNb7rT1phQ2fH
2d45Ucak6hfOuo7ViSDiQP3hY8ypgWE+8wT2HJZXMbV+no12TDBNj2oH90mSmbBUEJ9kPKIjt2+n
6T3xoxIzGf1yUrx6gEKleQfagTKqnUuWlLzQgUxlQimpn4ZkzTdRYYEtpgNL7ixoRJEzEDcTPLfz
IiEPArWZJzS8TjiQxMqrwhr7IY+Mo+C93mSNU3i/+RZoroHyiahyoQHtI54sI12YasbS6xkgO8Ht
f4/GEXul5tan7NvR2fcPRgzA/WTy+gX80DbcGtOBuBvjxnVnV4QwSkBWOGPGfNcycvuid7kaX7do
wDkWdIAT4TstYBrOf531NbqsCbf5iJNlLvOuvQ6zr47V2d4sOsgBz2c809v/85qX5I89sLr/r6ab
6ukZyQbreZk8LC1mmXSXAOM5wCq9yMdtVKNq/Iqs0qK22H27TQ7iTCbZ1QjHkMQOF+odqrsIz7do
Yg+n1fMadTk9hbzVzFQZkCmgDYAy6tQtyFQuDYlcL5oAR94p+RkzKLBl6mcJYUZAvYMnLYwnPHzB
XBrrZhNkN6JV/YqMsFgJEGJ+IME4VEQ5v1apzCpwEdplP00PzcHSFys1u7pD+dNYEhrMset6nv17
2A8h0rDt1kTINBTFSoRH3Z+7/eMr6gAzZy3eTqWkNZ4oiDr5IfToOz5/hSU8TfwEa1D6RC8mSIKl
aAkemwxq6ipyxXd5r3XKcHwfKWOuve9NtBwXnorCSGqt65oJqZldsFkpCDFhvSSUZU0iOglql7eq
GSuf18EEKpLuIwrJ041mKtKKO4ZBogxz4tMPQrbPpg2/wPqtUuR6fTxE+bMm2EVVCiUw0C/SmLh2
SdUt2jFFgo8bi+yKkYgT/+iCv1efd9ra+zNruTyYGAIERvtb9EwbJGW0XvrpqkaLAE8m5ISIiSqg
YwoKpXznwqm8RqOJGxM8fptWe7VxC8dS+jiWlS2vCBZE8/PP84QMEODGweqivOOOZpPC6BpIoqFS
8YucyC1tc0337bU0CuY2SjY3LpYWevbNmNprhFAq1f1HRFKeEOjVNgaV20rzAhjCxLRsqQGUj/Za
KGRRHbSrWaM1dXOw/IeYxdCuBhUEq+/6moGftSwCmIFOhWQoNK9dsAWg3nxrXNWQyt/krBpsqIHF
gdmljLKqrZEKtncn+VbaYMSBcp0q76mRdvKFAk25NjoIj6SEo8HZiU437lUiv03MusIVYGHkB+n0
I7uoWbVLXfci1wrgwRNbgDS/h8QsZCptqxkhxyf4Tp3RDWptBmc8tHsR1qskhQLZ6cY80zxHGZCY
LeZ+OAyA6x4kN6my3LWtn9D1bV9XIq0CI5qwbADKb/Z77jxt/I9g+HIQLI7ZKjQoHVMuiwQjUK8/
+3H7RkTY4I/95krhlr1tvW6GEjvNgSrU1YIQ0r+czdEss5beBLQpK4BWJBZ3nTKik63nGbGD7XEJ
S5gxkKfysrSZil2iP84eatcChyolrcKrZ1Nio95tpTHoGyN/c4pl8ejPngpC+S9NAJIDYBjI9UyL
zhsxUsD6XoQEZi5gP/8xFasL+HPZY7XJaZZ43n0qOWcuzMw7+jvr1tfVSh0JHZukkeY2zhiuRvvB
5qdLk0FIkDgeM4r3aAaosMoQDc0ro2ksES1qBslEvpUibAyLiR0T4zHuxHa9P9R5WeLPmZAKK3k1
Lak/iKIlo5vB+naqEkxxA3iZYnLt7o3wNKEa+5glo2SDU46ndAKVyYDRUyQJF9vo7L5ole5xEfSl
ORq/MYPXgRawLK9bwjjozDo8skbmjcgNESCk6ZHKlJRUe3xV2ayQfYtSJUX3OvKxVnS7MT4y9/YX
k902AwuLiW1v+bm9dJtgAiyxR4cXRt72BIWFQIMM0EKNittBy5uC1s5D9VNrcboOZAkHJo2NwiuZ
i5dhACyRu7LG66spFx5cVAqV4DrMuomijDR3K6hSTp++SuBzENmuE9+8UGOshBoR4lGyiIp1G7+W
bd6WhipFqWjCM55NJ5DxBW1BpR4grHphRkUkErt4XhQeoi2zjjEP8oQG+MC8/pvVyI7yjkLmPvPc
3iXMhaWma0AujN+T1nYpWR3WmLTrQMZb4ddIdX7OEzej/q5L4ozgbsxl+mgrYZzZHliHDLX6Ddm/
rutEzFl/F/6jTdiCDlWgBKZdCgjqMrt5HOsxBn5nHO/UwUp1vWJnlzB8xqnTf//Y2w9/bWaLuprg
Y+sqf1iZ1Knu45UQvWNghTPq7mDquHi4oXs2IyEUOS0UNuxNyYWnaY9w5up1nmfrF8HpHqrRce96
j03J8m7fJ2aH49uDpj6DvvpK+z8csGhP5e6eZ24CnbJlWRYBZXfAjNS3BAbnX9S2FJQRdxrbUiLk
HgAzHXa7B3C1EaxBbVBYbN9JSmztSAacH8PmDNCqRJj+jkJm5pLJzIlrpWVF2ZkRLHpVUfSzUenz
Bg7mzTKVZrheXyNGB+hl3pkBQit8p/s73pDSyPvQ/ofbJt2jEBKrxY101kkLLZS6Q3RoYQse2HLs
WF8ktEU//RjksKc8DOZ8813rvmGYcCuX03RheIdiBu9od8iOxsv8CxuiVyW2m3oHYNISnj6zcduX
qY+KehZzaC+9QYkD0N9FLcT8C5jpAYHundaY34zixajNZj/4AwbhcwkDPOORg1OOTZF2+iCzlBjN
LzcefroKe3ylvdmcTdP37EfHwj99N2XPvNQ82eFO2LajQnR8qYnx2NoXmzRQ8OArSij1GT2q5dKM
5q2/oY6wArfrISzUBkI8mbV520jcnMuUKIbIKlLWMZmuBfXWY+C8kqpdLyUzn5ll1oHTwgWsN9e6
MV4XXh3xzWK8s0F2At4RAAfGR0X8EoQGRfCux3febmcaBig0CYMkbiRkaCxQl/mpQYpuF8JeMnxu
wKAtIVKLGucg0UIC8MaEbDmjYk+H0VUkRdixVln2sjhWCMuOjSat8b778SnkZaE1vW2xE70t6ySY
Rq7W7maJyxeleOYNcTcGYQRtIrB/GdCGSDdTVH5ZDSfqagYAZGGV2JSx11GWZ4SaIrGkml/L7P2O
sUrfUe8gZH+Kv0tp3Afag/y4ZqPGe00VMIKCJdajaIsxwSQcc+5AdZ1Rfrvmc5AIhqimMqdd2IoJ
lO/HR4DXW+x4wCGf9qN3k3sIXzhdngV5VoVlwBAvdIw0RUqCdbZ/tvpt8NmIDnD7dRk+/QAWUxNp
nbJO049a5mfhVrnUcujRWoM/jce5b2zbRWPM941ep7LjjluRrwHZbcjDI8LzfX+HGUa9rjplH8iB
WF/i4iregwalrqCntZZryegMhjz+5ndmrdA9XUiJ7r+pdUOC3l+e7QxuHqUCk2Tdo4RbIDyojeKc
djJ1F1/UEaHSLC9xttl55gNaux5M2aWNHhLXIWckYXK47jL6XR6n//piqE7PfsJvK2Ip+dWM5fEp
IAk4Ks1c6ItBeVlOR4DtBDi7p+6qqQcsZadYuvzNbt0DlLEtJccE6R3XRnqsq80zMxtw818c3W+S
CK9/Fgn9Imm+j2Fhp7IH4/s9PnKUl1RXQgM4ZtsZTk3GKOTgGl/7ufIoUZqt0vF/hE8jax4+nNxU
PVOwnimIz80OHIswl032o43tB//BTNl+D3KjhHPL6IqHLFuxMUkIE73dqMSYJHpm4O+g7mU+4s/I
Y9+jjK1OXWQCmcP+mjsgSO5OSLtQJLCb6dg9SVIdtqj5fwh9NAopsLlFZUxExNH4UbTsfC7cX7CI
3Y1VvUw5E8131pj2+ysSkbQrJXVmdHK7/D91TNOs2Dey1eslYB9rQF+HueIbpQzaFTL5z8GrqKMC
t/E+LEADxx0CWZi+8BWc0VpwOfHgjYBsgTevHDMB6i/UDARKbZ1EdMYFD/tAJcPZgaC4ayP5yxme
wmPH06rosJo+PB36Ih95HcsucbgJzmsY1Zbua9LEP6blwPWAXwyeUntMhr1x4/T8b5oWeXnts0e6
jXJr6/Obhl7OIfbD2X8eb7rpc24fDBKmZ3DQKjNk4M+/37TUy7ssIjXm+aRkOd6fkDnAoy5Z7NSn
nBWBtvM0EcuAiPOLx2A+aKiMh4BQgUR+R0+AAx+rhgNbHVrLgSw1MG+S+4WP4oWUT3tMxpz6HBkr
YAx2GmiT71CkboGhsv8+03QP8IsA9Nz93+yEiKei3xS9K3vOe3xiaIxEhjRqGFCZrZ/0cutdKc+5
C31pEaaAsvkaN+Oo0Vzdmmm9BrEVNk5u2N8L7YTUi3VgvzLMYL9+95cyCqOZligRQQBqW9iSV3CN
yuKqShC9MMFHSvK8TY63cH0pK0PvYx/gR/4MNv8rpnZoyku6B0JJ7Jem5eFbm3IdTKzo1ySbXkqP
ZYXFn9ZrxMGgI2XiPEV0KJfQK7d8vTlcOLTU/ykgenx7bszLqZA2YjhzIV/5yJFd+FxKDQGAqaBl
rHCeWPUMeTMrPdelSkH2N/DYQlwYkLwD1/CXSSH70CSJA6rAxS5ZLBfuQ1BrEtRMNv1vJ5gLxOkx
xGR8Fbbf7Cc5zEt6mhqhRFz+VfrmBsJ1hMlnBgMyn6FWZlVxhQ+8F/bTtSn870SmKENidxuFvm80
/ed7hGb2JwIX32qBA1o5HpEH+WZfDww/ys8awBI5z4HH42wbuXTzHpESulwR/y4/mbkcKRaGCtd8
nerTiGyi8ZmF5mp8Xv1WpFDdBeleG2Q+xO0SXhdxB4+PPovosu97ArAX8/bCIjPhKno3KGE1Zvbt
zdddQRqi850/slQP2XW449AZgQNDOIDSF50H98zQaYVdKyCAFCeZS16vhJYl5sCS+EeqqwizimBU
WdNbUM9MtgCY+MmV3rgC9dwud0/nvWlhjQDsiNGW7oYiNTZ9TV0ZD8J35BJKKARijg/bNwNCai0R
+OUhNCm2C5nVrQ6uR4s6tF2IRGrmj8c3jBYSa9G3NiKu9YARgYuqnGkm2WLvYm9USEPT9q3Fq4EX
AlRfsBgqEtOSV2hvcTfyNjGfVkP+1WBWK6E/MVkL4/X63Mtfsh5kmLFSfSNetCuwvOk+bdf/j13d
N79IQIh5EniH/exaT44C18F2uYeRp598bkQBQGSQdljB3Iy7k6+enOme7orCOXP9stZtUC06Mq19
zudHMdmJBBI8SiHsJn7SRo05embEouamxM3sboln/YQjpBCYzaGklJ0MXvtAEG7/XTkerq0eJOxe
XLrYQ+0hBV9Sgu8swP+9JJx7jXl/8tpCQgXaxtld7VzHUHWnpOTYpZevSAJTXTbdYdRH0FjGZtiF
dO4u190hLpgPAxlD+NnqiyThOkMkjLqk5CLLHlTS9+UJxtoU14iF0bBe4HiREHkLwOFiPs3e6g3g
mlm6qClBLTNkrxrBDs6kW/jKhosDGWw/XKCue+duYudahgN3zJ8PFx+VYgc+hKxbDhxiPVmvTJHD
a1a+5ksebk4YYzUexiykDU4sc/XR0YA5ATq9STOx0rZM7SfRD3hvfBpCesooqWRfFIfdp8A/LANA
0GZmx4OyaE3swAE60/CeRzWvOZN0ta2JCnKzZr8Cymq966vJaV1wdlggqp5gSNRztyzzIpR1MCXH
sZv23nGxR8fHCjAN8IcBul+ywgHPE/miP2ncEBr3V4b06euKN7i8wQF/BKyppSdm7BDESHiaPyL6
QV+c+4mabxVFIC9basa84ekjdXssFT/373Cx4ife82mYQeQfUJhsuljVYw6BT4D8EshVxSy9xc6D
wkg0M+x56Lq1bVIGalvzF+YSB7JYhmTDLRX7jQOHklV9yarEPaNByePQaRhjr8e9pbQphi89IQva
C5fISRDfJ8n0YNaqzObwY4zyqzmYbFb3Hvadj8mpJYul66mgLXqHRHRLDWPvHr2wt62Ps4QBqxD0
fvvR95iSklgqftAM8tTOL4o+UoH9LRKcEKFeOQfD408a68/ybGrZEnvmyd4dIwSez60Dp+gB/pS7
/MaMqnHdrrcZ4sZr8Rw2PX8fNPUGquqpBTVG+6GjXihyyCamBdUQNeBAduMGwjgfO58Sic3UXyhS
F7ByQIP0Vr1IkW1qE0bA5JAF+0MCADlh2fqY3iywSI13KMIPQgQU/Nx4lugmOHGRKCI2k33jOwol
1iyZbFGWVGoGubm+gVJklU/I0shz/0UIGjhrREUOTaX6ZmVITxMfvfU/i4zYbLlgAX4ZizDg8oMW
nEBgfQwbLRXMS/mQ+HfthuGRDVxPwLWEpc0bYeVCI0qH+io7Su1bGUaumXP+wnnjsttKSTS3xL7L
p/vIXIxKkAKEA7iaRvVawsHLX7xXQvbsSX+HXfMMG0X0z98SpYjB6NOWWhur9e5VWZSoNK7wsmbq
4t+EYV7gZH9pknEtWFvbRi5igabZPn1QZUP23Ozfwo8FPwrGs2EYKOVvTZsvkhIcqQE82Xz/AtRQ
+WKlco44L44lT3kYCYKs0wSb8tXHY9CuCAQw6/dIGnw+2H72oL5SrGCIWqqIybmZhDxL+IWnhwIp
H/yTBmmf8kSGDM2G96gbFRQtclj0QFsc9pjTHT9pqLZiSWS/Wu9tsEpqmpnaPRdJzIA+JPfzts3E
U/OpGaCBfas8md/eGJH0Nvy8NgQAbftjqfnjJt/5D9DtK296KNFHmcVKOeTGXTzxcYaa/vsWrud5
ac5eZ+1+578geBwhVOyBtQwya+3Zi65x+Wl+b1GsfM6mpeGKUwp8jvVzFquD1I6iMdBPscdUJghH
gF/ZuCFRtyGpZFyl8hD4Bs6eEzzGFUOSYepYtwzdD7BlxAyxyyjLFJjwQSL2GzH56dIsAuytr8In
89KP7BdDvwc3LDzODa4UqT+2+RLPqDXV0tJHD33FdGI+ySM/H1MB5bpkGdsZUp7hzPDctNPm0crc
0U1xkyk40CeOWzxzkqSHK2rjXzW3eeHuvkD6I4me7WnZUmI1fNqMBlGBoSETwkOmkMs97bMLOQwO
26HD7GIBHJ9tdyeoP1od5npnljhvt/xjPKmMDgxHhbKvbhgaWccgifE6ij7YcMNy4Ayy90LHfkk+
OVXdRxHpHudY3dB4D3KcLjq36X8PxzSY6pY4MlmbpBpSDBzEQiSbDo3dRWtkdxd5gzkAuYlcoDSx
RwSGF3gm0KVo+upuzFpieGV1Vj5TBnWSGTTBzRqMAPM2Omj6ENCJuULaV7OyMe5GyjzJU1gPW2vM
fm1bORTdtmgDKdSQ+cE7Urgmq9rJaW5O6uaW8nsX68BfGeRe6iTEUG6nKpMY9yDvkaw3cKQdmbGs
+xGbBoj9KHBsGHXDW6XEHSjB9UDhW+nrNRRoG3CIv8kp7ydAsTcdmWjFCIBw9s73zrhuuWfPe/6Z
BOmarsuozY0LpucouEtIh8+P4xRmuMDhRDHVg+npcMBbaU75jp2Zc93IZA0oLrJZ8sV3TK8B7OT7
cUvop5Y0+AwVtGOoTYIxNds7Ws8gYho0f633smSaA7/bu0yuQiyGX4lJpvkapNIq5A65TdXAkgha
h+aAB+HZkW9rZ04kkqzQ6HUH/xEP/liIX6fyi7xVVBo6Bsw2DjmQe/fku7ZOVVrmeAA1fLWfdY2F
Um1et0RBi/VnPgAdHQZa88JzlAZDFbAiHPIbmu0Y3QWOv7C4jH3lYE9v1EBs/JeB5dqrLJ+TKxbQ
9wAdZzZSxmhbarR9KPc4tVpp4CS89SHJyhIfx1p9gdBBn8m40dZHj1Khki/9V3kZaQW54DDb34PH
Fl02/qG5MiU/xsQTD1nNzUgTP/3/ctZ1Zij5JZ93ONqsuYUgdraHczukleA65Et8Dvj1p3Z5YtCD
jn1r4tM331qBjy4XxyUcQGSS8XV3m4PpmmOx78yBQv+re5ivbIhBAiV44+WulLt0cRS+HdlHy5yp
rAZrqEeyX9kDEkkkbaWaGCEPcL064hmv1NK1rVieq13YBHDgs8n70dMcBHXZvraLLfoWL61/5ZkU
EtShqRV6g6zStCJp+Qx1x5KO7s44H+kAWeoYpWHc8zYSzTMDtAOglt7JFsf9s8DrhYoEmHwFhaxx
5vP/n2UsG/91F1WTfxGKwQTFNtVxgPBWyh4O2HqYeMzz39u0qQHA13pHLIQA2jIjZq59AL40y/K+
wP6yh6B+IEPwFqPmb+CjQTRnDebuDM5zqHighs+V3ipbKhcFYjbBC2gZd6k0YoSrFTqalVEZqSKp
iwk5ICWXpnWr+ZqcoBZ0EBwy1vu64Zw8wu9Yv3MpXxAunzflGCcP/6RZJDNnYmJB+qOOvZvGIbf8
P0R/22ktjbHWF6Qwcg4GLwcMmsuBfSrjgu1W1XrZ4XHCFJk97Q6tqXxdNfbccc0+FWqIs+w+AZdZ
hdSdmNzQx1FXxtPXCyNflV6CXHo1qzMjC8QUl0pX3kfYSCQigLuX2ZIV4ij1OQGszTAA9NYR80jJ
o1jONiNXCfJK0nUjFJAz0XxmSzGCTohJ+wXOamKQktP72h0vtBayOy6eXPD6CXuSHY3dE8eE05Ol
10bZXQM2DtvygMEqHIL4tngvN0yfSGPbW6CGTgcYe7UUWXEisDHydGUnb8lcC0qYDl4or81b3WCt
PQniOfgUI3LMpvzL/ICwpfnRRw6mNIHoTvSXFKzvTZaiivHKTjTVdo/4isByX/OlXTFUN2ug5JIT
fIqedSId/0GBKGCzzaCJLu0EfCGv06ev4QsBoV1Ea4XX932Y9f4Y9tm5dUacSppjiEleIc26C42N
QFN+U6k4t5iCNLNOW+CLPyaD+p5p7JKQmlJ4eQrZiOJdeqYbOSX96RdD8IGcsY2/Zy5YMlNga+kj
jvWNIyQi8DmTdS2LjLhkOE+MEQvHkScQaHxhCqV3lNvdeXP2eWxFzjupNxLdzHyltXLBe2SebibA
tfZNb0q/KMdh1kYoYc6QcnPOsOoB/Y/FU/pC108XDT3Hwp+/Loaj/h4G750wzeZ8tgF0ygT4tk9i
vqTn1fk2jmOLI99sCAEJj8gz+ufVJH+qfygdWVKRBi2WlGdEDzQZ2ndw51lGQSbE2oBHKCDHtDLe
BWGWgDT7GvOmmBAnZLvtAzQctrWAruysCAesuC06tsykcMGmBzBipsp+CuePrL71PoCeoI9pdV26
kJK0OPLyhbSkA2yqjHDASGsKqRORbcwaDh/F/MNYbxiNznAtm/SVaXyIOWRMYLq9Jg4pCv1L9bMO
21UrIwo7QKq4GqiJonA04MStjrxYcMH7nA25wuKzmGfQmyuH5Cfx6IEOYaK1fpgkdYslsOcSCxec
OYMfb4JhSuSWj1yADQpJAcZyy6pl3/u3N1GJ5P3mm6TGAqpo9dEgzULknIW+S5cgihBllJY2lDrk
WqbWFsdXVGIjmDvcVQpohKXywslHbDfuCbHvuMiA7fYtGfo6FZQOPcRkDs2K0Dv/IO5H4PbD8swR
AtOmT1hIPz/5LpDn9IH4u5ig3DaFkNpaiosj8hq89v7im5kZmJ01w4ccmR2ZGemWZUWdsH3MicT0
xE2HKjEhRmw1exJ5pKk4hI2QI4EyLxHwlWPwLXDiCuk4V9hFE6NmuHB6gxTxWGKk6OLc/ggJlJUD
3uNYCI60KbN9V0gz9OMhEbqZWHJVcinHt/2/nGh+2Y3Yv5sk17oEKB/jSJazHQaPtZRbljJE8DPD
CkaVnlyY7PvSOs2d0ycXyu7k1GENNCrcSc1xHBCrR/9wp3JIMrPRf+QrFuXinh5XLaveFI2hXlFP
RaguoxTjPAsKGd4z0+osN5TzfJ2DKb/8bTgJ0v8oNPSovdCVVB7mByKXgySmzIZUc9ZR3ANo8M9g
pAKmLqNv6tpDdHNqWt2UKfICqKLF6vEGoBUnu66i5xaJFKSohM/DzwtLwgHmxBKUxv30K15bbPJZ
4t+S51mkhVrw/fgz1MSX+U6aJyH5/DJyTZvgFq0m0Kh+n4GXeZtodsfcnUSBZTz2bXr+BbEVFamm
MOLhaosRabT1MHeXeDJl0wnc4XbfnYLo7ZA5HJfqnodh4wyxMMBHrXC3qJ3XFvpFEldGKvOdBtpW
U/ij1MgewPnaiLiOgiNb1KnpSbcFJFPJEOj7aetb2rqhjnEFjma1OT2yDZZQmO1+lFmhslcrSHiZ
Nux+A1XLpUCR2ZLAqQAcYiKefIgenTJPFhogc5bg5zaqdUn9bHdzmlwsza4UDH879TTjETQG91A2
y4HJw9kT/6M8Z+S7u2/XknrCJkTae2PizAGIsGa3dTSb1bgv4GeQD1rxHKifGl8UOBNeHDk/RI9g
L7I001YnklqBXsu9AOmLLKsu1uCqIg62Dlm9tP77kDy+MgL6WgHl/JBjDwTdlpjmHXG3mA6xmebf
wsKiFq1SiinTy4myfqJx78ZYY6xug1SQKdixreYBWzudpKMy11l6rYKEFbbsMfeaLw3bpVm3fOPA
Nmnc3qLSGu7LCbV+dsMmS5yb+9DMqM/P/pg/bJbCrKdpIDObekZMpPFeHH2wz/7GeW4x2B0pnoAZ
VzzpV27cJrPfYb1iMBUqBHCcGz+zJi5vwzkWXDFLZX6mwfk0f4Z+vK60Ys366qpJWHg21cH4E9HG
yK0KJ9me53yoWJM9AUgc3VSYPnLdw/U8nRF6hfg8MsAbPuyBsNoU3SjS+VkT+gExd6eKWcuarlOU
UsCwFQy3L7pEU8riB0xTpw60M5A70ExWZORcFw3aaX7UEUxBT6hYFasXWpmKXEW3pweGOLSkoTmp
dHoFH0X89+f+hI1EXIbK4dLMZHcdMYDWM5L5exZ6fFO63NG6ulDuW2gLADqcoEFam79AgaOdEkwN
MIizRRVT4c2EuxIXjP4Frta+S3J71BgWCHC/uopF8K//sJt98HZZdD9cgXtQVqn1cVJQGfOVzEW+
XWFspMNcQNADR0j93IZVZZ9bxoJS0sAjw/SAD0BQrykMouKdwQoXiSS3krKRoUHqm4LZCytfk6RB
nb1/zhJ2f3YKFZScFhvFgDmRPYU1PdtVj9sJ2yN9OgTXpr1UytRG6mBN+io9O4kEP6X75ueDWzVB
NCjKoek/WJb+Xh015eHwJtOHan729Y/305kgsKar6fc8JOimUaYa89tix1OuebfcqEUG1C8NSwfA
IoIoxpf2f36zXbUWalz4+kFW7o7DoLzd4p2QtuC4SMr2JI379IidR8R/5Ga05lh6UwpbCKV6PjI8
Vl8gtb63gpXpsenkIBW+iY5D0ugRT25q0oUQLAcN93UvvLMg/WGKTzT6xYFYxQAvApWKdAekskM8
nqHmUeiDGyg/S7OkMfgxUYVGyiuy+UpIP7ICXaCIFl1JKF7hFPC86Rmkj8Q1CVoDwk+IcpKnHLnF
Jj+Yyi4Fx4GDCWnNxrTjBPRXVB0LW+yBL1oQyX96UGeOOj9OInV0c8Fx3vlsNQZSgu/mRzxspTgO
rIauzCw9EiwHEZlPLeraIbiBtlaXwyB0ME3YRy5Qi5ywccf6bHC7hlDmpUKliwuywCd+wwp+F5FW
qpc+Joe+LiGyHsuohmnGrU5PbhuCnZhm4nOowF2a/blp8x6TJsGl/Uj05ap5nLJrVd9siKfEOoDj
U30/JlhHYHOMr11BWAtSdWi18XS7VGi5HwB3JihDnE+0UHcRqhdIuxU731Q6wTHx+vADqrjB2eBQ
GT/dFuPiMCQAD13W7dWxoS+W9BKH/tBLetoqEUrUZu3R9VkOpNiCRxNSEP3t0gqYmjgrTlWbAubK
8cETseseQsOsWE/dGBj6S9ANlsW7XhBmCmns+pTFn7+MXwS5ZktcfEbM1Z2dHHIqu5CNNa2cMI76
kG/KNJEQAhWwcvTenNx9elyeQTw8JoW46Z4Fqr0qCmZEO1etqaUcBEMsBkLl7CiAG4uKAcO9HiEU
zmeDCjsgyYCw/99Pw/V0JTueAa1vdcg45eTEjYK6Mqim7WNe3S4rp1z1cMQKNVGEw6jRiENTvR88
36dFOgfjEdZLFF3i5HxB/9ufJfdcUVvzWimlTTg0vteJ5h7DZd3KN6v/1ik/4E6wKBPKolCfroMj
d1PuvCOVGewat2RcsGBx2VZUcXd8tFOWYo+/Twb0G7n4uFS+smdW7KeMqW4z9vevKpaRWZeZUA9S
P+0tW/8E6LnWnc1bjFp4Zt790P3pF7sAiC4hZZhTAVP+VVejBJvIBpn4xGe5gtvnIoQyV5FvH6uj
Unl56WupGRSt70QsrJdyuQQE8uiNmsCl4H4bJuo2AZCEjcPBydMahNg2OWFE5c2KWkcjtF23mg7Y
DD1TC+KqrWKiwKLgFQNHBMuMGm4C4ENFooZxpXritJvNeRes5V4T7mOuKfKzmDRYad0zOGhgn54Y
sQDIlneHjtJd5Gax6vw31+AwRICI15rY7CHhSYX329IZd7gpxk/aaFqwDqLR+uHRd17z6eFfvA37
41ZI1/DhPp2Kd9z3lrje9a9uzcqQ+6kauiaBjcmviBmQZ0ez/51Ak3+m/BZlPG0M/jGSZh/InxpO
rD5hWnX4XCTFZjW/xSKkro8nruThyeyBAxRdhVuf2k2EBpNkVeCxm4KvqN/6oAxO4TtR4/wNc4sD
wuvdsAEE2YrDf6XD/aQbjdP4h85av8RI6X1xZKW7SYsxGNLx30jNLOoCbtPzQSwnokeKhmWC1ZWF
+7TY3Sz8LZywUgjkUkAPbp4QGP402VF6U6xmrejHI+vwW8I7DkWTiruwtF0T1tnouYK4RMfoVn6L
10DJB2s+QtmvJ+lPjV57GbwotlisqKgzlXtlJPs2vhbqPlLWrsWJq3r9OeDjRTSuShz2Fg0cCr6f
O2NR4zo5j/lCAW5C7vAOADSsmnaWsCBCzoUDvdHgKYvTHccDp1TEaOqRuG2+7khtmtGS2czVlsOf
n+eU+w++aZ7VYemZqaEDM93mbudzIWMjwryie12i8z0KEeAdSHxf+RX1gobyKxhQrTor63jN9u6J
vOp7JXDBhQygAfE86VQI54Q612uq5zBbLi8Wp7iHKoEaFtA4qGYkUL0mfDfIeHyu84JB67BIVc1Z
SF04j4hXitmNRibYbXpFN1gL2XnS14M1SDq7e+T1fylIoW5UVfARZ2HtiW+svRzeOwk7GzQqgOjJ
CG0ERrQDDyB5sKuJ42edoYrYjJPNT5pHHuSvt/dC1ULc7de6rtrEHKKskHt+AbMsQO8Z/nGT82d+
zrWaL+G/pI7a+fqRI/5TAsS9vjhC/CchId+fey+cjyIj8cqTgpHkqldtnk41K/AMLmjYGfEcWzjW
QPKNb4SCiZwNDro6www4i0AnlwgPRxWilz3/rOLTzsuRGtl4wTrMBpxXQTfzV1QUjHgxZFXoXVpW
letLXJV6UPd5xIWeonwRpL8CpJYgZitkZtSxc04bDhniqpY0PJxw5GczXUk5qVszsjMq8zhrGfC2
04bBQbxUA1yo7KEX7k3+WubN11FWnjaqFIbDEMOCXPKdjpcuKAHVSnv5fFeDoggf6pIpa/3vB6aB
5Rw0Ux/3LkwRP/OHLhJSderqX7Es4l+by3f8ni1KUTp9i/t3LmZ0z1NQNfAzzTvL9XzVFgR3eKp5
KhlMLf7RxUjuVDolPjTZpfH8JL6ltPtt3GUch8STruxqrYyc3tdxwYvodwr2zP3/RKENMKK4Oyc+
bz/lz7LqVKqQW8pAHSiHrdoBeQ9i0rmHWXamLtUtkUivkrZ+6QhFNlXmKJbX8pzRNPrY5Eco7Oma
j89w/CjBKHR712hkgUo9EB5WwCBusLSpYx4NqzLB8PtX5awEMSuKq+M2f5dJeOON4SKPEkjs/17T
8GNNXTaAoTrTONRIXjeO5EbZKVtEj9FbbdaEZioHkQBgEQxldn1eCdKUgfV7eRTI8kyHKvQ0Oj/T
EZUWW2kFPAFEmkXcgcv5p9EVewnyWxuQgDOXeAEnWnBG02DOOhKWOnM+Fl49RCPzi5weOuY6WcV9
gHbY4hSpG+NT1R+0TqXslF3EoEx8sfdqiyWkR3gtFz1cdnItLYBdBQmQnYOb/EfK4USj0AnmAHlC
KLnE5Z9Mt19tH8Dbzs6MV5I5uObszVzNKItjDduS5y0brIqcnZn2ZzXG89oU5sZZb0V7b5SvH/sz
JGTvmhd1LYoAZs1gJBEvDlphU9vlLpG9hGnWsyfbootOzsroduQboRb67/ZYQxIXWvh4xRbamPjr
PHCcZeg/XeNSb005nKcoWwUfzS/hheZSuE4+tkt2DpKkVLDLugvSg4u5eqY/hNEyPNdOwj6t+mIv
50frZt7Gxxnxbkea9ysgjEZFcV3L+1sGyoAiRYYkHU1DVcGN7DEoBoWTo6x8ROddOT7GA0Gt19lY
6Yakq6g0uJRSJp0MBAV+X0fozq0zyLgOnlnCHIEumhKL3MkR9dhNRaYA/5KSt8IGNVQH74jZ/EfD
y8OytplSIcyEp7BdhUajc1gzeaDuxaIfIJ0Qg9MgQBMPCHl3frBAYsmWeyuxqvpA1L+s8AkTUCMt
8sWU0yqbDuLBur/O4K7XwWKEvKDLevb4xLzjH3kfMn7eEjKj99Psf8IrPNKtKGHpySk5gm6oureu
eZXkuGYOl3ua8CAzLKgxkCZtGBXBMVNV+MlXyDQ32CMc8+mqr6ut3t0eZTAeoXJwH3CT7lLTmFEz
PFuE7jZgRb/p0T62OWQjIbHQPyv+TykNAMyQuAz/Rsd2guWsqD9cOR5Nx5CZHHkXyNOUsRxPnd5F
lojGXTo7MHJWT9LUqhErcRE6UeM+Jot2yAwgWGMQvXcKITuv/u9VtyZrk1w7sKLkBtOsvA9HnCAr
6wj3uLDd3Mx9WXdmMBsE5N3Ri+TlBKHWrzWQIiVowYQzSHC4a4x+xKgKj8rUgyQcxedf0DoHokmx
O7+27gWFPeoTkhKZdaMg1EpMenma5JC7Ke8gXFNnvj6OP66l+AillnGt+TNLX0+ZgF0tFbLLmDC9
dCH93bPvBn6DzhH3wqz/D7xcRoFlqpI0yiPDHXyIZrwZD4rRqEhKkbfcXerbVXKj93y6f5Pw8ue4
zKr67ij9iT17Mhb/AqJ9jYJ+4E01VbcbdIfLG5b5+02CRsVG8gcWwzqz2Mr38RaKFFOcl1vTx10X
VJ9Q2cndt26F2t39uJevcIfPJ0fTapYoG6OZSdoqStnoTS8OsizKAQ1U+zy06JjtDBkNBqFGHpBz
gFBWFXDp65EoM/FO1SnAlU9qjFdVgJqZz9PCN8oL7xr/WhNoYuGXfHY8a4jCyNEGNSL01iiQGABj
kGaibBRrenPecdPWSqZAnayVuGNQNbpfwtuGIhH0ixH0fJc/LVs7cbWDKv9JVDBbAteKmWMUs1Ba
R9C2jLfMqG7X/Oq42TKAyxT+dRhd8mdhnRh34+Ff5AA7hOpOEdsbI6UzqgIh1O49OPbw7xTzJ5UU
nEcYrIQsQN29gLwMZJoHoGvUlHOEtbyhBypW3cCy8Yqp5QZKndwjgfx4L8Tr0tYtVDw7fw/ZioLl
oKtRr2zIuD2s7wMGBriAEuc4HigwWpCxsJ+99qkW8Qi2tQSRDUUp8Yr3wvuUF/4lw6BaRBSQQsWo
NamMfNSo+3XOx1REXEcDuMpaopYzJKTbmT7dtSr/tRWcdEkwN6pC34jT6MvI2UFYeE3nqBZ89xGH
CkLHwIf4LwgcPEVi66hTXhzsZERyrg6niO2eQ8Fua8T9ULgpDfJDDmD0ijgQuMKmyLHwPmj0fKpw
xxCAVlsdD/pNTkilFQFQP6MU1oBgJ/KpP3E6zVh0VpmTsRXaGddCNV0lIfQ/8e7D0sFWf/52s3lz
eHVp5XUwMPipocmmAIKIZkkjAlplPJsbhp3aECcVgSbIbtOqbg9p+TNr+KdPjTmsxQLOgorc0MyK
ohVw/FtToZbY8iQZQbLjrPPGL3u6YNJOoIkCq5UXsFZqKdT9jUewavMX5oWdFFIgJWxVV616cWux
gAWGy4vTSdPN++GpxdmGFnR0TnCggElVHyyApmEn3UdQ0pFr37ifwWpvhMJeRYKEyPO5Vnm1GJ1M
p6ljqVC8q59cQnpnVL6JE37J9bYoa8yf+WwZ/P3cW9NWgXfwqygjixNMn9EedmoRVRcb/H1MIteY
9u4GUz9nXRaOctFvXHDlxidocPNRjn9Xo5eacfwtlhsyErvLHiS5nf1MJF828ZJYqGjUMl/pubjT
4Y+oPa3h/ph50nSjkPWS8EtDJF00ArtpaSS55lRCWyz58ZO7fCMHLWkvJ/sAq1ZJPcw1SXWaETsx
3qEryVzQoWEhK2rblnj4Vk0XimV7erlbss1WWJVnHyTf4hvSUhWZDplOCBYfuRxOBv3cJp3zfAEV
ttSOK9kqCTWX9DUTXrO6NNosMCegyDr1C8D3zeZ0j1XDx8B7BQOrZzQ9N+n4S97fwaBWTwH2stoB
frAt5yChqD4mvUWtk7D12VyAgdIJa4ewubLY9u5hxoGDL7gT2XJHegNSbN/nxjy2QfdtwRrtUh7i
zPD8/kEWDSIwnZOatIoO4SsdPYi8WupnYM7SOfxNJmZZy6923e2swFXi0ao9Jw13OwibVV8wME0j
TRMRpmeXOh/007WmmSXiV6nb7p3z+bUz4rq3PVHVaoCrCEvhtdodkGP5FuEWcv20Cas68NxKxFnj
wjIKnBrT0m/hZr+OFotCcEAZMNh86pZQ0sRY+GXssKjfO93idDcVI7QhNHTIb02jJSlu82pMqLuR
ZEXOESzrWJ+v/SbfiI3t21HAt9DfFZN1jkMuRb9m6ur/7XjBDu0krFE/2nAMUNmdIvdAM0wAVVnn
8X5iNnQcZu5I1fIm2htVeEzKNj+hdFjq/b2kjIj4Tjxnejt7oTrKNPT4UmUFecmxiMx7890ZaNHe
gyp06xu7VBGZGH98PFA10NKf4WxiQgTSBpZ40T2blSzPm4JFWYBWTLOOmCpRs8c6H3fgWn+MFZ6T
Sc3/TDaEr/pCfEDdlZn88DAniGKzsTr8yb2zUdtjFQH6FljvPxlV0/nrUuHX2cj+kGQVrQlxd0YC
BNF0Ot4dcV2CH6KMXZz2NT4ZCoQc+hz8UrwIQkEDrY+xooRlEb2pZUa+TL7vr9IvX+8ntM6qzfNb
KQ89Fox6b/n2y3v0p6wTLqgEBP6xRjvBNdT4NYFOjUWz1tlh8zKjQKmXlAaRwc/Z2Xku3oTDlpt3
POnekcxwXnVEp+Yj2asCrcEgvIpqulCEJH458aYplDHrIeGHYslZ/M6r0LsHEv1WUPOpc6USxx2Z
dvzo++EALWW0H6bI3xMPy7vnZC1b+BIX9uKDFwa/kd/npNxs3r0tS7MdA0PTAJIRxkG96vlPN0by
U0LZgdUYZliepQBJsmpjtL4zOt466r6aEOwlQtwqIRVNpBy+8TkgOQUMRAAnjUf4aAfFTCiX2rex
kyurTPuWBrM4yytrLDConANQpOQTUXHXihwiBr7pNHNloayZn/ncqMZtGfXGJk1j20KafQ5zbX67
o6nLmCPAopSr2wB+DNzagr7d7Sbc8TasifNOyuoFbaXV+nF6Mad21DEn3YpOD8v3V7DrBkN3Jdf3
40EwdWrzdRAf6zynrGTZeIvhf8KC5BteCT4OVeIIlKa7VTTrjW/fcFuoYKCnsfQmlqzJqPYsrE6k
xGc9nHRr49PG8CujgP/2/thVqNkiaHu3Pk2NT1mnkZubBZhyxrWXJJnhITy4NMYthT9+1yWNnWm0
sXNG884nC/yLDC3NSfMu0/H+9yfdobVjA+h29zqC03M7DOgqQ0/cHkqjDUQEHba/2oBwnPzu2/5F
IJocWPFAUI78fw+7bKXIysaHS6juMKuDGyS11o3cJ2qAMcchFP0a3YcwyiX6yydb3FCS7jzpxhXP
L2jNxCXN5n3FrTPWZh1kJNkCt2MEE9nan3NHNYKDt1yAazSomX9LE7XvgTMIfzJCBfhRR+zwDYQB
X+u9xO+kh3BkeCS8dSttA1wxTYxNWksfl3uqjow77Y9ilwpTLEDGlONHdXwVpNGow151r2TXlpM+
HDYACYaLRXPuFoBAEozxOJjRo1mZreZrMb3IojoUxAQ0mk+gS8cAkF3IScbXBTSLaksIISiBsPuH
9oaSQ94ED4ldaky2ecmBY7eG9VZhoEpx0s67leL4P5Cdkt+zPwid2py9rg7JNyPu5MDqBzS+JS4W
AKoB0vKXVnsBDJchNtFvN50iqM/wF1TdY8dcMLHH2pJnBv998pYzm5Mw/vYZwhVCr5YQ8z+IxXu0
GI6bnhuFqpM/5Co9Z9OtpTqd03r4FD4VwbOU/wO0CVh0uAEyOg/c3DN0nvjluGJkenDRxDBSirQ+
WevFlkwdus3dRYcnE5nDcY/8ae8DNHBCoXvxIZV9A9DQAE81qu4ceHJbVOBsGNaPhWQISY6jynpb
lB5GgtKKBe0mtbFtuHaU8n9CnqX5TFzSQJux32QJUfnb/ttaUM2UGGgY8F7VOdI/P9F9tPTUiJ/+
v+RYEKDbZax45sYZkGE4tq4CIt1EnTU9VXlkoN54mjswLwekMfsD4tRRHSSrNZybdUG/Dhnulwgb
HnfzlwKgobwfRlRc7H+cn3S8gP/d8UyDgrSsQt/WnmONYUtAQo01SFP0Gq3QWyvF/9aza/usgISu
J4EWfxzc8ZgsaLXCHhKlMPYsvidcs2a9wqPDD11r5Hm5+NN4ZjQwTYb8zdBIFvZsHo5nbs2bmT7d
cqyVQpYxXN4jGHpx0IiC4Nub3WMeWdXQVmjcma1js1nIsOs2JgnRJ5E55YvThuV2YofxWpWu2+18
XGtWo2GIty5WNLvTl00pf549zE3TAWAeCiycyPc00cLkXwG9Z0AdhcfuhlB+UaWne0ZDZ887K6GM
1hKocWpiGkd9FX50xROZd+1bU0Xx1o6fmKNbCUgjzU/2Fabi6sskggefjp6xl5NPeDc+r4CS6zrR
2Ps4SgyUmakYfLQuJshoZzCIxvleEb973B6KJeG07I9AjtUgslW5fP2evIbeyHQtXwAJdeG94rGV
l+V1ezwUggVK5aVbi51il05ZLcaxb1HHWEzPmGJodCL+kUrw/F/FdSk7KdKzEExlH8pIapQ2cPUo
erWZfxWPujRpFSjiMpvrT7rLSv2Nwkj+O1qgU6PfR5orok2zneUrAe4ED3TCbrShaWq1VR7ILPSO
6+4+G7/FYAO+BXeu69azeuNIiezUE00qsA2QUF2LugIfo4tjPV6R+XAP+ABTg1lWFxrYoQnetL82
ydovSX5egUpxHCf8SbBRZsRG0GQiIyChTk2Wj9CNeGm6EvQN82WWXcWPVb+ltkVyZMPDmq06ISDK
iIZhTDRzXXn5e25Lhs9Xm4Qz5TRMB4ffjO29H4L+qJatllwh6WK63awk4tLyzlxRTTZNIriarkJg
S9O7Eyp2aWNpd5iusnQS0KQK4A2XcNEwUrdJNdSkutUeMPG9Tdq795AQI+aZUrO2p12VuXqdTxY+
u5JGXgm4QypCd4wIUqzCmW75r/KIomsm0XyDrg9JDx4YdrvfFt3GCBzGezXZtAJ49thMlUy+hrDJ
nJQSlQoEylHVb68JCCrx24ptGSDXYmUpVuphfle0KZiC6uk93QXK12fhIToomRiuwAI1pDFh5eBW
RMU4CQofKsQT2XRhUCP2Cw/Qs3s5FxaU2luh9dgtTXVTRog586MR0T8+NdaM9WRFUzBGoVpGF/BC
8Nam+RgGN7EDLQQhoD0bHjxvKRmmSOXxleGzq4rI/5yDuwh/1pSbMUfPdGcwnAWcRj5WKsTz/LnC
GY9GYdHMTnYlVOw7WTbnze0ct0fkwmy5McMBQvrJrKmrKRF5zqR8+eEueWCea7yn0i9hfbuijXiA
fFazwhAIGsvJEW4kGKemSc4IgUz1iw4g9c+NOWtdNuUDTvkKMqhZBdXN3ePy1XtxRy4ZrTZmkYTl
T5Ulna04/Mfv0dawoDpWv6kc2ZVH9M9JJA+5TdQYHLjjjLCk5rxaNjTe8YMFzJlNR8gPA+DmsHu2
U22KmNybvkl0FMEn4WCBxneSFgWXutzai/ZtEkid9iSWuwb/a84ROH4fF9Cr0Al/BXT+Lccgd0y7
/raU7rOm50ZcR8WeKs6mU5VIrKTJNWQAfi5CHyIcHEzJ6ToQXIUjKl+j88dQDnlARzVHNX98Yk94
7bgccNiunnjmJnaicIvHNd8Z9VHUMqxTx/iku8tJ6hg3dleaEYWTnI04v4ughrYDGOe1SuhrHkl6
x7WV5JizWMAPTLlQ9Anh+pQpl8gex7PJVOrh+q2rRNMlEN7Yeo78EvCsVBVHrSQ4mh+pnoW4kTNr
oLLdagHa2tfsnCvhy1wLWHN8C7ztLIBRGlsvS6XtRRs5VH9SFIyA9p8ZANCG80akBAHuVxdk33VO
ot2kBLVpVzeX9RJn8+awkua0D0cL9wcBKjJ/fMLstFqYjOXmWZ/Tcng92RdvqahCY+l8B7NGuB65
zL/zBMV8QCwW297U/37ep2xft+36K1L35fba+Yi+xe6PB4yp7KFpJPIyWr5nRpcT4D1K5Z4bJ9tk
FeLabf8DngrU8Xg/gbYX4UnDDUcA/zat0gak9GTZ1Aimdd//6vNwOxnTq9/cJlmX/N89lqu7oxlj
UQ7xlhhWoyvS1p4KVqweFihgtIy47V3T4rnZ/sYndO31ErJLEnP0x5hMlXjZKdvM89Dp7MHqDCKP
Yimk2LrtC79cZMpODgELQpLbv541Ua/6QxoO95IFpu13xOW84fFlygYYzQz6KGtgP9lOAYVRdCPH
aAfikPIy21keQMOSCIklc31wUIVPt/e4tib5juxxKdqM8s/BrCLKYALdkr4mljS4zeUWpqNLtO/e
zBOq6Yp62siJxxmz269M0s7fUgCzKmlXK56BEEa8NcB72AZRsJIH1Eo7Fb9Vofb64Fh6psLNBQ+A
SHgZ8wjWcL1oCGmt5oGA6/VAbzIJNqXin0On7FSm5boC44JsGH+sJt5bjnm3m7RJCkVyaiEDbwHO
eYBuwFM0MEG4iTrYIYFh3VYussKg/49RHPYPFummFdS1OuzOuh+vrkxqjcS/EDJASDZXi+A4Jb6y
XhKV15o06r3RnbwknInLi4jOSEkWaKaOPS6/NfYSfCndsLdS2BmSanAbzdyH3wiJCLbbJMHSHCj5
tInmpf7vbffK/wVnz6Am6T4JamM5Jui0n4i13QG+XILsH3hzBAOhxcsi+qyKexhxJnnLI5DvEKrk
IDR/CPwFYbQAub/e88VgQwJbzVAZEc94y/hn6QV/nVwxwE8e4FGm1PUjGAF+QopLqyUEotvlXcE1
JB8IEuYDbnqEz4tKcrLcHn+9MGnD7ilWHDgihZ0r83VSuBLvvWxLzgAPjTURCfxd98/gmag5S0tP
E/SI73Byf0xIPDcCsr8sCYfsIkGatKEJdq3aRT3gqwbLH6xrSD/vV7UO4QG+ftGODcPCP6oo9q0U
ghQ9tuWJSpff1o1ZKGzLdp+8IOUcRA6V0kkUjUwm7HJdlHL+rA1QZNgmJNXifi+Y4EyGAEXQ7iwh
/v4rQ6NnAyRoHpDtN4sUBBhgzAbsmdgfPtLe7IShEggmRMkjI91G98hZYpeHqQshJOfDmGrqmCae
3dFkwsc6qTmmvC0XMeRvHT5vRPTX2K8XecktOGEjl81fvmoleboQkAPTAla8qyHKKWtc6P24fofP
1wPZSpv0P0EUkEhGHjw7YQC8eH/7yt5v7IbiYIHc6ayzbTm8JeQ/eRk/DdHGlf8H722ObO2s4JR9
8lAPRJz+7Hyj2hYhU9bxQDCYG93ZjaJwlUJ+ns6kXziWLhprTSh1LP6qC3/ewqR7Gjb5UvBKBRt4
y/7/HvXicepB95QAKcSebQrErvLGZK+TPpIGkP8IfSAs8DkWyPmmdNWcwQ0Rtz2kyAJdMGa4vWf0
0MH9goMdwWOjH3Qo8jb3Lwugg6U8pLdVV1huzyfFasIEP5m2wmQU5oXb9F6ia6hBfH2KWu4jhhJW
XGf++JlGD+dAtvLdlrLtoDgGkVJSHTKO6AFjDbDS53QdPWce/OHl7f2+79DuIKA4H423mFvBCTj6
WnBioc8WYT4qdIjrGAV0LME9J/hCcWBArbNVcLQgKOY0aTeuyTT7C3CM1qqFdfuuJopZG77C0cXo
gFw8pmS8JUiqhKz4nur9PdRpcM1KWri72iyKYQ2/wLpVM8YNMDqEpCpWiREi95q0o5D67kzIrj/q
H+L9ymbSKuab249rq/OPVuN68dbRPbBlbGEaGzyLQYJZ5q5EON5fNVHHacEoHZAcVUz6cg/KUxQv
+8tbUfbtFlNzhhas1XffSu0ljLixAYSd1HpTJxXMk1rY6nb2ggPjUOI/9lBVe7U6IUU4eWdVYDKO
m7XRMKombAAZ9IDKzRP0eChEs3JIVlcOL6Y9BUP0843zVrPHefYAT89jTK+iRZ/pdHMlPQXQc4fk
AYU7zRkzHHO0bLfaIm9rRRDd5Eoq1aCY3pLor8cBBvOYv2/23gRwGk2wS0nDBNnlqp870pIuOZmE
ABeWkjetGmAlsJ2U9dT09YYlzPYnAzbiZqyljJ1oBza76Nve9HD9j3paWL/Wj9vgRw3mmRRowIeT
Cb1evGGbTC13sz/lYGnB5rXzYGArBD311V9OMeewFhBSZ+5bkts8RIB1496helnf46Sw6qgAHwmE
PsvUUPF85SDowyMKvWNiKzX7aRHSoeUFJLpkT/W5AU4psiiDCYVmLXLTRVOvtA8n++3K4uOI/AqG
spV3lF9cgCITNb8AreeGxOIb1WRcgugviiz3J71xKdWLkN1m4Cci7fJ2PwyA8u51TtvGS+6Z3k25
EWCAli7/MHmj/7Zrg1FxAYx/Pd+bF4SXDO2yFZxDwxRrrLBmvdxaNHJZ+UXJuVJGgH3JNwb0AzQg
wY5BxHAxjnapRaqG4fnoxtJ+auzJrMtaPtCIsddfzK/f4dk50g1puKbBKRMV0sblwpoMaGD6H6rX
X66SzG+rmkzqRSL3Hlcc496a9lRMA0xFvZSIRDrIFhhydYaRGG7b6rdNi8h9xKmQ6EPDsPGl04eP
qQgFs2Qw6zZV9b79vZz88u22rAXgkdU1K92f3JEBFZmn/vmNKA3GNZHGUjZQh2/Wx/wVXZUkONIy
KQ2FL8GFPSWHezeAlb4B1gTkUqN2MQ0WvFwAreLUdWeU416cIJn/PX4Jrx5GozVk5zskqHZ4XpaK
tksX/vieh8lgq5Fn7zJed36EcSUsPl/LaOpuGoYK8KqL0thqoWVkK/tUShEuEaeO0uaAcR/GJ5D+
4x5a6FAO4UyKmEGh74fW62dKnT2ENPX+kjItm/1bBu5W3LGv8ibfbeXM+MiPZ9X/EIxSsKM4VcsU
wyN9j1fWF+FJaiSqYA6Ksm8Zgj3I1jmfFnQCM8Wljw04TvscMZUU/SUZ5kZcY+yusMLaY0m7kB/o
4uk2SvC7Mu+qLOPn0HDBw8VZJ8xwifke8jp6oTJDU0qSk1+e9OMWvO5tZ3exo7XFhW6qrFDbArjT
y3AyhNTwp5xZbQ2Fia03CDlo9MdHpNsbrc9FEqwvNd/Jz+wgWIF/mI61hknvfZlXlwPzx/0aiZGe
IVgFVKpDSS58YUnjTcWomPN028xbZv7jwl0v9ClUDI4vUh218pSrAGLgE33y0R8bzG4/Bqmq7s3K
DvwveN6mJXgQ8y2uT3qd+Etk671NudgH7fsAreUzNGe4co2+zQ45kg9DCgvlsboARnrWcWMwGhb8
QElNpd5vsIpDmfSLop+Rp7ICA6kv/cLvgfyyyjUJdrrxawWwfG0P26v0flHHMgsOcuMh5gnBFF78
Etezhe3Plj5fQlQNtYC5POOKZvHbZloB1Fy/p1fsdMA7KQciLAssKni6EbDRqOcw+pM8tlW3N45G
ldQMx2Su24QL/4xFnGcEs0i12N1YUnF8htFTpsoKcLhRGPpBKQnKhDC7Fa5S5nDjKTZVTspDlWSR
JChmif5XgmbnCz0DphbG6ziVlt8o+d/UwnJeb3bGMKPxGEBxb8tElh5czsKicBI40+eFP1mlDCTA
24potbBb7yhqbWhU0ZnBh0t8Bj03Yz80hQF/gAMmA7XojLOSGr3gUAmrNJgSi/lYW+qMze+kFQ3G
KA/lCaV1a/xUBV2DB5NecuqevUczWRfxQ/6UnAJaIUr3TdJu0VUS5PC94xL4VUJ0ibsf56vTvll0
voMvWIgMgBI7DcM9Jux0AiCv05sP/7ircOUHMuLEFl2JXRWbaBNLayyu681X01G4qK5FkGv5ZVd7
MynhiemSXc76YOZHk3G9T4MVdEkZInkgIi1h2qJB+aUUL2b0gJfAcoNZTktr1inYtonGJEqrQeGK
kM0jKISZ36mI6yLAYvrm0hb9Xk9sbT1k8BckzSkJGpSdDMN3Q5CQYYMc918CnUPxvx6vhVphdXop
hPNiTnGnHxslxAR+8h5ECzjrSAKuqOlrxX9rMticnUMmw6o7/1CFPFeAtjkOxY65LbiZizTSvya4
19549WVtJ5RBI07VA4sgBFM01ffzQMNSgC/cUL20Ckp2W6qTBpPKOSrnjV2lsDNt5731IA/iPvI5
uOkkeLIRPdRW1jSkhvxRWtO6ugvaAxwpk2MZaKWi4ROnxCJ3nGIwStN7RJFFmqy+YqXlpQb9HooK
hfZAQ2RLAbSCEpNm1q7d88CJOBkVDEywUNjmYDiwX3ZU8UpMH7JQ6geEeUMbkbkNoBlkCBdOW0Db
Wgs7zjGQP4BnjlWT7/vyni3O2/p2FPVtxZn2vboP2kDOyzirXmRtxrK5qcZgYpFWTx4PI6DxYt5H
fh4cle/wlb5iJr/QEcOvKTu3cZJPYPfSvW9i/WBB8tGYu/NRr9jAI/FaetwJI3m80dKnvmgDOr70
cVK+dw47JPVk07cRRzklrDerBK/dcFbUis1E4yUSf6/BdUrYevGSlttlcLAMzFVNuPol+h663BkU
KSAdFC8ffrW3y9xlRaHecKTOoWpuHNrVIE0OEJays6K9018gBBDgFh8Lj7ijGf9FWHephMIO99VL
CTgiBGT5mFIl6AwmEhsIZYs2Q5Zq9DlwJ82lmnCXIVVXmnmL3AaQPdcSw9pld3cTQaMc4uX3NnvQ
GF3rDnbSlBTbjtTu8+i5Qx+ot/mr2WjVMrpVrc3OVTrQ3nW7sRJ2GK+BXhZntWIvBAe8bj/wJx7m
NjAPUS7n80ku3fDTeVwuzsNDEVs49Ny3z8cQpQ7R4vBbVFEKshKvuy3fmMgCoKAFs8r8mjEgaiy7
YDXYStbMkr3191IPOyCz/XVSSFodNqWKgk/SA7o5Elmw9gVVzCxLXOGtHkrAqPNXvKEwcQFJl/cp
EHogfxxlG6pmSnk/7u6j+6t5gBfoVXygbN+DvEIrhO3MiqMnFsaMuTPMbYpeuBy67Knew4HuK40P
Kpnmy3PUnOJB45UpHKK5OXDrp1qG30f6iWbze+5ea0akXv+RGU0MBMZzA3C0M29AMOZgbrDycPV/
EP2j3MPU1fRQQ4BYuYAged88oXFqqP6FRPKx7BbmcAijBV9Si7jPWYFb3i258fiJ8jktNe5OuQow
e56xCYVbikE0cjiskF3k3pe28FEGahcUXTonJZZMLxIrHe/PXHJCRCTKbG79NPOcC7aYjA6jvDuI
ocKz66ekxJXtTZdVqw30fG1ahBWa3UoX+mqqcM4G7p2oI2ydNow5X/+L68i3nnLKW0/tdi4Xr3BE
yODGrCfGuoQHNpez7+QBhh2UVr83A0oSyndgp3sorsPqzCHwlh40oUSblS+9XvfaNx2tiW+IVbiI
k2bmIiBiPDbs14BtVdaBELat9dZTM86fFWAzjG7uXGf+7VdIBbwDQ93JBQyqPlDu8cGX7IvFA/lH
vIJhOSRV6E+7SNgv47Hqbr5Vuzr/kzW+fQ5cb0p+V30aetLzTPrzHBtaInF9u39y7waYd4dK49sk
DmuHG8SlblcPtoFeiFBg1DfkvFqboiPGmFQLF3cCgry1YxAIumC2R9wvDTXusFWd7MIBuzG5E8WW
K+MWGKfxtvfR30JADzEOjD7GGHbRp+UQyaXi/I0fQpagRdz5rDF+nNyDumy8/zWhK1FlAP4pbuVE
q2iW7YXywjxrFoaVvORpW2EzO1pG1ssWEBrXuESUp2eAyN4d5Gd4s4BOD536Po93tjeGbcQGUhzC
MSBsipw8o04y0ZT4zRQK/GoJobX9Vc92KPKzeLTdjClL9/MPFyKT0AJWbLVZB5YioVxqHsOF+2Di
U/FGE54aPK+UikOb4Q4HJREPv7ELrBUI5wWQQTqKMbjveXbHhYLa/W4UoOfVuSa7UIlJPd5a1ayt
7azT1G/Cc5g1lyyGVLhj6gbNlgSoLEfClhYRD0DWhVI61trpE0CnUeRkuixE5nQ7rhu1B6vwtmkD
QJfzHaaO+kOv8ZgvroisqxYmbUME9iP2yRyPHy5p479WJvMQFvRfPFZcxVhqK2QWCSbYiq90JYfq
QaZNpkE6hAoEoccNtNHgs5TB0lvJV6e3bQhvjM81X4tMT7angCPVGCiziQKuL9JrjjTfSO8xyySd
uLKERf5odCdwuRFSlrmdX0zTpzzpy1EmTI/xyO+5SNXlIfZS83BX7Z3sjJqgRw92/P69TxLyKHgZ
uSa9uAkkLGr8nM5T0461edj9aWhuPq55IXj+d+cfxfNOHddHpeJvBInLoy3NF4W0WJMh3+kh30mf
BZKzRPj/9D60+wMfiUCAP7cu5bgNFQ7Y5qYy+MKFKk8wmb6B40SfVYFRtWR7jobJ4Q8QA3Qo8IZl
qRrv8N3RNL8U7k/cf72CH53zMiY4CA1tRDLkZBsyZq9hZh4WX4NmyXfuPnBLDu8p/xPgvACMdhnk
vCCWxAIN5gaTD6q/RG+k6NrFO/6BMklqavE6jVwzya2rlnzY5FcRFmu3H/xteV/fxpXOOP17rwh7
n62GTOLMfeFSe4nXzLi4WtAW/a4NfQO05ly6WWMPoBnq6zOQ2OwLOXGQXlZQ9vmooxY3oIGHrgDL
EPATvxSqoyGtwSteXsTmN8zfrhxnKbxQfTtHfeFm9XsAknLVoQMCrPlFA0zU2hE4JqRrNLuNOTQH
fxRSTqNl1BAE7jXOE/e5c/I+idYdC3VC2pNeLed3HS01e+CSxeFR2s3vZofzzQH7lPqYCYNNcJ7z
vnd0Bw4ipX/HwYY+YdvOMQaOy6jKvCb486uTfdnmjZAgl2Y9PeP46vl+pdL7GCoDzyd/m4ihOwtI
1S3INEbeKGDdfHaV/96izLl+VOyNPuNknpOdgU/5GIin9w5xD+yNrWXYvLI9I24pux15FlQTj5EA
794FK+npRjbXxRkM/47E66cfPwHO4z6yge2/1zvszIApAFkcV/9WGLinGo8vKprwL7+wYC3YOlxI
AL2c84l5L6JFfSkf23uzEjy01+CJL17HHD4x+0atcuBj6VQg5yFIqMhpvg+MCfKz2Opk7ueSx+nW
Gk/xnOMB2esFwV0kPV39wCi9MECbx+CWmz5bQU2Hmw/GojlXRYA4krKNYEjj2Dje/eiEYgxJsl++
00y/LUAbC733ZTzVhfOVSKplolE8DsQshl5DLFpsf1vrglmnhZ2z2lZPtE0VSAwioN3aP+F8JGLy
IiInGdmp/X/SCzPUapvrieBOXv64Zp2eEVSuTSZU9n9+QnbHTM/AxQbjojA2f7mMCPXpYgnfkSI2
XM3c7cZaV+4gWXA/SnUbVbAyGzGQhX35zhXCBRg3+qRBKKJg1DE4d5DJUT0MK8MAcvxcrAKQfIzM
GviGwY5HWnRgTHaeuBKbuU8VBdP7TemHVY/34KvYnxR/PS01g/2PjCa4yEe8quX3qqKX+nJrXJIi
BfRHiA69/RALU1x2d2IEyjdno2gvpmC+YklbES98FslCYJI1BrHsCq5ZmyTRAGq95W8n5yfnRb7e
QP0801p8XKc/itlWFmHV/vDNDeJ0ne84QQE3l2JhJxcjwR7/eGpxR7LrVna3O99WIX9Gy8+EJ246
TDAFn+90GP3m2WzfI2uRxmBKUSNUjOmtgeFc8rrTiSSGNUZk5i0o5in/cfFxtoTwgu+wJqTMrqQ5
bVBUvGXUUpFLyNCs6TPUA/pVy0Pmxhevw57inrh/z7KYMYeMLHHBH5DFFW90oqrN1pP/x9H1Sp2T
a2jekfYgYjfVbyecj2cobuxJfosn0Ufy7LIgl6rxgzFXksaxn/jL4WjCZqrP5XnXbCDJ29hwCeoW
vfe+CkfbJE0cO2HC3FTXeHbWPL7Vu1xjH5P2u2DNLPkVHeq120hdyz6IHa7Biq1/C9+IRyV3l64d
VI78wo+YGpGQ/0uIPto0Sh7fCAee3mdE2ktNDMliEpCxMtg+xXBrCfaUG/TwgmtXmB4cj4KQEjBz
5W/J9Oh2wDkNaWUWmv7768KZ7XyDHaWmZlfFtW1MjLY1WmnVZl9kCOcxvZm90cc1ZGIzqObRX20S
axgifru+lnO/q4G/KF3DH2V3eF6YNk6aOmhBScC4EpkrH4y/nEGYyFdAZd20+w+cy5qqwrG3nOv/
qqwd0ptqGNkdPKTesMpsJyC+jt9VB5wXzFbebmd6MdkaDpm5VWWjQpxwNn0ZONQiul+GN6hjSMbk
gX7t61RgNMUBGfMcf+qQmEpQxgpY8NOEJoKR9wCJDSUhTsfcvhNnlRutovv/nYV8wgsMDla4rUuO
lVhlozDUiy7eeuj/iV+UOWaS8DsNZ0eGpuVS40BoxJzgyE0LR1gTLTmMbCuAzmRu1oQBO0LUWSJf
kvXfGylkxfUA8falCkBuTMP2tC9Ix8fvNspDuJibBaIQpgzSfuh0j4NNM8wjUOXfHeG8joe+MVry
lZj+UbwsNtvxY16ABi8WITtb1BB7T7cBy0ADDzfvFK3L6vIiw9PHH/UvLermv4yYPHCXZMuOLtT2
yY4I1aHdqMX2MnSudx8exsuy7t4pSDoe9ZsLpl+xyu8stsiOYRff0YLYBS9Hw4awdLy4PCiS4W6C
vwtIF+WvBhwXLisZ7X7JIeBxxvFpUlHn7NPLTnOiuQEAoZkWOg4ZOxKYJT9WCMfK2REgn34nhUra
F1MaecNXccr1NxGKk+tHR52w14g+iue28CK0x9bgermQGhOnKT0AIDywoZwHZwQ3YapE/lWxOQqd
LPWspwbucSBMzVwZuuyiNJ4TFKClETQl+i8r54znYSPZ1vBfdzjBlQVQtjii8HjCKKh5ec9mTyqn
grIX8PfGtJkT/Oa7VYBDUtgeG0EZgAzGc2v7+rqmhN9X0sRgkod6eGQx1xXfqG+OoEUkGDuKQ1cl
VVonyx+hfyQ8KCEYkPug/KcNJHceUhtKuVl2FSJsRVCfX0JXaQvEoibemzBrLqfTkAtI28J1IIC0
EE813yE2jVO0lQuW/M4md+XomhoTmVDVz4x2giqG++FDvNyljGeBSt/3p9Wf1wfIq6Gr0ZH+TK2I
JY51VlzBJdHpLCqB0YbFjqnHl+dRwm/ZJbDQi49vLDAP1C9SVycSI1fwi5Jz72iRBJD+bK9XnzNS
7+Y3uRv67nK6ij2+Doiy5JHpB4EooYJj97ASJHZ2wi/Sm7Zz7aQZfpLaxED+5sI/tq5hUcpQ0nD7
QQqP9Waqmp4UD5/bFKQ3yxsJZLqTsfggwUitato7ssHBxIY16v302Ex+6YXToMogQUQQ4If2ZXz/
3uxrBsbrCEunB6EN3KQXJ/CvZq5WIn9bLA2n5ngHygNHSusWSa9eR3c7L2sWomchfa8tCxVYb6/M
PYstLiTEb0kB2oHGAuCXALaPpuj/as0aI06X+iuQ2F6ooRaxcZAj7ZZ463R8EfZJVWdtdw3aduU6
CDPg5ARUAWK/35NOFEiwQFlFk8WWGJ2awauxu00GjW6XNyY9/9VmUooHtgyluLchBepcF5erpFQY
nHjSGijjphJ8j/c3qY8JBH/4buqd320I7rHfetPYPxT7rB0KpAebDMMIXMpAzf+fKKUhYEEgFVPV
UeBWHMlbXn7gTyt6SlEjDfN1saa7ncJb8ghSTj8AUyiDEvrYxmJpAsBhhWbTJ+0MG07oBu5jRbVm
UOQqSP3ZiUSgC9AhmsxxyEH27gNFq8jbi1jXoLHM6o3aAIdThwIR7RmjyYCD6dv5ljun39u95ot3
nUlvVBpV/nZqWCYgAs3mbUyPUy5AoG+oj+97AI70aBjhiWp9OWIfNSN+NExHI/bBLpawttF9KGOS
Qlb/v3vn1B1LPsV1knBR8uf19+Wy2tcmGuHxbTqCYdAkDfoGj+LezwvUMgUhMVPZdN1Yy+BwIQwy
OEGjGw037uT/g/GlcWvUV7adAVA779kcrW2O11y7wDsg57qbH+BvJ15QybpIhIS3BuwYOr04V7Zy
8PO0imXLJ5MpdWaIRFGvjlYKQOhP28jjqhQgKW9sHS1fWZOiWO+paYBN4fF2mmbkQG4Qcb766tqj
S22OkyOIzcpfXe42Qwa2cFAyd51IvnyUyJETqJqZvugOy6PzkQsYTzHxhtPSrE21cWdnU9EJMNON
L7mqEufOWeY5qyeZTVKmnBhJwVvs2gRb2EKlLjZjmvIWOb+tUi/CV7egXgIGR5Aa4x8hmwOKysYM
ns8q+8WmCs15KrvsvaS+7q0bUCM2Kto4Y9cUQvXla/DxtwWtuj7Osa4QMqUgp/yFTnMAFF4j55PW
4gRNSaO389Y4V4aC2rM1updgwWKolRYyQjLGWoTLpG57aKuvzKgXH7FLpmpnGOYHkDgFc8BO0D0Q
d7FvHWVDaNtUNNsbSzPYYGSPRpdPPxLFzfG5gwzWlBkbwxgeZuYNfTpftbqDa6k5Js8eBiZ1fV0n
fwh91cuyIv6lKfN/bqpxZvpRzU6QnSmGsfxyP8kWMPAObCIXsrVn963CARXYlAeMo71/UvZDv3j5
MbwTA8Hiu/igNNxOjHek0atgLrQhQavjxyRrsRR/fHGiUqNyM5kLmU6NmDCjacSpOqN/QdSrA25A
/uCvZQK338YdNcFN2HBBan6bHcHGY1bI93YnHccoU4CCeqjJOTXMZCF/XBuaJe4wakRMyfNN0Iji
+/6B0PiJwLyAS7n1/jPB56x17w+v1leDCjSnAklmfz5EYWK052fdAmh0+w8Lx3KBM7fqCGKf2HcH
yyhHhOSxH28phnHeBEmkPe2vRQigofi0aorvRZ1LA5zl3IVHqxy/wK8Nf54IBGjdT0x0iJTNxHSS
+i0eaSOOOMrzdzYqmaYCmP9+qpccy/QJte32tMupjE0IO1nXaHBz69RqoorXgFdAWifw3xUkXyZe
Vo1E0gA/qY99WyYskKgUmGwvw67YB9GARMxi6ZCwTzc2kaAq1i3KyDGA1tcVs6pjz9oV6cWbrYKK
arMZagC3RZJ5bYLJwXbhYN3wCK+tyP+oxDfFCwedH5GWMrd3swMONBc8AQLXfpk4UxxHIzqdJnsl
2SkZHNsJfr0JHFYKEDdsv2/Leq45RI549MgQAT0Es6cxWs6JSngTOpKuHxBGrCVv0ReXVe0lVOtX
UCQJj9LRsKcvOWtyXE4g0YcyKzf+S3kKHJVo3nouVdE+b8utS8XmSY651Tgg19HelnZ7n20rvFD7
2yAtN2hG6I0H+j83gtJfYyo4g3+b3gUtvod9L90Wr4DTE68Qp6Rx6LVsrwyOxi7bPnto2HGMMUEt
U9WaYKxFFa7VIElrWsH6skGHDnQNSF1poABwi9IvHgfjtYcz+UyusL1wAB0p69JkZWNL6Tj5voXl
tozJfuHjlclbILprEtIT5QzaXfl7PTOS9PFCwdwW0JyaGRPL7Gs2UZwXHFforD7f1C4wnAfa/rIw
B3sRKe2fJyt6YkJpWgKWt0NKKvCBrfFwM/IcSNQHcdnXc0hkzn7w+75n8nFfDKGvUm6sXu9QMjiw
yFFVyY58BXjYz6X8NBt045RwyxkW/3EaNjPdn/rUSOt5masgtAoihUe6IWM1Tkkt+k0EsKz92cuE
TvttbVIBiv/2K6cptmPknJdUgrFGl+Ne9CnQF0yxIQ+0RSeHakrxMbua2KDMf9ybTBRV/0tlpyF7
IflZBwevUQTo5yYmoZxti9lQegchvqntOT3M8UWyL17ZA+7vd9ZvuNhvzPqZdX0oPC8awSEuSuP1
/IiGsWqqbX+89fL/ZdYIEMKQ3pRAfrIl5yCiJfXniorsODDFhgvWeLrv/C/CP1exgMJg3xWwHMst
tzGhpChwPTzcj0sYi/WTU3/K6rC1pWl+3xdqQ/6rLitRA4cFZHvzGvHZbLJPUH2MGkos5HCfVZeL
ArprKoGLGKnl6Tck4BWFeM2qTB5lOqKMuY9/K79fqQ6EzMbvSeZIm6ogvcw2wH6hN6sM06xifkzr
Bdtk5UOx8n8DE9VXC3S8cz5aKdS4s+ibdQ8UfNc3pDYSJ6WFH2jnKZn/L/lruUgzsO434MRxznsq
i5E2xOSW7hdIwhOtfNxJVRkbd3hKLhhJ2iyxkBq81e68SEnS0v5cm5bz+zNH6n5RYpe/npVnZun6
xwXLfp588kzKz9hWy9K58ZpiKshTvuf9Sq1zREGG8uT1IvK4nwPMVhCR+fBpUpogj9EHn4IYleHN
ay6XKUpW9/c6xmWTDBXwHlJfZBsfz58Pv8kGQOziWWK67RRQ9LbsmKUGVGJWU6J9M+BBzwJV1lDi
UIUf0gePs3+rZsF6ttRRT7TUNHy4WIykKYmAJYViZttV9xxXqWPVzeLkEAUxSvTYhCfeQC34dR7a
8JyJeDgTbXtt3ktimSQWa64wLivWgOR/ySHBfe6kokDXdgmTv5h8d0kS++oJ+YXk4my2kwg1lFRD
lkaVqClLb/KIPZfiP5EtfUZJG1zP0ekYxn6GYbvcpb8q5ZBk3o9w8D2m0nna78SGtVZw9pOTil1n
PsqgO+/OpIz0iaKUC7VXL98f017xfGOMT6rmZIEfmqqbmP8bRisHW9UGnjn56IN4XBepzyj8pn+J
uDO4JASeRXZZjMfl9l+lvk5Wl4ELcYcWS+DY1ZAQ0CZaptpxyxw8XGhikhpPXH27hHIVAi33X+NV
PpIQtoj4bWjNSqsKPIxv25cAHGXL2Y9e6JB+hBc6RAxRjQAP7V9kSc8BYKn9XjUVquDvk5cJ1t6u
WBoY1WsK3kraAcr3dPK2BcBav8AqiUZtGpan+LGwKrxXVwpaTcZBf4dLIylLxQDgCnnfTJ+i7pK4
DnNJ6QIjyWmRqzcZTQKLMWxwRleBGUvjQqnSUmKTWAFlQCv9oeeGic0XlS/lYELPdkhd2sBClynk
BDcqAdYmwc7sGMTR3Wt7wJzSmQDTGM+EtGOifdxexm08lp4CBX1/TKDhJEFUVcViKbIVQ5Q1tLhY
XoQtnWbOc95m0bzCqC85AEJvD65gZja9d5Mquu3+VMFwRMpR4VcJhJdffplgupKgBVy5rcOxzl9G
1x/HPw8C6axp340LIP5EnwcByk8blCb3v/HXuHvoCTLqna+r8mgjKKwJfvH/R26K2V6NpDHYrH6x
A0XbaLDd3wn0fCwNmv2AKvBfHasWci5sl+rEFl6NW9vpdc0YIZF3bTft4hEpbmegcsh+WEE/wYW2
xVVZg/dniEQiq1TEGvbIGLQQnAhzIvirpfWmEm7MIh5WwT8yIZqfNmCUMtn/yN9WiLTti1//voHw
X6sceBWDzK1ANbsap9nm16W2ZrYWKHLc/g/JWc01qypi8rhtdTnsMl224Amsu73oZHqWTosIvfCO
a4nJW4CRGSrcy52fYgwqnNlktyNryBqeTXP4VcqRVO4kdOV+UWG7/ThpMIGOnCk0WsbNrcY4T4xv
iH2GgcTsNkMzGa8qOBFwn9V4qwoddqAtAIJK+nBhe4jnSXvGGOpXH1bpBrVhGpNhKpcTL7j2lwH6
V5nlHtDSeGkIFdCjzRPuF6fgtOgGhxF4Dvh4tT3wJKuarBBSJ2gFkGpw8RK8UTZEfDD9dlyKcEuh
ClezuCfGp6Jn+pK4QiIYNgZIyMHvbVY0b4yKNpUT7y/B33ZWm82l9E0Lh26pSA7HC0Skc+0dut1q
jVIvyrbhAsRDtWMjq+bjqePZuIUj5gLwLkCqgwYKmPZto6d+Noej03f2b9KKEuxQQru2T3bPQeB1
BsiifpN95Ogx2iuK29OTUYCPg+t3yAOP6Te+py0dqzwkxhztQ5H/plsewGGSx6aqHxmGgDy4XbnY
UUwoD8fi+E/CHYLopRRP8ejAcjP2JGvoSVQ9lV05srLcOffvPYVTI6v473BIo6y5x5Fgd/PCYbbA
NSTb4t8Dcp+UiMPKFp68JJlzrnx6zGvYfucZWEMCkzB9tSdZCdEmro/o/Lvpee6E2QlV9E4Vl5Y/
NQtTI10UUHMC9qnIO/eB+3gQHYY3HIFgoU/bMNs2oxxj87Kd4lN8xiKguo4slqL5tKop60e+TiqW
eENwUUqeA+WJY5vrklbn5ceP8s0d5b2CzyEGKNN7RMc/WBW8TAvD1OK93XoVKysLWF3MbHpYexyS
Y6CpREqc9DQPgE9Bm2dDb9LBVFthBpO/5MrwcH8ga4SGZwvgU0UljScBD41R+UUBZAftqZYNrBoZ
AH1V0ZudpKy6U6iWxUxGg0W6eGAxGMNg1y8C7srB/S9Cufuy6ebmXgJgyIdr7+bFjcfQDn6eBwzK
r1+brE/L1uQhSD2SZAD9k8SD1BViYH+f9IV/gH6JAHHiVPE/Ayov0uY0/W/JKAhG3BPJo+7+AjCp
9KzsfP8GZIXI3qBtbTynkJ9zsxodwJuUVvh9TiN8UNXRM3Bu83Gafj/rpgRF6pqdtpOrTj5tsbXi
rNxlnSBmWJ0xiAzDSbktiDH71kwVKl6kmEPJc3rn3cTVkwLoJLzTYDBFSaYf5PUieboLxuajkIqq
DwrRuogbcc1wTcf0kOlpxguhxCHDF4dyd6vf4c4Db8PvVbscDh9oTkpGpIo+c3dyy1vNnT68DtGa
TYSoWHJqg+k1XsU6jiyXryAFfw/VHD8bH3jArrp/5gwPx1/Gzdzd/OrYn4VbvyIkOWXjfhe5pkP6
9/Cl6Rn6H0RY61flszpFYPfPg/CaAuLOGurDGL476N+Nk9OvmiB8lSa9NHFNdacf/GNb8eEqpEEl
CLYbHiD6pQgWegazPi5VgVUCUTF1krMKQ+HfNuLCZn15CKLbwzwXx6RHwXuKbiM8WxlmErSeAc0A
F0yj5V3nk5mIIkszG7yKHvSIIq9iloSXeie4HIWKHFQJxIUUn4yRQqDweGwD/oeLusWDCgKw8yNh
KJ7vs93fBF2fabvh/FsoC4pdvqxCYxQueeNuMI7hkLQiq8BTTMCOwoIOuhSUriyIrEukJMbGYjYm
O41tricowEE3ADMteCokODqdqlB2YmGjsZfnVWzQiYSweNcvyO4mqe8PNY08viNtz5Vy/YVTxQAs
jJCLPR3hoyksvb/T0OaCD1qfWWQDnjXtq8MIU87d5BPmgVbEYBOTQOz1fo6gUPrNcR8DpoUCrbuw
W9B5r8i4FbQT7OTXzpEi/mEjjqrxjB+qPHCbykQD9fC330GaKd3HtC7tcSGALzafDnxX78abnTtT
MYeopIGdpaU8qvG8KWHrctj60325vyTA+ydZogciOPwFDOqsp+onr9qF4VaUceIXoEi+DgaGXo6z
ZtTq7z49uAmXkzzu/5QaF/KH08HcBpTYg0eHFp4mExB5YlklCe7P735Z7zGnx+beXqRZ6PR1OwFk
qHtkJvGOFnEcw/YobMveObpCpSk+3izpAF4cauRlVp2MBFb0PgSEYidCClDz64Z7EuVaLPSXu6Xe
q8a7zXbMT85Eae3RHmO3vLjtXQgtZw2W0f/TR4vnsgAmPYkpdNRXJ+NUQZjeJwx5knlJcbhZVbkk
90/2BUR/3rGbj0KTmbgXOCmzAeBVjYwj7ugZ6wwKZ2VtwpzRAK53tpUMwI7QRoE4lbfvTLGyWbbI
mNH/sVbicYaMSN21Vj029Trng9Bp6BUpd81QF+xskA6Dt3k3HDdRHi6U2r054wDPJCgSp9cOJAkv
Wjq3RxdCGl6fO9JfdALhLpqDUMNHWtj9iouuv3XtQrsFDiqilywjV6uykb2cQNRvolMJcQZKtXzy
jsxG/iCF4RWxdKMlI6GJVhX1wVtZ5C7L+vIBGt7hC+B8bmnERbmEMnkkMSNHHoj0+pj1IZ/BZzvN
F0OIMKZe8eMxIpIgUTFQEHR4IoV7dBBbA2zxSBUVLqLpILmXYsArcUpOhDQHGH9pEgFZhQp5Ivlv
Mq7w742UtVJHoqBP7uFsWlmQDQfp5BKnNTFpB0p/YblRaI/1q04ZME+Pyu9bK9g8l4cMu0azKeAT
1yDSSx1Vg8B5hV4w/YBJWslIowzywMenb4Dqowe6yJ3zYbRvkgRZD5ccUpVsSYYHSd7qTP6+j+75
FczryCpmiEIL93SibYf69LMlMOqQD/Ro9o7AQmwfsM++S0E+C2ffNaSo05jIvL0DXGlqP6ubmKKK
kYTy4VD9xpW7GBN59xZRzzeIARYEvm1FlrgDHi+I00i9HIqcEm8iUD6fnxz6pU71kRe/FiidPpjo
vuGTCJaWkcEA0wTM5m2VcmDzQJilTDMNaETI0qICPQbT4GyrNTm9bL3t77pWa5Wg87IDu9H2X50w
BWgWvND0NYq9fjGsbSj8UERj9lsBe2D2FqBCMQon58bL7Z4xfk0K+6kF+GHNtofpNNJ8Z75dwHCu
SigKdVRG6eoHuaUGuPyLTRGNjpZG8kV5DGEA/zqRf6ZVaNRUfsS0G10VWMh7iPAOGbB6thgVu3K/
lajOFP2ILPJJlE5yATvUUCSlzvobqkYa7tDlHmSD/l4o7MUliAGVdaKrnUMBvWGPgJTToAGN9qML
dw04CRULEv9jm0lqBdZrNIoyy/Ud1M4JkpN0EO+HxX03X1mg7vYKcAuVazKS471/IcPeYWn8oGuD
/cRu4YcCNkpJNRUnTL0dK4nG8l4ROUHrL6FGI5m/Uy/kIY3a018YxqazPwmX8WH7EGMUnahpzi+A
R+SQpBjLPdtGifQiTivquW4vDxRA7j3nJM51Rv4/nTGnyxaB6f/SK3KG6fyNutkcmFsIgjAtklWz
XS1sXD963IRDTZaeV2skPHspMIItaNIxtj+j2T8/Bybg0TPyO8BXsw80r99/EeZSl/y1N78H1yCf
u7P30Qcs85hbzQnAR19UBEqyejT+qY3IqG5GGDlg4WJNgq8X93ShWfZUHNWesajLdiZNntaEN9ro
bt4gmoQi5YcJO0lgfi5g/PPfmu03XVPRVAnMd944Ps3jbEFjvpf3sB3FMkbkJIezS+Tas+hpvUiZ
mnqRau+P+MURdWTUaX1TM3E0u2XKnT2tH7gLJolplO5WF73OuIw0zbRn+PkS2cyiWLR+g99IoyCV
6f/sHWUrml1GkhSmYhYTO8U3Wp3JO4HdbvJafjgoAGjf73H0TAH8sTa0dtvwwOUJxh02F27pAlQS
WUAq9ZXHmwzGd6w3qSr40RXpsuiAMSlp1ShCFk6um4avvkaqO1lB0abjpIBbjSFrBPmEQazJPtOg
BhWhBXAvzntng/xsCEiitZ7GhA2msnyRisUquHr2DwyHC8e+Rqa/R3LlhQUgwM+jobJGrp1uNbCM
u6pLrcPli3MGfcXxrkJSOlAKKYzCgVZvyUfZR9MU8jGRIjitPuay0sMSvpzZ2DBFc7DgZqmT98IC
Afhrz7eji5/la/7Javhy4a8zKGbJ3Kt0WmPQL4FYl19S5LnbM/N9c958OQAjIuWohClydjBznHb6
ALy1I1wwMm2bJWz6GM6UM+KI0irWp6J8VuP5FniKrimkMYqb/ATD0vbxQCLNvAaebfKj41eMR17h
zoRzBfcOR5DQdoaPWD0tijb2uA0maHpIjD5fQceT3awfGpouuxiQaMa3pz36kTI9lM6MoKm63foL
YNg/ujXgqtzAlrbPR6ldLEthTof0kwEKRQyzKurgyCPJTGGj8/bVRQP2T4DtfBbkxmSXrRfl5qS7
juOdTqROugtmPJOzjpQEb3/m5UpohNkjHMQID2OVIao2gyO7pJ9P+qsC0cJGUe/+3ex1fiEkb0TM
Pn2UPKmB/QQ1geSfgCLDwDU2YSopM4p4TnVsa52WxUMWzrrjhQT393sfJwsZ7HiM6XQb/VJCKaQR
V2YDNB4qUW6M1oTv3ExmqGNsKLD7VotvmnUze5OhitQzCiexfdjyh74oQLXQPjK0UQtsKzEclWMC
jzc0RxiNVcHXelSqrQjZ7pcyIx0Xka+42pq+VJqP3BoONvlplkhn/i6boq2iNAkyTpY9K8PqTAVh
RwDV25kZSj6vYr72+cl74tVAheHz/KvBavwK4YqtJMn9B/YKdWWwnWMLEVd9nyJVW8+hUEX8mSMb
qNJPxN4W+vAdaNiHq3lxS+HQiXS1Texdzf++jBe94ll0nJZlwg9yiSlDrpLaxK3wfmloUQUVku+F
HlUVpwF2G2HROLhXClSn0wNGmJCJEInZ5Tp5kwF7zAnvr8ZhLJx0YPF8dqhKMomz+fawKbj9wh+i
AWD2PeHqA2NALcCI0so7m5tPNWVfRgAQ9+2Emkss9+EyHvFenTotubCaiP/tNVEk66u70rjJAYYR
7TOUbJwlK1+dY6EmPaGmbOW5aFB+mR/W1UZq39sZdZ9EwlnXQVLKiXHlbFKOeZyLo1gJALXafqkg
cglAjlzTVREjXGGjqfc26BnyrwKYs2CiVzmUuiz3gDv4IaAoAsT7/iE7pfjqswV7C+0JCvWLCSMp
cGFvn8N1hwAXjQq3tlzhTBZ/w02shv6jSndl0jiAoFHUESc1wfbi9OvrrjmvlC9yX98K1T56tl7I
1cRYcVyFn0g6sJdanYta5U9D17UkuT98tYgEzRJnlBCh4Kt9tQTnLDDIn+OeVvMhhZVhcJDqwWT1
SjtlZzoudryixVB1WHvuaqlAYKbvdXzJAItQOotGRt69K/O+QdifNYBzSvziHsydyL9RKB/8AehX
FhIpNe1tQvXyG9kP/yTxVQgt8cy9TEhsiNNVe1l3F5bH/WIPGi3zNu5p9YGSNHDJzw+kxc7tQ3QB
19pw9cJK0WUr5AOmmOUM8CSWT0HgurBjnKaVyHWvFyiC+gacqsbKoqNPzu8Zv2P/yNlhoViDut+8
LAFXAyCpttT1CyGtIn86Md0Jgx3BNncZtwHNuEb0LjlZbJ9hY6zyqdsKcomKoKoEa5xIE3ymgUSG
gkCqXjxNJKkhn0GDsI2r8IRSNDtxdKAdj7AOXYD3BJqo/jYjSih8vGAUcFEyo8yK/9vqj0HX0qAe
tnP2klD9cSAqQFlrny+e3GJD5LdDkaJaPHODAl66r6tgm/2/Lqk9s2DF6Vo+vYe2BsPhkYYTG4rs
yR4XJtsPfQ9BZQcH9eraYDhl9lDzzsF1V9Qd0O4ogujCt/G4jRxLeda8AtjKTB4gjfX2Wsy0dQX0
9XaoHiQBmO8nUme3Votdtf9Asx1mm8ass3mmEqJ8TCSgrtFoqcog2jj30pFn9zB9OTTwFmX/3zr5
xRcIK41gza7nSdlViTHXNE+JZAXYFQske4IegzfnLyLWFWfeOL1D+00lm6riNnUWIlWrkhzmjTFp
3fp4i9ZbPgol1hhxdULeBgs0hL9ZOZiJmN/D0ym0lXUUO+xkmCvijxCwR3vZFBIQWmq1940jnuR6
3W5d5KlVXurjkeapdMros2ipNRtjjEJltA+ftiIsd1DE5Zr9SlSGTZ2gXR5yncBSqklHOl0yGwj8
HRkQUTfuRVD4mnqNuJOtz1MWiCUt0VITbhwFOIxdYsACbLqt0dKshanZ+lHe0ajplcLhg/AoRMdh
vNUrYEzClazX06qyZy/yRk3brhKsRs1ootI+tLY6ByakTeVrxWIAHa8eizEglVlSmpBdb55OtVPM
WsP43VP8ZSLuIa3KcVwVT7kSkm3i8Q3/SBetrBGj9AJJHcHt3sl9oDyw6sWdrvYKDGcBoSbjisU4
Tr1vPkGL5hkLW8UMx2cY4PtwG4U5kC5G1OYR+FRKsBPSOAmdE5gx+nqTdBgA8BZhzhekSyhj/k0O
fmSFFU7Qd8f0D3mxoPVAgAigAHSxJtJRK46ddfNDq/TZyFxZ7wzYF+8a9Q1R+UsBrinfl+DXHHyF
CkIEnQ/wgPPwT2wBC+Nichkz+FUpiwakn8Rduc8g/WKWbqxKYFUSZ1u0mp2n0PjUbfAlWki0/UXG
w5LTvT0lhK3bJj5B22XER9VRjNdx7ahAZ745+3xXSPVn/MGnSozciOe+ifw/G4fGjsSlCzqx3KAQ
0JqqdtIpGsw13axrPOUt/R01vbMzdR026LPiQfbqzxioQ3mFTP7CH8ps7jCIy5sXykpRSFT8A2iO
Ww+wjym+ROGYTtlKSkomKKvw3QlQ/4YKXQ4mgXjPh0b84MXC8WovQZISFJM1KUahniD3SrE74pNv
kq17+x+gwzHWIpYhn2mKcXvQchmxf0dHU2TPV2btXEQNrfJJOc8OdrAbnEbmswlhzQU0LVciynvL
4VPWiTDeDRMTkIkmyEv9MSe8YrblH+8LG11w06OW+N6pj84HRBUZIrZ0tiP46E8QAkMjw6mLyZlj
8EJKYmSF1HgTu+rLqBDoQ92eDX+2Uh1aiBhIAl90mzbcobsOw6C7HRocUEN//sxwhRa8dBqAB7Wp
LEqPO0W0EsqnJcCy2SNhQVbszMjmzNAA9Qd5cw59eT/S0xva3nlGUUzgCN9TLbt8CKbfmZflBZNK
YQJMu2gXNFutpRVNPuEeRlkT0aHXTgIOWrx0In6bQc8js+lkYAgfAsVtpvnCJlQq071qdlfINE2f
3C9qm9ST2ldq3zZ7vCzvAEOIUdvEqgiwucjQBa6sgfzmEc0D22Q6Onu6yz4Yf+YpEThSOhc1qfSh
ZceLOYxW+TG4mKxWHpXrUKgKwO9X/sg0c6zfrwQ+s7k6Pra009+6wjc3f0MmdcnwS7W8Xc8puXDq
A7nsLgNc0ij3pzvh3OMB3Kez1jVczWrFlo+pFFAg4dXue5GuM4cf1pJe9ZLKByysHnNzrHY4X+za
moCutxzJGhbVfIu1YJuQzhSKYHqSC03nclxTN50J2ZM3Okdea/yk6Rk96uCtfBwZ1uPYXHJSClUS
SbINtYbXuStn67RQZhU9YHb3QMCJHZmEnsKpfBo4TCM3D656Nr+02ookCvUZbclPOuE+9KFKs8aA
h4YNAf/VT6c1P6IxviEiiR0AONNd1eOMiodwdGAUcDm1hfJ1JOzmycr7avbBP423fgvUQx1fYi8s
J375TnekuxOVlwkOr3j5uBFFWSxRrzz/762aDTuMJV++hvhYhCgY9OVxx5YBOIqySJ5aI23GoItC
EneTDgj1q9ggEQEOFppNdATQyCdOu53e4SyN3vzGHUHDOKJAO/xr837VB+UcG70HR0gxIT++OMQI
86hY8+qQawv6VPsZ8JhcvrQchb2/NksiX6UMiXVH7I/tl4/BUGrk8R+mvZBJ/f14VA9S0SUZY9Nm
nw8z1SEWQPdj9jOF+O5pdTmeVi3Us/P+bsuXWGgpZ4rNOAhy3yAPd1JaJjiHMUxPSVMxt9tfhFZs
NfdFF4IXd028TnHl8sVJpyWCoXOJMFjkScw5LULOYmfiQ18pCvkTgMuLdsZBXVV7D1q0C2LH+DBU
psxNeNK4KWpcrCtRFLviTVUKPVSo1mC3jgbNlFYMoObvpic+pC3QzIliJh9Eg4WFwWonDnFCHWje
vJUJAapYHlPcT/9GtxdGKJQGO79+dOG10AI//vI9dj1qMrJIxQna25YV1Pg8BVA9TUnNbNNx1FTw
1Y7TKfWUq3+ogiE0rKqGf9lI0s/1gqHwkZqDivmrvL4zgB7lDPJfmga1vjXtmEJ0tsiINNU4oMED
BinjpUiaRaOMmk3FCz1/s8MRrof9WzsJwGI69YZpMd2hawSVSh3idv2YhkKtgPza+3+pFxwwbkqn
+uLxBqFuZKpB89Nwty7Y0rX6A6m12ehw6YSIEmC8Y85WLlSO2M5qomNBe8fW1TSwIzd84Z1Ndc5S
Ia1FufUWeoexzIqnGX8FOJdzojwc5/tVrudOkyTfmBYrJJf+VFJAnUUVwj5utjkhIfDbv07BlESy
u1MVLiWYu+ooTO55OCuZ6i2YMf0Y4146Y8AaafGzyKDv2hiJOJStNx5/a0vBI7PwVLGFTDepJLxp
83cU7iQ9BfS3aqoTqvSVnYvFJb9/b8rR9dhed4CsjUNlIaguoUF5F22kmNJ0FBuvChHymQvO7lCj
Q0fxf7xrX6td8Ece0mVtEEr9fkbcErwQX4fnbWpHh9O9YzoK7f+pVk9U3NmH/qNTJwCWM9DuKmnm
aYiWN7g5mfOJU0pwPihIXCNpx7ChJzIe3nb2HzAe5a2+hdW+NaeLGl7MNoM2fX5j84mH3FJolnMM
fil0Oov93vzNX8uJtpYhVbNNjb38R3j+UF7GApI1f8CJTMs7XpgV3RvkQ60Ov4EOzZzFDFlfKQTi
fqOlmI89B8QnbrlSO5c7CHk/flUZnW0zWlYj2cbHUk8wv5Cbsp3lrYeDFkwnPMtHz/z/33dJHZAA
RfGml/Y3qv/tAKbCaeXelgwjzU/NS8wjFgygnxM1hX+i5TYsEYZhJyYnCTW4vAPV/VELNkiEnVQH
huoClAYVGBV1IW4b7+80jDt3a0n8UoibmB26deQEFvW+Bd9sqB8pUfVWKoP+k90vjq6OY000nYK9
ON2aIv1LklvzXbHMNZs8GcWedIB321Q8cHqiH+wilv96KL+MAGrIgUsK5xssfobolKYxRAc8q3tU
tWt/F5MjeI2sKTTTL5hSV3ekrVek0HiwtetiKXZgxLo4Imc3pXZSgk1PuC1LmxDZDuaDLorTN58S
K2iitTU6D6ugr+CdBph/fweOkSRLSMETvaWlerTzb+177AGfMVjffU3mphpv0fHxaK1mFOq9qg7Q
kxwyHea3KRMfym/JaRuxegmSVuQTI2YZ+KvwAEeAJ9Liu+KxPpjlmVziZcBL5aBo/Kdqbnla4gwm
U9jV537io6zA3zD/38Pva5WHsKbhiuMzZYkmRkzd43CTxsGBMk0GHt85aWOqfltUhBOH+vtweUEN
ynRU7o8PLPR2cmoVI29OfegW1C7bQXZYYUelVcAPgVTIGSWKigbWU0GtFEhnTW00/w04pT3z6TLN
4+UN0/0p9PhdTeEg/CoC/91C3kaiowVKQLJBKafLmh76l8mvlqVFcTkX7EsG81FIo408ftQfvVwT
unHiSvjZAxPax3ZbXcl1tg3pljI8VlgzzJtkOWfKP3bXtWJU3JbxFFGdbGXz1nXBIvNOhcKDgdPc
UxsMJjlpeC325kOZ+Yas5o1WYmhASldy6SIEiVRC960XIlaA6VGFIVxO/XrgP/EPP4FLnDwUqUqB
2J25NkcGBOxbS5cWOYzWmxWR3UQf5yABVRrx5Z1KCBorfc5wmIwK3IV8rrR2YA8b+z5ms8dk+QGk
M3nUT1LS4R+31H+XLoD8HhqOb4aO46cfALW1Q+pXjH2sAT7mCvFwt28YbDA5KbItYJ5CC8FXjEnt
9fmAXqIM20P98LUiXTTTP/9OwIorwzl9PBUdVYhQON1L500jyf6HGeBcTZdAxH5VNxT5MYikAiqm
U+KpXBC1WG+GomqhBF+jkeVdgHb/gtAWZCgkx3V697BCIIUg4AZmLXtFB8fVs4HQ3t5vnSLSrBvM
Ml9eqBHhcfANnf4SPWCMxPSTf4dVJ6Z83fd2pmuF5DiX9//OSk+f/mVOqXvrTX4lec1Ns5c5l4gf
75j/u1F23WQguAK1ywD6I4RTAwCP7oyau5+3aoOyAFET+sQLoy03BJBcRb05P7jgD9WZLFKHlbn1
AqzaajefnHb80GQigTS3ZoOzhH6Vri0T43QVgK3v7UMGRq9rZxIfz0ygi38irO/SSuVusz79wsfr
JCvLEHpNdDr+Ne90qujaWEH3+U0HNkOtyPvpyl/n1PNQJ/SXZBAUPBXb/I54SqRlH6X8EDFO+tbs
Zr4KOQmCm3qI/HpARqbrvjbwSfX6D1sG6KpYqxMlJ+dtzaBGk1j6ZjlKyZxSXdy1nYlj+IxEYIsl
eBriMdhFqIySOu/X7AiLO/os1+GiiWSyTeHG4D3vvLGuK6HF9WOxl1Gf6cT4Xdi9tS2bZthaLnMw
YPpRhX/uVg6LejOzWiUs0sJbTRIuB7RZSXg4lYZLZu9UsswsXz/1viD1tHxgZ6nPBgHLX+wA7yqo
FKOb7ohKnSPxMtoeTEc1LTYiLlDblIJykc48P6ov5rtoUHnSBrWz2IT5rrSqFQvw44nYOcOOF224
KyAcdg6j+JgtiHynoUWJtnpy4dM2QYLZ/f++ZjmTR1ILKoJeOTFEbJ89ok7iXwkz7Fm0ZqnaQITy
P6/Ub/3yWf38UueBIchrG3lIZs9l61n1p0YE9ht395rwMtBVUtbLEnTJG2oEEi8sIxqLGAwWKggT
SxSvp528E7GvbVo+FB+/TNVxPKetkPDOd/NS22FRtxea/7pbh2Omw5vdLrYdAu/pJQSWjSTdlbck
Pjb0/z59jC0aF9PbMTJbBgldX++wEqBQmqJ4PjPTNLYukB7Hap1IVUfzb/WbJ5Y0cddWFvA8nQh0
l5+SCrB0sAH7GxqXr4WPdpB+8vehS3iVGpqHlJGTOjYUSX4r188WppbNfCGkpbpF1dC8f+JRyzE8
JNFvwc4jKj9EQV4uaig6HVtQEwb9o3QAqur//zLuaox8dJSDuSqT8C+ti5a6fp9x0VrgHQe8P5+L
e1wC+LmS1KanqI64pG5qpZnlfBAmtkouRUuL7SJieaUpEje/Aq1FFgDo7poAIoVJAxUc5o1DA8hR
4GmSGiKDeV6huz2U4z4qoyWu6rOAG9XRC7XOwXDomSenhQTjA1P3tPBSfrXD4JElARL5yYpn3poc
DRz9BYjCXIrH64ONf8EU0SAq04Iel5bYbVeZXlvZ20gc0gw5TfTY2Pl8YBjh4yfWDWf3W+xT1Tns
wEs3paK198wjBKbKE15tqPRykFMpb/66ynY1257JPjbvSWmEN0n7Jw+4EB7ESQWtHWj6q06MJl33
DWfypO/yJiCnHapO34HeREC+GlcEO1ZV46kSKAocDuj7Zj3JnaFkfB9rK4cIg+uQpCpj3B4EUP7N
to3pyhrgXUOBnmsubu7GbDt++qsyYzdCXBMkAg4bZ+C3AUldF37WHm8TV98N3BYdSPjzqaod5Lmz
6MVyUJpvYeh99bvfLlX+y2I/NTsAVblpoxAD2Ye7rOfNnXxKY71la0Jjo9bBGc9TvReEgYFJCkHG
UI4XkBc+TTlT/xpd4k2lGiJVLXppTTujgO5j4PAW7WIiuuBdH0N6dh6xTl8XbTWe99HnvB6WQPOn
0QRvZcix4ZkbMKL4AkjdlIrHbXqZ9bpSIF8tj31mFo/HPDMlAicGlZ3L+K39tCm2g30Aql4zkCnW
L41VO6115L/qMn7B/RJj1ruNUqXHgLHgBUaMwMZrjKKDNaiLlZtBDRnb16Ix63QyjxZwAc24IUfT
7RmOOkAPg4riyaE/hcsBp6hvISi0v+Lup53XhZNpAxBr4Nwc8tBSiY8rjVE7D6VRk34SIZyEBSkQ
I5wGa3hx0vbJXRO93Y98yoCVEwgz8M2T0aGg3uYq34reGPkxnYF4rzuPyVK3EJ3IXcBVEMOYbWTh
CvBaiJPbm+noi/Qj86e3LAO7iIdMuLCdTekVE6J7iPzQiHkLQ76nr7FRTUmW2e30/1YIBqnEcCET
7wllC5R65e9AmYLD2mq+/NkhWpDONO48Xw/uRTihk8DpAZkpmuSQxVZeMRsJ1SlEC1OWTlxfIm6E
QC15PTIZ1LT9KumOybBFX8M1UA8NDroJDKrVPYdJsR6v4/+9G3UPm2hvSHadGR3dfJeG5NBgLU30
EEaF2Qp8NC0sjgNK8s5oDgQ40ubD4bXKt9IjWXXJ8mqqaDgBfuUkEWnGwdir0fab3XN70tEO3Bkh
+OB+aAPlKeB9/+7zJFJoi5GN8VgqytRfpfwclI6eQdeRlyKQj3P+Gcq0txKnJewkvPl7IfPXpIc3
z8f2fJxmK//OC3CFe//06+uuhoZKfBwnLFPeiZ14nsaWVBowj/6aLnW8/SZJQq90idFauQtMULiq
1bxh+BVHPKB+0zGtudrBa2G9oB+c6RsKossIx3djssVjk/v93xIGaT0TEHtgoOFXLIYE12yoUxUB
T8TUzcLx57mcUG81zsfKU2EWrgkGBTet/FyBUb6ocqHjj4HIcc0mmld6lDpqmwXuYb1UCs2wmlfs
YROzU/dzrG5HIpumuUPPJD77BIAknhClyiKr6ORylmCmaGzGHUK+iXvUDUgL+HPI2NjphBaijkiX
maALLxaUm6JPly5t2a4JMkF7jCvaywuF1lU4j9rKtWXyVZOjNcLOZv7V7cQqfN0VWypRH4VIY5Ns
yeljgUDltWFptqIfRFTtzzls7p8qYKokTvM41vq9C2LIWgc03v5wEmIYrgGDC9ZRwGF6PFIp5j5a
sVgXA2YDhqw/aBDRH3vwuQY8nfUZIjttB6LElNi+dya/B+XHWT7Lo2miq179dxk4ih1385NF42oF
COHoh8Tb+KifcQ/sYIwUwqiMauf1xQoll2N520bL7ThPnfIFY0Nu9E+xGsy5+BurnqhrSxwOcu7S
Oxqbs7M9MevkhD2Pwb+yTfIaao1/1i9a6D79/L9+tR9MO4UdSww2PyRVcLaBoyxIrfKSxHflhoTr
85ZkKCWEyujcvuTItMcwFuAHKVpBuDrnl9Bk3p3KTNMlpOsOMPq0oe8o0zw3Oh+5CNK8FzUH9pra
twejpCa3N6AVHb0lQ67S1Dq2FrjSnaL8uEqJyJ03LzpTX1FtWHU2Mppe8mUqs2p5BczGJyvXy7/S
+P+z1v8DqInH+wzgTINVl4wR8m1WB8xrztYCFO9fD09U4OJ5w4gT0z4fchpjTKu3UqZUZB6i11OR
XXQ38v4jNq6OiIO8C98GLsk3+dtFaFRzT7aEm+tqDYEb5/jG+7Yg0Nqs0QZQU1GmlFXWRoZcaMVW
dG7xDjQLntjvqkrBtjqfSvWqqaRiveUS4gM35fc/1htrMxLiRwZW0MLq/r69g3lV5thGyS3n8bh2
GNWGExW3tP6eizD+Vnn7NH3Uz0XqWWnAa/O4U+khXNqk55HSTYmVjtCCGg7KLBohtIq50hRu7PSl
MCXVR8cnYgonmFZfUdqQX9RQES1eETE8mmImC9fypE8/H3KXThDVtTYVl6a1dwcE5QpB1gLblnJw
AUTR9pUKtv3rrprxP8/9YrrAj3g+ZQ/zPUwTayH1J60xHJn7frPcGDis2hlPboVByUj6bqLHGHAC
ou3y7i6xOgPuMyGn12QmcBOaYxLgGWTJedllcpKJbay92CH9W+0k5Xvdeq0ALcUn25do2WwAODQh
4aLtovKJm4TledkETPNGbGxGSruqIgtzMrEF5PGLMLUjX3SZmR4zL4MTo9IAwywX6hQli5AZRB7D
RokrgWO0Z4pjB50bDr2jWZUbcvGPAF+fueFrEFWAwAMAN16mpokCq12dnGsubY2emZda5FzHrm71
F+Uubbv8WLrp+4+Mqt+/IZLsRA6E+zQsYFfDIesgz+b/i+/ZXlg1/ajycfLXAkvb6m8FkmWFEZWl
7aoN4QjjJKOUD9tPkUVJgIRQdCNXky6ijphqHx2CL+AoDtOGFqbPimZh/u0nOsdjtPPlhij+lNwN
ZrPdU/mgknfEZa9XVJZbfuEa34Ev3IAus1XZ1L4yFqgvz1ch8iBv+kAbtB0+YStHN6RmV8tuj/xd
MParrN3TbNfzmK3uPk+YFpwpa5/qZhjZAqpLa8TRRC0i0V0TpS79DY8Ck68lx28o2Ju/M19IX8Z2
DCGdqkOH+K0SKl/vn7KGfZF2m3sIOUtyfJ8yReuYvgrp4Nw5Jx4dBVnopCNf+AdVODtkBsUr/lUa
bOPPHLFQjMZjQFtVEhl89QbzdZaeKZJtK7BughaIBK8DZ8LSsaxTnvf/iuXzH+i2yS7JX2HJ83r+
pFhgVPdbveL3zqM0agGErrExJk5qUOUVSEia7D7IX3SqMstHkMNZ9i+LmNgqzRRcMsgpO/cC0odl
lakpFUo0NdqGMJXeVNWDVFhS9zDlSqvANxaA1uM4JckoN0gcdv5RHkCs3WRSBJ4eDOusStCXwCKc
24HRkpqz4D35gWpVcf/wX9TdWsQJIgTEemaK82yDUH2VIgr3U9uqGlt602Z5LcsNLr5qcrrxGfQl
pgEpU9WEoS6iuLnHiqNMfP47ZG4A64SjvcuFmhfp2RH4/SkmHV+dzf3fsgQqLDOpcofyUi4CaYq6
+gINAw9/RBN5nZjfL65kwbtCmY6H5lsGc4NCnTWjBi1itFKu8JEyjOaPblfhbjqurkYWKp2HHLqn
/CGl65l+8DODf5EBAHrxwKxoOp9X5RJj3SNNPOSFhbrvU9gDAamaQktUJd23O6PQqV0oW+hOHQuz
eolPworPA3ku/h+YCltrVci6laoXqSpExsCU7gflubUDyksUAPSoiVpRp/c4xZRSZ89qN710lUuI
GcZ32VSzvUO5VFInEkH2zMKOetOb6SVVRxNAeZTLt8NqNswiKbMLMozRkPcNAdgMtpy+2U/mIB2l
go2a0BtzRyi66J/XZG+WMWQYxDA/PnI25M9z8otaP/j+uwZaFtGQ9LXIgA5bQJQye6EHV9ofcBK4
uJL8NZtdABNtyOC6Fm7kpxnZiIdvxKPpCGTDDeADtpauH7i8yVXvJX46KcjTBAeDX2fzC8Cssb/X
xLxIeTXreaeyCTOW0+UdWQtP9XxzgkkikDd6t2fJ4uF39wJ4xX6M36LAM5hWCCwjLE1+wlQsWyU1
z4tPDMzmYG/w/YA3rxcCwE3O9jU7rKEyP/iSjqMPy0br0LcDekTOqKGLZfT9aVmn2WFo+T1UJ2+1
6akSoB3r5K5mZ6xC3w5TFsWk3X7g21tdLC6kxucNqQ/KXnJjl85y1HvWtfmrhZP97fcAt8qendek
Sv70JA3abhPuL4At1VhsW0xN5cjpr8BG8mhwckvZjAvX5YDplKVVGREWKgzAgOEREj5sX9XbgzlB
vE0niugcAnrmrxDfdOGkcDf+UN15nhMSgEbAlILOIerCQL8ZAjYb49n7UrKi4tIj+6N39UBYOkZy
aSDdQB3ynFITChoD6KAdxS4DKmtGB7T/aLqWLz8Mx9AJ543w1VG+Z+tn9tRpNLuS89RjRlv6wmXw
vWXCeTw9+eAWXRaAbV8EzibVhFhDREgCZoy/hsGMOWeyuPBL/jbS1Gd+EH7pQG1eTKOyJj0BX6D4
ZGnFsgE+nfG4BBl8P8Qi1ixQjKjgUGRZyB5233J3py4oZTqZOK4K9RSbU91V1LeNTFNbVTQ2OqLn
E4pfAAHfjnnrGHcLM1sPtxQpcyB8WFjAhY/YiwWxW3uGFrcXSmBjcjNC53xMu/6S697GaappQBqY
c/mS+EZKla62FUCK0dX4/ULgI+hZAw44MH1lcncKU3hoCfznZ1xC3sMXkqvb0UB8l5gN2vwWQyRq
yGfKcM6Rm+HSfo15zDcSKCjxf9Nsp1PnYphbs5AV2cMLA5BgRsaLJ3/eSxqj6918TpA6V3YVjs4w
W9PiQ/bRnF1QU3HKHJqHuWipaUwh5le8TmIAwcDN9LEtCaszL43A5fBGaL+f1ILOGjasgIH1SMvN
AghiM29MqkXq8PSX6qyB9Ic4gRN62sRrAKdODjWmPyLH1YjwFs0KQJvWrJCkdZxTDcBYHG68Qpmn
a94OluEuN3a09Mnyi0N3wL+xw1pB7MMifcGbwZNmNDIFiTKvlz3H5SyDlgYGBaj0W5vaUBgobwlj
0/gRfYZ14nnsAax5ftwB6yRkg35kzZgnXBj0KOE6Hv2jOGA/EMydkLv6zn1himjXoWh9EJOBmZzm
TcP9ji1ig16c1p2OF20Cxj+KKyiwQ6Wx3wRTXRZBnLG9XkZw/zXYapH5/4jK1l2r9y2K7lQUvfbi
23+AxVgCAc6Ik7HzcShjHMKn5gh4euQVFTGaBPajbQLH1lZk7YVLxjxEioqcOYW44B/7j7P1rTcr
QVsRhpL8UFLPLtOnj3e70C7cA4r4PR0EXLr9N8rVZDzs+nhRKjEqDXNzk+DJsOdKLI5Cp5exlhEJ
K9N9Ro6PaBV+qabrF97CaZGPdwyKGrai1LURNC6B1OsDAuaGXu/Ke8X1Po8FjQIOte1nyQt69ZEz
xrEoLP977fvMOvbK6tYmCEZ6XONIfx0y9yYvQazdP2qIyH9E5/RENCwMXDeYHbMbiAiTSNePh84A
IjjLMgiDStgtUYTM5eS28CettwiBLzD6ZjOAthlouQqXxDCic0fpV+rfSxix6S8rYlcIeMz+rUT9
f+Cv63kdCkqXtVr5Y3TctkErLMHBe4E6OxLKbY/a2Fgqm+S9vCe3wFxOKUKHeIUpuYQrBgM6/mUq
6V+oxGXCFSUB3HkCD2CuXjC79mJVjiS7DiLT4Klgkr1FS9ymluy7IJTbwM9htslfNgKaC+06DXZM
En4QlvT5MQej0yce6rCHufjiBJ3Fk9QGFbzVg9324NK14rOj9QOXUtR7bN+etSECJuWAup6IR4Wu
r+5Oa14lt9/BL7IXIIyr/98e12x5kxzHsZNZf1SHJ3xkB3aZP0rIhX1hXAiVVM8w95rptllN1mjt
M5NCRkWKo2L4dkfAdW709EHlRx/lcFSnfCgUkmm+3RPJIDqDmBWaG2Ud705hpp+wYoy5WvIBdDKT
Wrluigi3YjvpcFWw6cWGWYIj8EiKFTBB4lJBcgZSp/NjjwqKyf8+DS4A3/LPDjWWac/mbX7x9fnV
Gxw+m6KHaBRZP2CIp6pNt8oURkyPeRUtP6OB/7zChiiwaamn9q1KE/WeVaQYEQO84cl6QCJ+KYRM
eAGbMonRUbcLgJIIFeTwU6J6fHgqOc3cpbYNGAuVRmuFUfkrAhABwHmai1CILJPfe3uDsMjEzgwQ
ogkV6A25qpwgpRgnkC8pXGl4Y4iYB/9qOUo56LIH6I8OntCm0GmUWBQEMOH2gihv8rVoKZWEUmFr
cglVitkpQd9zwQOuarpVAXv1uXakJGiILhyGT6eQdtMOFPnxvzS5/SMkch1XytbjAb6KCe0dkkQQ
tZW/baH31EUIoJILAk4IcDF49Umk/OVex2HFfzNdws3tD7qu7busrYMQAllcohJRRxVh6JWqKgyG
a8NvX+UnbNmJYSvTDDCgXZzfQcw1SUZL0kfJtSUzdTYhpedths4scM4KadPZCLobQMqtfqM1qwFe
EgOr/b32UK1Nu6KNgPz1zwh1O2+FCW1B41pDTdCqlZqWO7YowxOPXIek1Gam5Ub8wqyxJUb0R4+E
nQkSV0xSmmRTrNOP1TM1WQcLbkPdnolUvVs7vrMCjbCyB3juihVdGFWe7bFbMzJ8+KV8DSB96T5y
BeH05p5qhD56ck/1zvf3OT9irUkxwn4jlbhWtrcVPEg8OB4Owf8XBesf/ZQB2b5/Yic8LyQ5SePr
NyucihDrspc9uzQKvSonU7syIXWyq1GhUE2zKYt5LQvfrz534PLndDLRrn1ofad4Wc+SKjOiY4XK
wkcDR7dBrcvNL81T1u+2bUGJ2CosJlXr/3s9uRWBLZ8DF1iPNYxs+IFEUF+1dnkDo7p3fwspB/B4
cs7eD0ObEU6LRMvv4J61g1y1s2gFMHscgATsQaPatufGCe8Wm5QOeo7lhJVkDFid/PezGlF3p0vH
8h5HpX+CGL04yBDz4ttXfXQsUrIhqvWA6I7RC7LyKyBiWf5XhSnz1e5w/d2IznbOCPzgbJpjErmh
iyBo6HGr/1gYQ+Q4/jGtXR7r9IYNzTJreo5RCPYBzOZDbgTS/AsIs5SU5v+G34jT7luuy20WyMbC
GGI8IXdyFbYNe8UtuS2DsG2mOG2eMowUmVfDVGWSaBw+V+GV218huuEE0BLGXR1uUKdI/8wRZaLA
M7QzvLS4lTLZIKUGxusFF0y1Ij7DRvJoRFWURHHYvDvPPnNnBw3XUUq5lvbqFKaYu6p5JtcVxLk/
gOJ3g309Xcz4WaXrSQfri/87r18nCJ8ey0/1FSxV0Y5/e0TGuH26VYU46fUYRlO7pGalHARm2CyP
UH4Me38RNKBQmsudfg6S5i9ozVCpJ1LtDsoF5aoKNM4L0zhhJkngcSmTHXI7nM/viM9x9EIZ+zZw
760+fZLIkRv7mQkNe0rFegFLE2dZty6gMj6PM2BREssGkBybSk5pzA6VICFulXtJfQpeiPR+18q6
6X9/fHYvUVnydG7i/7fELmXxwhXN9bTmuGVuJXnqmlno5J5p3kUPa1Ghcw52alnhW5COWD3suXOO
pbq1A1Xw1U9RtkHFZ5KMmuQI1jxbwO8AQyFUFv6G6kYByMIzUheMEWNUJ+1Umts9Noz3IitVco3U
K9osH/joHdWg5vDgmjWvkCkFNt1YYNPKXW1ohIgCVmXHxOvOKoYivqrYDj9GoK8zvbQHFw3r8PsB
vDgStdmKbYY5oKmB+hQ7c30lbwVCl2rtq+u5K7L5t7YGdlvFf33BPeaZvxysZDioX0pD9xD5xcaP
Z0MZhSQkfSBsGCcjBC462fr5e1SjqW5Y7pzDFkfThvyma2/3Q4DEeVD/093pRLtJgFwqJeG7Wl/z
49HWIpg2FFg46cCZRFdZYzU1VUiKwqPO9opO+4b/Keq3zgXmab3qMW5nxQH2x7pFjl1jAuggiBUy
L3nGPPmQI8+70Tswpd3gYXWYgyYkySk++XQiKllBBEjtE5tKCnuqZ8UKZYj8AbJGgZRf78TF9w9w
j71koRlOfB3t4D4oa+eLbkQEPu1oQv2ap86eEvgdgrY+gy3++2Oh57lmor6EE7so5kDvDbFwLNIK
iE+Pw1oCQjcO3b2xk8bwxJbAWXEc2xLaNRwUifiNu9bzUpikRFMy7EZOH9gCUhCo6iYFbJqBmfGS
lddyS9EAlRnP7sOnOeCn2klCyvQE+1dxwRrQH+8oIFWoss7Ea/V4v+YJR0VZ+oe+fcwJqYynd3rK
D5NLGeRVbeJ/vCOMiljVqgT9xDqbwWzwPvvSnt0M0/E049Abn4L08rek8TJl+xa9SAv6Kt7Klh12
Fm5ZZ8HyhrQLFkybzX9+fXOGQN1+hAciL/nP4+qKLGES+plRiDpkXdf7QcwseLuQSyMALeY1X7HM
ab3gAlctp2sKBCf18gdPgULVdxG5TbEkhokEPl/VbGY6pvQaqq2du2XFadm7R2eskJQfI/UuCNRp
9wKmojkPaI5DbFxldh3GkSuGvW2TBZaBcBa0JKwfhFhyZdeieA60dh/7tv7ZIgd6mDy7CoQ57Tz5
iZD1yW1DDZrounxF98bUUDknV2C+XkyBf5+13WosnadDgrGmnG2Z6f0vf7MkMgxGmVnNmb52zE4i
xc/xGG4tzuHbtlVye6BtZvM4hn2pCl/LzFQhvtMIzPpm02dtZ+m2Ng5s8p/YIgJoX2Tp1J+P7xcS
W16dJECzhCo2WnWwG4nrzaKxgSPgRip5lKRQEjCZM9+ex7Dm+HEPNHERwXpe7yBgvKncwCmrl5Dl
cM0HmfF/TjxVtsRrHrbOhZ5qk5XLDqYsM5obQI2ju+WiVaF/RtxR4NdVn22pPURYbF5vEISvX5b9
hMquzc3DlWgHgwrXW4UDwIcnrYG44QXEIjO6hkjhp7ItwIYJ3wUB3eS1XN+MuCibJdPRupt6P3Th
O3MSxitViRr62w2ST6Ycg+HV2uZtZkwCPue4aI6Gej+XcAS2USDNMylP9/TDNHTUK5qynpdhy+2o
8WxwH1IL1McPdAR6YCKrRnKAA+Ozsb8hW6w12INy7KoCARW2KbwP2rxu8b6aflZ4fVHiYtN/swtt
2wkebhJLrilvktuVIK2CqX47KlJ149GIUxlGxNeyWqehItdCF1Q/rYoY7wCjFGlVwkWZ8nGhECa7
tMM9mUWjPGMUFG4g+ZaoJTEnAb8gxlmu586HpHpXlZNbX9Nb7vG483m60gMakkb5fZ3ry4SJFMT+
8lkFJQXi9USP5UhzQXmNTSRJrpV72ujuVDXnLXbc7pLoTi262X2PlMt1NNumjrWFt+oo/UFlDa1E
HHPib/enOmufi/MqlnF4CFptT2xh5LvNTHZwXmIU02vovHUEFLT1V9e2JXlrXwvwh0xrs+YYJ6sQ
vHzYG5yRtxhsF1FY+FUlMS7lujzAUErkMMsvLdWCUIiKOTIKOEaMVClqFK7aA4bCsGN7VVBfh5ez
v4gcrhHv3iRnGPYwfSwElRyG3z9iNVC/68aCIf/MJ+l2an9HPKprEvBplx0TNv1ZkH+9P22c56cC
TIwTI4vxPKFgFwZMJl3Gjo235LviDPRu7AR1x5sPuYtzpg6glfmqA/8pUkcuI8f1QyNtZS8AmlKU
Lqm/tllf/b7Z4VV0vD9kSe9ZZ4kJwPnh4PpE3JovQ1gUYiV9/ZjKbqd40HfFStuWRJ7XS8VFBA9O
2aljMlq79c9fGg4NL2xU4bbwn5PambBMGVy3xVOuIG+PXaw1EzJoUkZyufOAO5qinuihoDgMBNHe
syZOsWzTR/DAnRNvS/GNWUKCHin8Jknpi425KTUZotsPpkEkUai+192NkT4ZOlvcodUeRtJH9W6u
ZuDahpKE/9bbH19uSnrtB3MS6aV4AnQ0xdCSkKqqg4xlHyu1yiRnzQJBk6GSAv7o8AB5m2LW62Bu
H+V0TP3V1xXpHYBqukmsfxl33JtRI25JX3j1vi/wNWuowhZE7oZqcUNF7Fht5T0ui1qiq03Rk30I
pz3vc3qVIlcnVHOx70TScqTvv3YEWw4M0Go2tBUA4+d4iLmKY1QOUXVv0JX2AYesHDjRnFQ0Wf2R
kuEzzqfBwK+7zM8A+ng6vag+HFBrBA3kxoDDch/I/h1u3pP1rwCKDPsNprVlWMG1l3TCCsLTbib+
BGMxXyDRtcY9oWmPBjS9TlORbMtsoJ2GOeA1a3eU4yxfqjYPSO3Sxlul+2hsgVBbET5OS2p5qesD
pg2VuDwYxtQlQpYkIqwO41gzGp+tLVtDfm7oYjljO75Fsfm65GR8tV9K4HiAfy/z4O1QaIDIcOWv
8fNNfbip6kQn5bipboGbzx8PXwkbMyGhbZhAb16OwPF9CQ3f9+VIBzmv/j22ZXpTLny+iLcV2seO
Cw6Ixt9aamH4XBNNtjKw3V1j7GvQWK9GJ0uz2sV5h6Mc79MTLI8rECve/4VEd2WeBVgDbxuPgNWW
RqalfZeDh3Xxyfhrrx7e4ZEXsSNLLTkU8gfgigusfDVjxKzZq4hv8kR8so9FUJlDQW6cdSHQLwmW
+oerZBKZ50zLK71Qe9hmY4agy/euDRPUjDv0Pl/0vThv9PwYH+xiqTFxsmPIE8S5FcyyL5tA/5IM
wcoxaXc7Y4A9HMO8WBdE0FCDYGcSUwkuM6tBXQwi+8u5U5y4Hm0g1jR8BtP7TwS65d6ag/G7cgZX
oi+4SFHSoxrEty8eUt8MqhsMnlpqa5sAUbjWnByG0tlafzxG4lCYJhTErQ1Rq0M6rQSSdQ2axhPV
X7/ImdtbSLphPEmvdiDAaMLJ2dds4euv2knQgEuFxGU22fO989X5dzxRzPAvk0Zj6KmTn/Y2mAv3
gtNxezgiWIHVYQ0oKmC6SgYNuoq1neY+M7UURx+QWqjH4ZVeU/HItuB8c8VM0QKOCVMbHvMGKOkO
x8Km/nHe23xBOEb+BtkcKZiPn/fOYiz7lClO76vXKZy6+8bl6wj8XSr4su7SOUKpfLPYDNICPfOh
zli4F1z0tVEzOreudhHPeYizqTgdDMgSrC8h5IQLQDxepK/Ofhbuhx+1p+5R+MYgvKIS3UC85JLn
b/I1638cDgoTS/gHOOPoB/M4jcrVX5YiFnb12f577KStg7jQAOC5UW++3014ymOlK600EleUlSyO
9kcnCqKPk2EEeIQpMTGH+nU2JV0QK7cNQ5SHoUYzY/TSup7LIqBGZjoq/q952lABARTCtExUqdOI
KO4bUL2hcAQbYVPmqf8geS2KoYzVPYS78qXClPkbxq1SxUeku4kwDr9JjDRSttpVgk2FK8k1w38j
JAGhSPw9Mu525k6v41jC7BpBXz9h8ewDs3cvdFyvYNJ1xe+OBih6GaAlUh9v8KrHEjrky9IsT/i0
Fiqi4z78L+jpkr/Ahq+bs3v1A/A7LPhKw3V2m0IyX39w1Q33hXHnVE2KXaVt00xcNQOlfGLmMcmN
oRS/aiXBmZ7ahRRmbCRTRM7ZsotDTcC5apAylD4opH6LFpcpVf+83Qpmon04hXkoa7aKxQHPyoPz
QKQ1Gq3vqAwrDCm7mkd+YjoLkXLzHzY8iJ/4Guhz3lE52sDJ1GHyBLzLozQQObZtxYCxLGiJA4Ds
hwrZbX/NlmfhpMkujbHTU9uFgbxPOwlwqrZILpgM9RsFVVdDSG76ouj0SB+B20nw8ma7pNtBR7Ri
2Yvrmk+jxXdrzBKwOw2+FTqW7SxsRADIIve/BCfhS0CFOd39Y9x2Z2G1MDkdssXaSSzaGXqrcOyj
hnor7/hKLwS7j4Yzvfvuo/jHmwtWFdLdMS6pLfvkiZ2L8OgiAfInD5PA73hnfNlf0cX7sxyJmxzD
sjTvMlLIzsVtFeVmQdMU+5bAtMsAfctxAE56cjdlojOcOVN7ZFYJuaYxJXCCFf5PUq/0XhE01bIA
TTPBcqjHKWwY3PinfI29fD+t7xH/YO/v/z79tE4lpzWiclks1CTt1XwGmyU++fHvydVVlpGf2AJO
bN7BUqK0zxaNMUxLvMjnAZ0g+0tfb8ODLppJKTqkyusgND0DOSVQUFA1E6KSH7UGWGfXM9/mURCz
6JukxS7iCwlnFtxiBFf4YUEsiDfXBWTO1zRG3s3BLycO/Kpv/nANlzmXyqnfmvncWnTZthYCG8yh
PKXUy83iaZ+486jT3MCdy225+o90Ms40ozKDDlDiftA/A+Mp9H5NoDy5z8+4SZB1LD8goDu+N/T6
xrwsfuWc9z3rAutNB5XioT6tKGzW4eSZisE85TcXr16CsllZfO4xN2a74EHD+YyGE4qXSNe7xfWZ
ob7pBHobkR/Ede3wOAIMaiXcTAxgQxt67ADV6SMjsH9/ZHdV4PxcCBD1CswoUX96if2rRyEcTOHH
1qxzs0vmHmyiLzZeGzbpGX9ZUt2SrUNkLXWGmuV3hZDyjQjPPsWkJ7RIWq2Xub7RdP2leWbfu09O
g6Uh1HNy4EKwhu9NViZ3Cg/bts2i7OqbAJnx+bug+mzapQWllgi2B1CHeNYgyOWpDvIg+CIWJBrk
mKuGAhU1bz4xQZ16pdbYRHOYlU7LAJMx2D5rDvZ9ZCAfBofX9OpBBW7RhmSA+WBBe5102CW+vCA7
jvcqGJRk+4uiNVBJzMcAhWmSpRKEfHYsgPB7f76w3a69xDfrNcO1+LIiC1NTnpw5NEHYV0J5q2CB
wEJmmPBs9hfxpLo0gHP3eqnQvhL7DnOz24ln5h06IRH3N+/ew3IPReSy+mQqGDZ7uXc6b1L+lRKX
VLD3BWKykXE3M4QEd0nI0QOo7+IcdSHuH3VF5KdqjJQ3KXxHukNT5DYhY8KnUHlmPrtUhO/dA87G
TDZ/AGwS7yh/lpnmGf4EVUM7PD+7fascDht0PDgeo1LrPMoS4wKCBIwQRIX7pNJl+MKaisW4TU95
pQQssepkdL0rRvXCM4tdNHBK89nYaM+qq1+2skbTI5dXABVx6RVSQdLK4DaH/vn3O9tWC6XZYo4H
sMV9NUs4Mkf5esyUSFIkUtkU7OAWro/Jf+4t+nJK97zqQV1yy3iKSEppMqfg4xKxOHFQqdXfEtzE
7ydVNOYe0MHk1iMeFIrtlrXNJj2yFNyPr8SZGcENpuBt6PGlw6lQcLpfQAJ7gefJXd+hzNrivNAX
tYPNz+QbcjFNbmhOp8VjrLoZiLPoQ5rvG66D59atycmlzXa9D3qox1GXu+/M9W0XSWOJNgcmeDsG
vZ8cFXE0J74taH4udANYVoUI2yPH6C+63/0IfNRVW6AB64p5Gq2ciYpEWehmuiNqJvk0Eu8OVBXY
Gfcu2McWWyyOCBLIHXxZzFbDtOJF6tbCkglYfGM2vUk6AoZnlqaErl+QzqfWxjTsS4snqO3DQ2Xk
3EhSyJdXQv5nvruV0tZODl4KOTW4W17hjwe4nRJ5EcYkQGATa3r7apkGgi/8XDarfQSG9/0iqtjK
3YesH6YDIjI7vr9IqJPpn17QgUSAY7GFZzf5G9G5esWIz5eTehA8R/MRYYL0ynvwuTyQU5kQWG73
84+ZXlmZV0AFN6x130fHG0Coqgds/EwKx7CgwwXQQEGpX+uGJPNQbrNqxPtYVz62m6JcFwbTYb5G
xasENjQY0g8thPqJbRwlio5m4x01YUftxpXC6+BuKkML6/VwkwD4rMeWm4APzPMohUIwEDcOC4HC
bXRpoknpedLhgz65JSszGCq6st0sf4Yy0CWunz6Gxxk7mPLr/W1WIhwxPlACWhnK7/teHH1h9n86
N3QBcVlh484z6yGAHZJt035ffuocJQmlQVYMS0OSnWT0xGAd/Ul83ci7lnCg1QFMG5LcQiT4/RDH
f1/ZhP8lW4xHyEdeR7mUw1w0MCf82f0USl6gVCnT26QpAj/wvBRM10KDLOfqtqzp0Xiw3+JeCR2a
1/32+lzvnnaNwi3lc3CuiFqQjkciKTvRJFNh0/MrGie+aCkjwxpVVaNMD6ju2GaN0Zt6mP2xZQPB
RL6RLLLW+GN4aRoN2VLX/AHSU/ipl5jN9jvv6tkBQII2rH+oRGFPfINAALGmSZRewwO9MshEXPis
yoZUeofA+iXDHD1NVciS8lqM0+rdMy59UvpV2Ly4uL9kH28f5GWUsJlNlJsQx8QsBOD0oGXoTJzL
GSRMNnyHPUDI0BR+8LaVaOv1TFFl8+yusERBDpzeFv29xTJvSeLH99djuOP/b5QkFPru9IFE9FhU
b4uUUW0ZZuxe9t8qowG/qSRLvH5oRiy/xdCNsy0echxiXDv74K3/PeBmxamkEZMpBW9iNsTgvPv0
77DsSsRCckXKLMJMMSmsQOHA0OVapPMNl7KkhzcGpN2hfQ45i5WIOtEjBowolAcRDxlQcKKGsqvV
dpAd1GYnnktELze7BITLp6HC9wyH/4unvmkKCccxU5NNPLNqy6/errHpwmub/as+lVe8yb7BnJmD
ZEmciu9jFQ54Gpz/F1hnwqvqSq8tILzfdcm/Eb1Y80P+FaHp0XBzriDQo8GIl/5fBiV9dd/t/csl
igbQDxOzZsQwrGeU2uHo4iLxQ+etRseVCmgPt+PHfltMz1rE83wJOX9jpRUNiYJXOVu3ICEjHYI9
6jHVMwestx3Y6EU2jmjYugOTM+TgB5eytmbx0kss1XBxu5kvTI9loo72BCpvHvU/vQoSY1kP8gnL
Dk/JImblp17Y1lmpvdYmrp9wG6DEf8k28ltN5FgJ3qJ0a0hqVIPCxeQi3BLD9f6kH44PbPmSccdK
SHz0BUmEkNYzmRiXCji3V8oqM1MfbMDszUemhoVJq7t6O4fkusI9WF5VNBX7NIDcjLcKVy2GIzJC
Ni9K4b4CKYe45QRedu/yD1OL1SV9V1fJwVxckD6C0kr8WaTBK2s0u5OubUV2N29Flt3gDpcYf1mO
BMfCX2y61/z9gryP+Z7BZryfxfWniLp+Q/MxeFNfX30nnKShsRDFfJKNSyAi5xpFtKIVi6LT2VGE
yEF7yb6yG74IufDu3Fj+nHSQTEwsNbEp4A2QsTsEJmzE8rC81ZcOHjcFeO86cp1ULi01SBE5shOc
ABy9DEp8f6MCZ2h2lcvgLJtPDFRb3FXUKrpo7qTehQ5YhxNfnJfYiiCG8ktz4626/tb7at7rIrkl
P4ujhuicqk4hsGkv+8wLzDo6VSufAERoclLRb+g7W0GfV521QOqEb1BvH3ErB6H9+K0DIIHj1Jvk
rVjgMOlf2NrQqLGj6NlkYB5Xvi0VAk19JW0Blld6mQ9qTJTLRh0WNwGM6EnGHafaz6pW5LJeAww+
frrYAcDS5SKjXJ+wpTRuI+3Q+HhNSlxUU0hDlHXrzzb8odpTxf7+kUjdHs2fqdcn48afSb/zM+3n
xzkfF8oDz4ULwQBm/2mwkWZWmYuWSDsYYK+AiwmWdMlVpO4LmAZm5TNRMA9KRBCC2YHYNFgIoAO4
BomLuRgNN+i8BcfEdogaR7TRxJ2A0UuWSYokewybadhVNv8hM9d6iIlOgmaahL0RfZPfyKUleFmz
JarEacEdlhaiPWSYfOFSk5dTgcNJY19hPjBSPLXVKPcQcRoBKGTILFfdRCgvuVYsJHQ5FuB3k5zu
OWkEl74rSltt5Vzq8sJtTJ7RbesyBf+O/zotsH8dsw787NvYsBaYhTPP3Fq2/02X4Hrc+nN2oAJB
gpChbciy0VjdTIlW3Fp0464YjBB3Ok1vA/DVVfJi5X+lAIUR55PwpJX+FEgNsHoiDARd7ouX7vA2
4ercBg3WC2zJksDa6mUZK2CyZKf53wfw1TFxTm1Qg/luspj95tnkt+Q52wM8ew96fKpQUITTlLo9
QBc9sF9GD4Ly27uac/J+zXAIa7apIORvZfFe6OZ5+YFZ6XAqC82K8rCZT44TvnJ0snTOj+YqG7JX
muEVCfwo7kg1JVjE6JJaBx5WGHHH30V4qmCaeXmoIVvNdVMORUbo45Jf/hV60/RWCHbMvHoJ/hcC
TTuaHlvQQDBuheSRMSOnw+zliLerS1ScHQ/qiR7s5mJyhay7LHoGV+JuQzPm61dXFgtfnQg4dWMs
ucW54rroibqMXWQodhs3SF6dyfHWMpMpZ0RxDlG4fcVNFv83IdBatEKlrKZvsts5Qzin/PhdW7Yp
xWIubHYwD3/l6t02M7iSOQMjFfvSLzSEZKZAoQMwjHCLSw6VcQONXa0B01MWECdddN6b6zeAVURk
B/EBLK5ZTInUgNfjB6ix3JGS4Tf79FHgjZL335mIW58gJe5fWlUegK1ZUpXy97ZvP7p+la9aBYbT
CZwKFOpWYy99PwB/mwbr2LDrayD10ILpxWbMkA4KRxgmeti6WXSsy3Z49e+3297bZO4K23NlJqEC
Lyhv42t/aXaJW67ndOGEY1mnVMqC8vsjGqwIMbKQhhjKe/BLhRoAtz8qRkGz9CC2g6m0j7qW5i/t
1BAjnlqJ2eBduVZXIRD7V6P8FbK4q2EP09vAR6efcXGvg5nInviDnysUdN3z4YUqCYkH3vxos/Le
Bb/VtPx8yARUDhxjK+OaKWORh7qnys0Gs3weVNjJ6InYWCCZ59zq2szsS+wIacCSG3NGKdCgngzT
zZ+/nkR8U45cwjJswqoN8ZUyE+iHDabwvbAO/1wAI4ZdE1bHY1XQ+idlMkiClUABWXaDgV7ZnSDP
YV3A11jN2gzYwMaaQ5iAs2Lk/P5IXk5Ksm10sVnytvsSw2iy1n/b0sVZRxG+mSfR5Tu3DJnadu/y
9xkgZUUQPrF+Ng8wJfv8K0h4wSIjmvzxqQvHUkvyBqIMBrXLOz6Na2M0KiIKkluOC8y8D9W2frQC
GX2JGh63bRSbXaTezYeFsbhe8l0aR2OKztGCzGTlLoIefLvN2fD2X5MQ/Uz1n+yh9ympog700LfX
hw7PP3U3lGZ/plbmzUCypGTcSvnrdc/wpVde9imbTeUbKlsvF+9Vo5bz/9pxDuzJUtkQ/K31iB0V
9UVmH3JhrbUz8k66Smx6E+NmGH4jXQqNxSap8biVTZhBFx9+ylz2W6HadecuTo1uHg0Ni6koGDmv
AXQfxz9QMeypHeYFPfex42RgjGILPc08GAY7lCCBVcK7VHuX9VJJSxvjSwe373zn8cwoi+1IVZXP
hkqtMCmOF70PpfaGDXOzZe61VKy1M7LdNSnFxwaWjTY7mvABVm5l0YwiOhmJ2H0zIhaJwsxoNiD4
C8Z6yoKCvAaJGcIXKh4werCaOSKSoumiqAmzD1+ztkJsxTqcnqvT/hZ53G7cHjnLltghSN4sicgR
Gdi13uNNOaF/xkQ4mqcxPneR6kNKjcnZF2c0u65jP34jhFZ7dXQTHrWTXeTRrZrK3ejuG8Bk7OmF
GapFXGXHhMu09yfxlmRT3TMq389gHPdCfhZar7jy0eyoFvSag+yhUPHUxs9VMIUkuf0dAbtN3ak1
np6/Yz7aE59YAgcODusvJ8DEFx8YVWIKzdkVZl0kV7mF4uHoWYz8GRZyFeLTbw+KX+4/pjaFxKJm
XiinQ8STbZfqVsa1jxU32FCbsPTS+ltazyi9RYGYA7bZmB48E9TXxz4wKB0xUPga0zfxWmVviFec
8rFVjy2PAQgR/T1F1rI16lG8SzZ/BuEoHY9K99NkQ0wUfb/leMwdxICtZgaDhmNmEo9No0ouhzD4
4rVvpHNpzfGb4r078umDRo5z2jX1n7wVYfTqdblWOM4MM7P9eMTTayLID84NB+7t6g2iWwLS24UJ
4DtEfnehPPFRStH66KKsLpXqHRLWaEWi2wrBztpNfgyEYCzch6pjjvX0ZmXZr2CfWEJYwzmddmrA
/s62HFVBiH/deFD7+hhDWABL6FoH0CvUYH/0w9XI//ra9lgskgFkSEeJcO3aWIx5ljv0onr5/GSt
XvQqpUB15eccsXs08XuRRh9mXtjtJx5baJn33wR89/UJchUqH4r9iCRGyrCA2NkQr3Lb3cAiyzw0
Z+lr6v9DxWMGsf9BorUkoPYSc0xnnz/qg4f32kTDMoQtv9C4izwHHTmpXccN2+Q5TV3FlWnwkJnx
uzyHC5w3aG0lybss15vKQPsVSl+bDJbwuKhJEhdWW0XZzDTFZDzbiZFmrRWk5XrPsqAbYHzlucJE
hrGQMUMwlSLVIAGBPlV9/YEQywK0EspKBHZ8YTXUkbtSBNPsq+CGXQ0JDfU+4WC/l7d9QXUaI7cV
ben/sj3xsAGTvgMTAZAhjyRkcn1N9EuE3htZrVuCQJB3lbBHFaUKK4KB2q9RAT+6xj7Q0FuMs7lR
RqmHyOQX3//OOC6de6jS2WRzKNFXdGkiMvJTFcCu3rrWqWk9bfOCXQsPc7VGrVPTXVFx4M4l+6Q3
k6Zo/Ul7Z9YCERiz9uNMzMRfUB1vItJHduZqY1nBOpubDxIU6Kupb5v7f3+Z0N4+3hrbO/hslhKd
f2mpQwqgI4ONjzuFz9fmGLh5jyiopBU9Kv1s/ag1Mn1qloRJlMVZotmQ2kZZcpMfWeOL8CZKA8nt
Cct0BJM7DWk3GY/NuSEvaO1iLVP7d3gH6Knlmqmc4w2ue+/gCSHEjBlUVrqOgYhzeEsq0kfXJ2Ho
S43n6e5AglDpuDszXJiYzizrMYGyUq6Y7ysSMxaAOJBhiVH1yYIYTBS3Gevxkv3SQR+LyISHEo9y
ZL8XMKQxUBtao/eZe4rZW5e6JdeSwF71V1CVgOfHjXJYDz99WN04Gyr//KizCHolCd7ntK4QyiMC
XnFfSErrJEdnOvg4LMmDd9GnNw3OjpiFLTJgfhmKD0l1ji08XFkS3Pm+G0Z4RQPRLXtLfAxSiwcF
4ELLsj7w553nmgRyuqCVE/JO6bOdyfF7ldtXKsxWEXdtBMfG2T4hreCIG5PorZYvPYbokFSL4G/j
4Va5zXDA2GU6mlRIjyuhh9uYM8nwtQeznPcA9l54C5S2c3vCLN8y0WxBirX8gHCw6Zyf7meK8MQD
OoWHP0VFh5xcmHiesUAxZEMNWp9CUij6Iv5CH2d8klii29yzlN0GvIHsyCFhHKjX1ou/t5DP+jTh
b2g5PGMDzl/gpMomLDIoQFUlG1x3V8Y7sn8qckHRVcFvcCSPhIowxMg5ak06Wa/0Lk54PN0/zADH
8pFzuHV68VGbwACLcqy2/Ikni77+ftbpVv5ouOEMJ3hc8/azA+BUwgj8frWFFOtpKK5eutQKfQpI
CdAMnaOy6EkICRwLJzRKu7eH9Gvugvs35/pIRXdEAb4cm3B4b8L32N8eNEqFC+wjv22CMskHeTBu
8L8QtvIy1/KyjpM6U02QzFLMNcqD/X8huhCn8rpEBZ40airJzG6Ha4dyQrfUfobtlGiB4wcAWPsY
i4idgex/bLX+Qdw+EqYsZd2KpxnU7Xxj4p90hj/gdmnDq+O1xPpuBT0ysdyrG2oKTEvoiUQgfq8G
Eqf2hvRdslq3gFTQ6NZ8nKlRSUYu0oCsF98v+bhAoq1CAWnnh2sBl7FuYzR5uk5TmAQcN7qKpQrc
yNnzUL4aAL8ytESM065z7VsPryMvnygmdLQ3BOddEPX0oNUORSuRtUbPwDbsZHNA7PIQSkxW1l2d
T2X8+7bixWWHOjZ15pTyzhcMCMzxb3RKD+jW6zbp01zzZuAV7BN7K7M5gTLxKUO9bJ392KXdFrIV
c3mDJ7PzscO+jGfuqurXVmC3HDA6nA829FBs6kKuG7LPq74Xif1APDTa+ZdZ/8q75d0scXUBIZu7
SsZbL2qVwHnReQ+cgtnlx7DlGNA3xZn/eEAm/KwqstK+qJx4RVPLQt8K3AqhnYkJZ9r6cjdr21F7
MNzoL7MdkUzCXLGl7EFdDkE3w53W4yylwExjpvcZbiHZoUHdzup4ymMCy4ibAmh5WVx4XWP0WEA7
Zh29PCynXbp8IAGwIX16cp66M8XnKm4rkJ0V+6hs8sMppXQQfERf59ftUi2p/oXrrGYXd49KVUM4
xqbT1rNyEY0NWz9PLoiAD63kp8iYeo4XxyF62+Bxrfwz7b1yfzskaF3GsFw+NNn6/QPX8F2JQ2p4
AeqxG6mZ6C7AJ2eQA/v0YZzfCMSqzx4FPeCqgr2fIfloQp1DHyOye/EXrw1fDhpti35nsyeZbpTt
bpGqtvuwLhWqPqrKvk5CZ6qNtRskPcAQlkyumOArVPNRLp/4Nn0TB8uXAEIKqXaKiQk9bUVsxak8
tPbLl6WDVcdqaptLEeKjXLz1c+DgW1WX1nAycLvzUv6VYB+dKaxHtYHve/l1J5hHNz7DDmDn7AMR
GAQ1ax++7NNnp5Y6wGFqWlIJ6JH++e00gvHxTFh6jelUKm6Es0PVaYKrX87jj9lOC4jkwyV4jDo5
1IdJjxOOoROFtI0c+VM3+Z06l52/UaicQ5Sm87vt+0w/on4aH7jMcTwfhAA8p2LXcjGgm+qqSVrS
2Nromuul75ZrI16E6YFL5VjvufIONEJOhgl3Qzu/+Hpns8I/IuRBisEvy7oZ/8JWdo7yFvmExQdD
40cs1oQPAfbKt3srNj1nev0h1a0hNno9O0mha316FME0CuA77QplTXw9KTat9FAgxWE7yies1OAZ
yaYMG40+Ti3Uf/7FkioU5H23Z7c44xqTj6pZS94mhXe+3iOSj1qZvKZjlS35L+h/c02S//fB3Fyh
jc6fbK/i2r1mvqajUNlhP2BwkYpy2FwpdQ7jbY95V8wBriPoQPlIupSc+bWia6/o33glRErIHeM3
W9cTYu6rxPaHRyljrhSma5Dj4pWtlj3d+TqNQhyyq57DmstI2xf5zzWxnPO6rrYixZadp6zoFAD7
el6Arqx1svmc3pKqx8Rd/uY2LBv6dSHAM0v/z7yfg+J7bDGKQ5DliXI+JPaG3kXyyUJQDUAUjztU
9FQphx2aC1iXWZ380Zkhmx6GY8TBH7JyKZR0MQnaQid8doRTF8L/rW4zkeSJVEF8H3uYc3uHekO7
W1C0NCTrf5eGfDKgOt6AjIaDhspD9Xvu5SJwJ5m6IeqmOXWsBVzJRq6C7SEvKHZB4b/pMO6XiTCa
VmhsN8n2SIPrdkvNBRqmqg+FVo9yGfe3Lj3cfFswgp3tVARJRluwYCHuz4XdJxONn0BVkqkh3DLA
mCiiTF2acUNob23PNwY45OaANUALSt1+DjPHvzIg1/aj7aAihZ8t9O1NaF0KFJCJc2rM5SUpnlWl
48obSxmCH0LPh4brM+XzwIvMxd7hwnTKY9e+ZfVPeBDLlf1OyDR5Ot+jD0rOrn7wLKzrqMNoYgy0
e6xbzcrCA0h3fKUvXGkyfvzLlVFZfM9tMAqShqiWJZNranNMA0g5k7ccJ0jZDTQQD7wxV4b0BpVz
H4YEAkFcQMksm9YkH6Oof4cX0NLBhW2a4IhfmXd7HMQFIzDdTPkrnlCN3Hic1nRL29DhIDycngLX
cKDW4YKThpP00DFlNHltqOIGJ4AejCdZnv1cKA9hScNPDd1hntEC9PIVrNqByeM+6Qps2Vm7LUt/
8YjnycyCkKfgVeXyJx733Hy0849q4cyniDyuDh8hjOTGQVbPKz/7UxU1OJ7UG418aaEgsBSNDGCU
0ePlLcupPoJI3Z/9QpCmLa0zwkiB0CENseIDhgs98vYIy2YHaWGDtgQvfvNcWUayzcho6fiVjUAE
97BckJ47QedGoG7hv1248uSxwegAzT73ooQBjXtTBcqSHVriZ3u9KFqUaZ5lCffhglO5Fb3I5zQZ
XsdCNszxiGeZA0VcaO8nYPD0B2vLabURTzlQVz4DEB7WthHivrLecb/ML64N2KLiTuGTKN9gINEO
79O+FSTCbDOq01wKZpahwYIKM85MAzQX4ow+0f6zCCDNsjGYrlO8Iu2L83YyoZYQAeFU699N57Nr
Yjz7o3CogdR/U23QucLjUP933dyalfVdSJY/Q86ExUrgu1wJHN7w9/knZGODLI+Oo6SHm0lK/aKH
bkBlaaz9sWFeQyPLDDKyfgW1kneGKF9Ij0y/FOzUXQsQVDC/taI7rdLI6nhUGVuMWsQ1oRXN/r9U
pdssFFQGc9nuDZQFc4w++p0k4crUwMUlQCSS3TPyX0zszEuz154E0ukwOAZZ00Hj/44LbTFT3F5n
OBYVlulFlD6IUnWaelyVqL7EC107lGsxdysE5g3MlQso5BZjYOMiibnm5ezSN0ReDZBK6FWrqnzY
PpdWd67B331/WlfNHREQunnp6XYeIEcwXsjhpNo6BhjBAa5JhecfW/YD54KytIwnB1sDIHiJQVrG
gVerKujtUt//52m49pzznTt02Oj/A9S0O+Yil+c8Lox8PhbOfDp816nvl3r7TuKYrU1VLvROrHl5
/Hi02uPZeoExnmXfuWULJzlPz+7z+qoHSLSKf68AQOHL6BrfzZA9vcQEixgN4Fm6skJ00LT6EFFP
Q954bwaGLqpfAWhHxr1GqJSPt7DVMjGubAN2tVnGHojD7vK08Suvbru0Xx2oz9vYfBZxT0cJzzkS
Ghe3iFkDsMU7pma98YMP3wetWugztZKgWWZIDCphMbie6a8BKgSjU4hmdtzGb7En2y1mIU3GYzMP
efsyOA3SCrcBOQe8z2XSfWaAV2LLowB0ZPorXFDy/c0NiDFfqmk7kbMddMS3Zehj4n+785czBuWs
v/D7j4fhXqSNuyaIhq6cOpBmghk96jNFJuVhNL4h+cv+PtXqkPXMzbdaCP9H3W9MxZSGOG0PNQs9
sBDJ15+cf0lXOR7/K7w12G/0D7SBNhkqQ5uUj7p6ssGxoyMs4bkWNea7nAUhmfjnyABeVwLBVDl5
I0dOQOTGyRCnWwNA8eiyjXwnbVpKX/lKmV6Tq/noheALu73mYQHzOAmqse+8mXSblTdDn8YdzfQ+
nUCsj8Ps+76eCWDsrNu9UOUcO09TWgdol7zR4ordI2JHK+gkNIjpljyD1hgmmDp7D63vCOJbJpxI
d71s+1fTmO4qZamO03tZSBAXa8PTjXHlBxlMvyZ3YagpvbU5N7q7sf9dq5KwgxvK/F8dpcNcYYuk
//JTekovkWdeR3/yLyVBvBjBHVVfr0WUlYrs5xbyETbv6v9U6uPH8DkkYPjSojIdpAeo7tRCSfwX
/TbqK3S3+fRroGbMpfkKpPwWNvLQ/yuvlvBqqgAGGxZiLmElXfXnkz0kuPqI7ghglhlOhq95iXHX
UPxYqTWYEY7Zyrxov9llDNr2Y5PgqwLVM71++xSK936Q4bUkyHoaKwrqlNFPfZrH5tb+zPpBLWEf
sKE/LBqzRhxbUlgR0jOf4e3ucc37JvwPGXvOLzmMHv7TrT0FCutZEOZUjB86YzBYH2gxlcIUCsg2
HfFKftkknjK4POZiFs6vGFCvwWMYCF9vw+t3jPEWZv5GNMKGaReeClD4u2cvtxDLu+FO7gUpeU7j
uViVUi+qjjDV14ZIVP30bE5mConuOSlnIm9Zm8yTxoWGTUU3qdBmTsw9VM3EaePJwM+61x0hu4zV
dlG+dWFlZxdv00INUvzRYKQmqIMR/JNkYzVILBcTPzt2BGXuoO8LjaK41QNscsv2z0uIcLhPDqa1
hM+wSg/KsIkC0xIFug1Cf33Eq4dB3MdWPmJVnBtRea+E9ET3Wu2EP79RaS+lOzSvrXqm9drkWLpq
aQHNBH5hp9TyvbpAIgh//dhHtlgurzOztpc5CjAVC9wWlCFFV7u/kSMig4tMhfwj9k2PTKSQ9rCA
1bxQ25mJNsLLaiW5eKemRrGF1yMiUHJOntUb33xZlvGC8puY+XXk/dXuwMkpugwrvzVwc2vujSYK
z701IdqMAPwp6/nP0pxOibY1LpbRfzR6JwuQyCeVcHdZmMLlQeqX8qn7ArqAWtE/58tdgUoboHYz
lHc1IKi2FlED3y0tWC8yl//oOi+qZfhPliWmf7XE8bbm1KQNx4LOYVi0AWZAvZgjFmi91vPsuo44
HN6NmyV+ER/h/UNU7WFl/ZMBjpxpuuj2+PujoAoVLm/QP3y9FUV9GRpyVB04FSdPzz1WwVx0VeKI
GInB9TGJqGwfvZNjJzVREkCf3yxK0s0UU5XEIm0YrhGD7MPEm/mvnxaD8L58G58Nx1v+UShV8ZX4
5GKFQg7BbxeaMyFiUlJACZmCxLZ03CD5JVOXbmv88iIq5yzQrPglzZZQjewGxVYRpmui5AdrEWJi
CwxCjI6C3DSzhE4bmyDaruZ7Ne8TlB3Q6ytVZ/aZVVD8tjkoWxcZXKWVsk0XbelRd/JkFOq5aurI
Qthj6OcX3RVn7d7e0AONLGReLZCOt1M/yE4Xai1NJQFN+RNiB0hyuiHM1pROkZm9lW1xmzq0cpef
S5xGgAiuk/4QlG8155pOtoPG3tY3gM/GVOZZCnr/vM0OT7exuhRm9pPbuKL/tD7IHJmTU3tFR/F6
UM6dwj0+69D4kfopfHI1fWvYFbosXVQngJGa1jiuZdXmQzwn5Y3mxav+P0HwsDc4IObSiTABrvhF
WGRVmlnN8skqAE5rYiAFIECG74Um4RFRiDjXcUPt81ZvAkvm+hxv4EJ4d7OuBQetBtUSEyo3nCXo
r/32s9fYnhX53T47kngwRLObqiHq1Fkug8Xs3c5xEokVe8DXRyamWnZDgv0LVsVsDM+p9is0ldyX
ksQiQ868DtIRJG0K09BAWMQzg0FbRfzCEatq8E4G8nNLAK5gZ4JDhAaxfpxWgRYbQGZqs6h5Pi3g
e9yjR08LPJFjGkWxVGGk6GTiQyJhkbGjuhWFqTU4Ra0KokwcZ094AbImzPTz44sGgdQP9fYrYlib
0ioCqMGbYwrAHAGjyx8t0VJkca5L1GE5V3pE8kWIIOxG2qlEKdym6QRZHPXRIUEEbB1p4PRC/B/k
3+MK+hl9kAd3Z4jFvQrR1RozJND53oNabwIT0VYIz16+Si/5MZsWRGJAcFhGzIVQgQ+cljDPgqqg
29FgFubqvcvSYSFwNatc6zSXAJKPk91awAoZa9f/ufNn7sZMjTTWMOUAw872Pb4ASlv9f0YhvDQg
TjdYmzZ4CqVD5HX+qjm5F827StltvH6n1hXCG+oSjQptK5sVBHEpbT+U9bDCIpsBkhI3GhQOGztj
ViYSvKp27KJwVL/mhvSLjEOCXw3J0tSFJS7qtndRbzTBbUJE0CQkFNi+4js3M8XCkE1gfcV7MP7T
ZS9/2sD7/EBcfFat67kbTuvg/YP2JF+bbgy/2wm10dTx8aJQ7aoqusZ1r0/e0Yng/m4Id48dT+lz
7iUt/HsklFpHQRtdqoYt9YNaono6wGSoUr81f1jT40Mmw5yfd93nkoveb6SXZdNrHyskhs912Nj4
TZnJ3dh8l1nKlOs11r6r7GnL0V6tcU2XzxVNbUVIC68dgr5qf5ZQzTqoSYruspH3YPKPmK6okbqt
cHX1VrSRMr4X5Zt60AxX7UyX4FqLLiNfzH/Sa2TK3vXz2yxwSWaxr9o7tnHOWeRNROaL5vpa8lcz
2A4hgJtW7pe0IYdYXBucs1E+NfDJxc/R6Yfgh615eMLcePYM134sQIDcxdxqrjZUaPvIpp59fslq
wlozj9xgnQp05ch7kuMo1Yi3t+hyr5AR/swwiYCTbjXk8prX5BTKEa7ohRc2vjYekP6YEPnC4Pbt
EFzbhoKMUPXG9lxI2u1eVXe8zvhaejw7fYwblESmT9wptrvYw7UuBvbkPWD+AtC7inNK5bmyfKYi
srASsVzedIoLRTVv3n16bSTfXRicdonvCv8KUL6R+EhC6v57tXpcIPTnzy5p3LpFuBmBfKav1PIV
n0tS0ueKM7qHVsoQ+6kgLIebW/Ecn/4PaRRFWGUczu7T00JKA8aykgxhIxIuPriaSSTUVWOi7d+V
ipuzRSJOR3Fywi+BTNB+SjkXxfBgA89AIOd8p60qliYGZthXdDrilgouC1PP7UifASZ+8APLHQB2
v/4sfN9zHeolsL5T210/SdjTA8qeVgQx81SBxlkOz7R+ocPRIovYR4eJKBYuaSZEeCQyfqokWTCQ
MtTpNPK+cspJMT+B7Oy1+F/OaPLmJ9BJnRiPT+pYflv3m/LCsagPrJJoKGY5nq6CCW7tqlz94BeJ
qVskqI7g+Ay8UBDpaqoJaudyASg5LibbPG1lDY2PIv+/4LzzIjli0fanUu23+8LXjrTnMARi/1pJ
09fC2s9gqsz3MWzSEp2dqtM8epW3mWsRWSFHp94T2SJKrbQj4sTbqKMWSAIoPFpZ4vpfwpYdgb6y
Ht8XsTZ4XNOtMgdafVnRNNDrFfXJedQKbZ6XsC4tdYBZIGwBZgdAHqobonSSV6St233bJ9n0cHAj
CcWY/w0JYFXv6O3gn+8u2WBR88juNqGeinZHY/m4p+qyvvVpjkm3cZgHNvrqHTqmhmcT7GLwbapD
khP1ZaUH7MWzz9dwO4JhOiyZpVTDVQMTcqkuwC6J1mH6hSfyqIv9IcUy7mLINW2eJ1o5zsUo9UXg
B3S/3MbBD7QaZFKKyEhf/5HoXaXNAu6fvVuaO1e5wRFxd/A4pRqZJ5jbG7+To7gJYojNfdKdSEfq
nDQ60masYt+EheoqvTRuG7cJnhziM2oRRZk21KAWro5tHEnpC8oRdMLvyHKjmYG4RuA0A1X4YntK
y6dRHGij5CFffiS2jXxB7N0x3BQMhoYNagSM+QqtM5jKAmVbfMlQzpy4W+Ld6i65/4NnQBlKEXlg
KFyjwyK1l5bNL7UO8crzPMs8MCqlEY4ZqFtXe90KKtuM2Q2ldkkH5qmKqe98K8hjdvZ33LQafhxC
yiuhfLMKKqc3h2w9TI7IqGGG4uWE4vkNA4WDpMOInUY7IpMk3rj08zHXs2BkjL4k80VRey2a/UHs
Y060oHU3Iq4ckdgw9ovG4Ukhaaz5KTdyCcP5SQN+/penlxztk4KK5ag9Os7MtBxgczFxAng+iDAX
Bw9gv/Wn6UcO3uwJmT18moC6CIHCA0Ic2HwNzwez4yhFJtRTRZfDoP4HCy2EH3DmmSoiJ3OnxXtZ
Xvo9jVYoiVID/PiQxtRUafZtszDfoLbxse6DrmRtT4zIZPE6d2d24eURn71926Vj4JltLliIgUdT
HuWOTTIsHGNyuvrlZBicsgMpmSvCWeyYD1uQBoZ08MB/m6QDHzYNy+53VU/EIPA4mhtbEHoMsW8h
nV64RNX/1ZFr0E35ZjMAWL3wie3/3O3/0o5BqLN/Gr5TcJfGCDmrSXLgKTh/iJv63nwUTV8WhC7R
75tqcfk49xyBY4PBSb/rS+ZxWHP93v9Su6gK0cXLdDuWV+HBViotwK+MeDBK26pvn0VOeZjBWDQi
4e1//hJQyKy7Sf3PzSbta63B0/yqiPXbkq9C11ER/rFvVOAiyDe5QmCapbn4+6jlVJ5SkV2CzIr9
ZwRJyStWvT6q8RhyKW8xUQP7ANYUIAKI11TFKgPAo6cGmFlGTpKAiVHUpVt9Mmfzwk6brzi7ErRl
onEVTE+KbA7dgsQgqt/o1eEhacj4NnCsjzc1FTpuqzKs0OlI/aJizs9MH2Td0hb+RJMPxIHUUf7R
3BLSSnPYS9T9AKg5gbYR4OaFEXJ1vMyMdiuTUt4kOoC26J2K+wANMbD+6nHWUV5SXqY7zpg0o1i1
7LCGDsPe6SP89HyuLQog5VOKR/lZccwwaJe+OG5uL93F8mZbcjuUaNBCqcVrs1fnKl9rQRI1ZwYK
KAMzdtI705HjtXAq3skQrrkyNOHeGZZAgCFu0ADi7aeKvuFJt3o3pdPFvFD/EhhEgy0QFPvwciy6
62pxYywMyyxMkV9Fw7kGKzNHzwElcxvdUOVN2Tc0D89YyRhTxnq2svMwvf5e817bQGa7wDH1yq6b
tmDtEPKLU1l6Op79viWyURKXeAT6zpp6pqXUgWa+VEtABIkPnsu/QDNtCK121GEHKAh7DRdckEKM
htiokNJcXTzPQZD6N8JRaDojC/OAaT8az0VaWIZd31/IL5CZE3QnZGUJgMl3evGbOxv21WT7KPuq
fjiuAmz4oat1o3ueYtxn71Us1HLT2p9fuN9kLuqQenbDJW4L4rojeeWLeFKEMD9EWHL9O0Bmerx9
UM4fUGM+/SIuLM1Jwh14tuAwk5lNGmv+HbRmJiB82dgvCCFkyFd/yWWwcD/XNGQEAKyFG+kw/mQs
H68gXe7zDviXAci3uXbB0wbPcKTnM004qCRDtUek/9w5xIKGeyE9R7Amf4QpwManyp26lEjmGN4a
5eOQ7LypNYYMUQLBieCXpQah9RMcqZOQR/37NBoQYkU6XID8ybRXuYH1gqtZvrmeZzxdOAbO92zZ
kjWW00IqSFMdjI/o/AlpG8QUTgpkX3BEAHjtquuB3+Ide3OyYlXpgi5ivuN1oKHK7XNwsNeV7SoZ
eyPpM6wsBNr8kGjURqx+fWMRGhsL9+Ixm11oLmu8Pi1cHP3BYhtVXiHXjPxl+RyUu1xJ9b6RJN5F
0J4so6TW6qTkyA9QXRKe6mYzkUwgddbfJolb6QLP80IiZVPkF+t2I9sakGYlk9Wg6H36qW6+raSh
+I8iVa8UOXMFa2503CuXBJTtQyWvM1Tr1GTrB5M7lGP52ThnQlj9ndIzjdmIIIiAPib5dYtpz7qT
JibN1YfQfvO1cQ7TgB5o9R+Xzw2uSCG8g/W0/w1ydR9AT62TqdUKPJC4UQGaTKaMplvi8oqhD/+q
3kjwEDVZjBHQ4dZdgxtD0ih4kt8rpPFb/SY3aGg+iS5pvhMdMWYFS6P/DzSFgddA/0gYqGYzImJo
jtq60MxIVQra0nG1kRKnhGXh1eH0m1rjCCJEzjDCu1aG9KgzONx2wsWiO1cr2DI+hnJjIlC62exT
JndRZotSbKqJHtLf1hgm4dTlh6oY4dyUxQLLqxVDIez73YQGDSSfG9oMbtfSwwDB42kW6laA4LOc
l8g0RidMYrx1u06duMpciO/DqaoOWCe5oSJ2FGwIXuXWz2yySAxtDrbUG1wlMK9ymnF25e6awYLO
d5Oz3ManaKaZkexjYWBDrdwl/xCXwGtI08HB6MhVz9AGvU23xJw9+JHKi6xFgWhJyeaQbU96K8Tf
VVfmwyIcmOSMbABNlDdMILuewcHyyDjEoOnjoEDQAlG1nvVeY8EDi5R2dXvtfOOS7jA/PNAfC8A0
e36D8yTg4yvMZwomRK9EtNN7bf/gM/D1GlnBT86HH8ftJk8CU/xu7m2rc2DZ245Or6NR1KYRFwxx
Axl2v/Lk+5VZ8Z9yQiJSXTq/vv3hugAwqrZAuges/aPvMWfdkZPnXaYdULGu2E3QGHp4+j80yCAx
bCTLqO75IYBABTdhcCl0N7qdSbF0ZOGJYAQ/qBUYy4dTZaErS/ofncqqzXiUDGDcIxD+xFOn6ekP
1Bj7KK1BgY5m2lFUysg2pCSTqQ7liS6T8g7ZzLNZGmrSrpFHewCswPhmcWfQ7dR53afXVI0JttKk
xg9G6CtjRGB98pvl0RslEM4egkzYlrCTCrVZW9bzINJFrWFnxFPlRlLHUaYDVRxOACEvCwajn7Xv
P4NsSFrZBd/QJjzvsw701kZa6rYo2vzFR4zoFngOqdkn2uhWs7tsTjz78oBJx7sF8l2b/pbdpc7P
iUGG2/kU4Xe9paANSNEbYmqJhgieOEgFSFVE3u2P60Xzqur6jyIKKUcln3Fii+5gSKkBN7U8DHqb
e9GsozjFNwtSVJGHQseA1gtJEZaOq5RkMTAzbv77Hm43AQ+ffUxsr93nVf1nl7ajuoKAJM33opde
lbw/YSy++nkN2by7RqVEct5v9EtPndapnbyXiFP00kbRsI46DFKaFA5JvDKtxPT+yctG/n1Dpt2h
rhg+5SEXiCXJjH6BvoaS/GdbTFjobSrJ2hWEMLFwaRWg6qiWtFUa4ZfwCfKnLlL3PdSzbKLnHiWb
CRaA3rrDjtgACpPltcIA193sBqoZsmZQhZM+xMZvQ6aQxFf86+JZEi+ryfIi5kYeQtrAbCBF2n+p
wCuHYgAXg8UVtRRrKAdP3wbj4y9wfrXNA0mRqVPTZHplrTItbV8Y5DDojigsy3yHvrZAj9f8AojS
3GUiHvRE++JJTh6Z+u+C+XHPCmmUDLxDS6yXjz3wy3RAf8qFYub1GoDg2137axSSiCpcu+/K9+4T
YZtn+hnwT54hs5wghNym8ngB9LE7KQLtJD1PHM3xEg/t9EtIT2UKTCbkTKX1o7DUUg7v6dS1P9dj
4nkPZGsnjeVBER2Q4+m/2hgHW0Bw7lRpJcxwMxCSZodjSE6lSDI5ZY8/eUjfZR+UILKCZd0pRClE
QBJE+tgHTI5K/mQCVffdCj61F2SCKKp+1DBxEQOUrVxbJdcVspBM/G2/MPqBKcu8KDFfVL5XfgBo
RFws9+0RvqeBJTnBWGT3/5R/sr4qdOiZ52LzoWcAQCOdo9qTAEXbPZMsaoyiNS4QvWVmaG0KiNAi
N36Hf1gNoQsu05ooQiQBUBbrz5c0WK91CepJMMWQf+GrVourXNBf3kIo4FqSE44bj5BektknQkFJ
JsAvmUZUEybnnlO4Et89eCVTy9SI+I0uK2lqzT9qwCwRKSGck+1nrHQSngvOMK+6r2dtYXVGqTUv
T4BRSQpT9onr+eoRkkme6uDAm3MZYzhI+fjyg3dNqX65ylCW/il1UUtwjk8Z6Y8x9DAxMZ4CxDTO
ME3zJrFI3t2ksc5k0px8Oy6c9rkHgSYmT5hOJEK89SP/aBqxPo5Gr74/7enENb18JeiEs03mqzBb
OY/uliTcNW+yQQxmkniJAgJVUDYZ5T3Muwh6nI6tTFPH4m2JPIYfusKXlmj4NJPzR9kKJMgTGZrI
jCMWUGcpWOm5DrGIKy+OnBHdF4ebgz6//ZwAg1on7aE9dwzn/RmLdqKDZx6i5uIaJUgqXfalj4gK
UJ6lbqZnAc7jQM3z6klVDGpIzr3xasahKpoPgfjXMmpWhiwu9OyN4BJ9eKi/t98DSnDNOX5q0ggj
O3PBEgo3mnT5IQ7v+v00CzKzfSoQoWmvXpV8mQQawKKUg3ntRACBVrtMMn6UV3gETX+74OP8VtNl
90MvYM7D/8aDh8wPOiDBX6XCh4wqbWv3ocym2Z+n2CY6rW78sri/tAu8DZc0jLFzZpCBqa/P8VVN
ULzzg95iFaL6HDmMbM7ccWebkVGI1uip9MfYOiDOBt7GJhGQix6s6y8IreABSYQa4KB1whryxQ5W
w2iXFijDL4/UOrGoNvHFA86f3ycl+1iUDSHiIlc7qvtYdS30ip4KH5aRZRXwVhH18ZQtFGHGCmz8
yWQt+LFk5MajA3O+5vXp3BApIV7qlvnrwbqFf2+iGU0xP3glHfZVBifPYu+aY/6hJHfh1WEK1jJ3
QV05LK+oMTmyE36M/RNIUorthPEj6jLC4Atpoh+fN/miZ4nyyvMCJ8uRqkFJNH4cLhWca1VrOn4A
zBdmS2D6rPfLQ18N/xyeIGXsv5/O5yCSEotDBqnuWkPcBqgHqCDKE2kqXlbHIcJabrjxd/1Jftsi
+KPJixN1XRMTN8FgXE6rpxL/Vu7+msSMdLHnz3oMnyD2ak2jEpK/HbhL0711daggZ8OreVVpaa3m
s27h2SYlzc9B0kA6sSgwuIqU2waa9L3utkD1IkaurFZh4wr+5yJONM19uvIH7dMhd2ScuHVm2jXq
m7hP8aG+rfYteyxral4uZXqf0NKbPcq1cgRAfA5sOb0F0XZlSgAftJ6BWaWiasotPSik/7qjbCKU
P20EBfbvh4LGK6eT4nrA91zcKwTFs+vbmFpiYXPqoVrKRnVZ5W1pSn/uj2c9b0xBzjlm11tVEOTz
IrqEskAyg5y2zjfxw9TIUmYUhMIi/zVtyhZwCnSYKKlUWoTrnDg5ShdTv6bhOVwyVPmGAHfmfoBk
wWNE8vYWoQ5VtbfP75tBfXzSRx7lH1JYeKHb1GCKXgAbyIqlNi1nMn2uVR1AoaKcAypg4s19PZpz
3vgr/iUOYVdEXXWJZNB/kz6KGW2oZC9cyNv2YO0biqxUnPdiPTz/SUFNpuh8YdBJGMOgcfKBNzod
CMwQyTyIwGw5mEFIcxQDY6L9rEWmQ35kWWOQwWzJozv19qany9raM/C9MWDpqlFWrmaRQg6/nxg1
rhTsfT3MbvKE5YKA89SKnEG9AxY7L2rlxTMHPFpVPB+/VXl1p9AM28xG6YK1BvuPgck/P8tTa4Cp
QdoTTVjwQ9YLNmFs2HobQPYhGHJ8V9FmuInJFaLCwdHLBQZg8pcZdKPnVmrJOXveciPobsSxp7KJ
K0Joj/rqAXRF1qnfphL/f16EBAe+xygtqIaWIu6ZZB0X4cPNF0w0mx4aOLG1DfFonQe79pLtTqu6
AiVVPH3F6vLe9Z3ASdoB0Bj5mHjx8ElgbgpYnp+j32b/yxgzn6DXGVhV0JzczSz1cpQCnUmn8jH1
iSQ5+mNChoOLMReaiIac81UCGI2iCnFJTVIiB+M/jz1dM+pXXL7xlGhagzhnVND8tmM29BiBAx8s
22c9ESskNN6N2pdbmgg3P85krLFuIBLe+Qr/rfKNjwhF8KaJVpbDxzrzxhUPw4Rj8FBSB7RjURQJ
z/w3XCQw++/qS6uh1PdsShVFXGMG+BreTavc+Zmdhuvb13GPTpMLFIEIrV3spQw3ALxocV0EW/DI
Hez9jFUMPj3B+LUF97/7b1pmbVrBWEU9PMcTEjq+bMMW81qYRRaLE308NMUeMndVZTjGaL8/pk9X
W8iQLq4FsgD50CG+pzOP2VPtFkE9xcof4fktPzGSsDf8eDooJl/4h5AXNwSo1++jKsY7Yh6RKY1W
fgvgXMq9je6JEBS+tBHEABQIqa7QEoCWKt3hETwDG8xjMe11iGqqJvUA/lymnZDzYQZonoH+6ufO
ar7XpNLsKfCCV1B/g7QLsnWFLm4fOwizNrypxOVtHaD/5avpzCu1faAHU2vNA49Sm3niOpB4Iu+5
VJDYLXQ69Xm6Ao7pKu4ZNkXFXWGmQb5aCf4lbMbzUFW22KmZ3NwcvGv7pcSpYnIvbiuVgWq5khcA
DwpOa5icCsdITs8tq/atd+oqHwPXoKhqkU4v2aVQGdrj6D00eUNapSbx/kysKfoXZ11KLFFOYf+K
hAKxm0USWxuNJ8s9DsRRQDJJ5PExWUp1rh7pQ6UMpHu8Pg3yT8QQ8zqF12uLZn7TRC/U/jsqo5D4
ewv4YpIKhKK87SHE+lur0EN4mfHzTkMEui5ahyKu+yfxP7w+CDwkE8LTyk5zddhdLQNnLYFuYtVb
8bfMJwSdVuXTv3vVFNfDk45+nfKcVgUf8/fIX8+iet48dzrjt/jGTOH2ktwosy16n2ERFnOFAw1+
iqvfmqoUCRiO2mN5+rr8SVEfA9DJuRKO2HgIu25nmIfhSjOVwzSeE1RIVMTVC1+oyWkhQ6JeVIyB
FZbwz4TfT1mbTzzdBmliQRYXl2iM3d+rwzntXe7qQnRSYYWc0UayTuxTY6xzUMC+YTgotjsnnB/5
q1SuRWxFH/pnILepnjWSOp82OA/bXWE/ha0lkZrE73b/0ViuDixsVgeQdW7bVK7CG5yiidtfNGh4
3efc+3EcMFcnmlNcdhJ0jkqCon+vfxwmCMDQLpjzPkYdxKmgy0O+C775VRY+dfqbvTuqS76XJSfv
rqOJsxHZFh36ykELEjYgfqTiwubUp1ibRulSczL10cwhpyHOs609fXbBFcdLFHzy9hQ6USsus7iy
liV+axIYzZ+G4uSST0nTmxAxKTw39qFZIcquVz1MZYXg4aJQkOBEhuspXVaiEit7IOYlnapiaVYz
Wcoa2ZYGY4OEbdJuUmHTH8IzQnRVMKfe6kjFP8CNcuMjxT/bwT04g+8nCOMx6K8pL89bHv4T9mMl
Xtq23eA9j4GpbrqvviU8vVl7Ym78qZaGnGSB6rwUpGLJJuTMUhoQOtCobErxpd5S29ygw7KX4akY
fNbEGCsoJkhfTxM9IaRTZfMA7uuEtaWysesBylAU7AJcpZUZ7kVFZFzJPOfAxDhFlgLZg3/AX9/f
B/348SfnuY+81urmxxj2WtYumWYN2RyApTcN3j1CJ4y+v3fLG6B4P5PWECEnLWMch7v4kwA4p8LU
/mwk00bZSUhq+f+Y6IT6Hlj3NOb1zBUL2Q6LVnskNc1B7jTO5Y3l3c9HDvVdDIoFMoZusLkYxeQH
1CKiPVp4BtO4pA2ULBAOjSoWt0sYLG80TbgvyaYvEd7/jNSwF6s9mzqTtFB0OtfkcUsf2matT55B
BItjcKb4yguP3ojIdtocmxPFTbtG2tAIOqqyNfYPrthou2qz3xRNi9Xe7+NPgVOgpOa6Z5sux8/d
L0egoymIdXOXt//5oWKS6fFPXiJET4wP4T51qckepXlUCIbJymBKX01CchOeW3Zznfbo5jh1Ky4c
XPrzvWZh+fwPPuLSoHN60wOvvkyddISc3UFtv0Wnu6QuW28UVQqI0KsPl2al5AWuIKfwb7D4lJ+h
XysNEhmyIPdM46pqJNzzjb2QcL2WNMg4gwkCHeAQNo2/V+sfiVtVpoM86d+0+QA7WW/QjCQRUaic
RDu7VkCBb1oik81BxTNoye2gtZTR/OxnpQbvfswarQrm+aInIdKYwpZqum93Udl8HcsED6iDdxfR
+/KdjrdZAU5P/UcSZF9nCjSLiAwb7Ym2HZmVBD36USMYhXYnD3zVp2Wr6QZ+lzk8/WFbV96NOs3J
McgJmqj4zzbFbElKqeIdMkmkEnvS8xpThpY3eV0Qn8DW7anjlFdCGQjJja4G3GF/mjZv88RWvzrb
W54RBPZYaMUD3CajE8FDVP74/sVnC8Ng2ACo4PKDBPj38DC4e3SYTSPE6ydLzFH4doEOlSCBc4+Y
ch0vuJ1ewxnAIUrqhcpdk8vVIqH81OI6wULJ0VqNpuSWUj9NOyVP1Y6xd+zFHtWENMcLAPYQ7ROl
Ntr/qQc/LKLLZnHXSo13Z3844+8cgVI+DCs8N8vKpCOPu+iSUxluhv7EGCk3kW35Ay8oK69oNj6L
off2oWsxtquwWHgEdLi7i6DuMzYHqfZZOJ7lynGGcWN3uDR2wdBiandSypdi7uef5U2jfvtDQx62
G30iRYIV/Pzwseol9xZKeQrtIV/Ev2GYO0AD/RxcH0dqyB2nkE1t6GhUMuQRfe4RL/7YE8sFLD+h
S/RUexz2wZp+SWCDde++PZ0EdSQUwwV0xdyzkEDoQhQQQ5cr6iM8JNElpsmGqxd9ud5Lkmvg2HhO
oYRQhX2m/8nWitQYLy6oooA/iEq9KZ+LvhS4AO/Zgy6M3OI36IG1qNEgwvze3H9D3bN5cc/lpic1
fyPIT3y/nfNmo0muIiSLCzb4EfuhcgbH1oYUdtZHItos519iSR9FiCi6uhRgaTNjrQ4/ap3ZtVcc
s80u3JDFPwjErXjBQBA6yiKMLCxLszpB6taLOnc0M1HhKr/04iyqphsnCGLw1FrHqpY5LuVk1map
EK5+HLBxR0IRPP47FySqInwJSWhds2TlSSRg1MqlRYrs2epa9ASeACdgN9+Fefa/IZDulD0lMfFZ
aWo6GkXNLRnnyjfjtxPBA3imqZ6BUeZvKM2k/1B6yIjdd6ZHUIJsMmuWovkVl13d3sm/rh4OWT9v
NzxHvRLX0zJTJfHQ8RSyVYNw5rUmmW3eOewYNMJ+6i+bep55atZ/193VF3RsCVGLfVapd+l/sF60
pbnBk21SijrCS/l7jmoCXFOKhgiS+Rb1dP/n5+1dYoZ4WGgS4n30NSqpWvIhm2KGJVWC3MiqMo69
i9fL4/0BSThA4GVj39zLfPW+WcnhWmFJGGo8ZQBsRFpqVWykjsy0Mu/SIN4LDgsGhLPdYjV5q5oy
0G3imWmsobhoTJnf3CiFQVn1zRsx6dDdQMnkzaE7m2+DrWAFjI+yEd/NX3vKPwSevNzI+fzeh5Wt
sD05XIaKcVPqSZnBvFvJSHZGYsQ8YlfjK4/mQEZo78Qoy42NkCRxD1RlAWHfhHN4HW6t/h/yUe1V
govXDn2SgvIErbzDi9EQv4+Nf1EhpWcj/DwsDVIfJg1dJWmoLRs614XwEmzMTlQBYBwwsAYXz79A
SL1fScycmAroRwv3y05tVbJ0ptX4hbjplZvU2OaDvYIQq+zaACspwzwkvbn1KQNU7yIy1jL/094V
Qn6Ls3xRUrTw7XXObniyykKDM7PinUmCgXo1SUkBPmTFrlXH7xWlxJ0PowcddBc+ev3Kiu8GLoiB
U1MfopHX3917otRwtcOprHEKmLBwQHZ3vAzKGwIhD+Nkn0bwoUx9WKCvIVJaUkixclHIDPIeUh6d
cvaM0A43+Pvum6UhvK4j95uruwHpl8M+A+KMfsYGZFcYRj1nuk7SK2SBJ8u1ADqk62zagbpN2wB0
BI51Iql84LR/kx/lLk2fyjUmqvWgAHCLkSxtZCZ0osmi/37PMJXFI3VgiI/j+bnKT5g0wh6vTsNz
vEB2/+KLrOvmKVtU3unRxqJPQIWXUbWz7ZyQEZ63IMQd/a+LevvyY6jnfBU/IDiw4YnZ4LlU+I+M
8N3DGfCtVgDZ4G+kHuch8c96V8tVS1fSyEgGEr94sl4SanOMNy5LoWj5wrvZr8WauedtnPbv/pQ8
yHKSTv3b1Soj1bi9zK1Cl3jARAsXcuFWJpT59WbvdENCIhQiZXYCUxQjRMsgR12UWi8JdHfn5xx5
nV9xb78Q15D8dkScNl7CP7e65oTBa8oF9kiJbg4pTCVLeLAI8Dbkir499Xn96PSuZh1RQ0fVMkai
xgcxl5txQ+T72vciEdHuewjKvJJTCsF7skSTgkqneKixsMUgu5e5uZU7Ha20ATx+t8KeKYgoBbdd
n4xA3d9Ul8rlFv6uVJgKkBciWwpmq6PbwyDHGKlpXyaTSe3NVHG6W7BYCuLnT7l7EnYr/J5WdTrc
SyL2L9/5GF8nc6tmiMiN9nptdor3reGFQUSWa2MDqAketBjiivd3+LqiTAikrVFYU5qtz8jW9jz8
ZTkV84QqmAQxneguZwBDK0GvfsSZaUJqhnSo0cpu1ttFLi71Qe8w4pnmVkVUkXp7pWa3kMw7FPcO
X9aFflVQD1ZGAHgBnM1jS0s9Q/F84P/cp+Kapz53jZnM1Q5nhv6yhYse++Zk8Ar8lK6atdrUMQ23
PDyHwAT/RBZJ+nDuciCqVEl98nZz/hznEV7+jiDeqBYbVL2K9Wi+ii8uXpdo1FH+SJrhsQ28Pjd6
GAryUogx/Um/D2YpwtY72mfvfCmUxjzHqz1Uofa8LpsO9U2o6WjsuVXNG+eHPGiG3ZDpHqlUdL8b
6bKLvZt9/iakxqMk2FOJJUALmwF1UkrRZOjWOLngamSKxa++FnlMKFS4wN80jG6BExrVx4GRgsKX
GoIZZDLq7CSE4wfF+GUlxFotYUzHzQfOvG5KWi+cj3lcYie8YPO9sokyGubfYDwMl8Slb3/cu+sE
fkPNGwiVqwxy7RY8wGEou9Zwz/uiiZjNVElVdqzusAXw7k3wrOYQByAyg4u6PPtpC0lxfp0u0aS6
tHRfL18F/RLy0DJFiezsF+CxsH+pOEUxtpXY60GC3KzKyjeKnBbCESgf4uDP4FlrkMI6y1rMKuGo
HLry1WTPMrWPlHJYoTamaaSa8ExaI+AByeVFxxuqp7rUJrN/Mai56WX1xCmDlb2i6eTydHkPRpdy
5wL7Hfu16sudL5GkvYNU3HzCN/g4mIhTJp0Ebv7UzhV6iHeO3iTZ5b4ikDd20JGmvX7iw2dB90FH
nfUV+5Sd0tlw1Av5n07nUCZivHGP5HM4q9YOZ+YzIwSRabtDykKBuplfKFF3pSWXoioyFNpMiUBe
pgOw0XME5CNYmXLDYQapP7vyAsImn8s0H6Y0tGjaPutaaAb24I+OkwAvRvEVv82/vb5j8WX/Msa1
G5ovM4r7YObSdoYdAQm+2Ab+FvVA/4vNWwMZtByIaTRA7/kqUGIKdVM40uiHI/VheNiDfT0D+DhQ
2HgXBH9Spb9saKA/TeXwwXFOjC+xpDhgza67Pfr4yixcKpwNzWvPa5s6QYCnEbu+GdJFLnj2BHLb
I5xkzO4DJrNqUxJqG6akmouFfN9CvWkXc4tjtGtNkUGkB6hG5dkTuoB9xBkXmNRpbdY8f7dgkzBZ
7SOkexIeKCjSlqJJe1yUUnFSUH+cENtdmYvn+HaAURFjOOXBKUd+XDwCWKzg4xCtkvrhinZOnPdL
fLo9LcHW+nxrhnsSt0Z+o3WZ7EPdRmppk69b9FRvYyRLctkjz3yGCHVtgoXlYBoBjC3V5ecb1hhx
Nbd17SNmQ2rORHxPh8e0oz/ExLHz/I5BySOweaWBhmNm7WBsg2U0H5C9zfXHt3AXKUpv4JyyA/yK
SA+qEmYEgOcv7HVDu/c1AYyw3KAnZijWimyrXmcjgkU+qWdQ6+nV9W5GhG2AdABJJdEbO3UsTkfF
v1LbWjoFVdJQPxD6enKWQams5n5L4wF+9woBgRH/Dn1EKYTvEL634xO6ErjJoxCczKUjBEz9GD0q
A7vauutM+LUhzVrrQN7krdSnrNxoCg9zSEzAap5HZdh035jimtGlD2mofumk+lF+OdX8jRiLR2kP
apiu+8JxDpJ54z3xswyouQFGI0k7vdkj7CmSYbVfMixpoLk+VmDiQJfO7zj1Bd6UM+cqr7PCisUO
yKuf6LmwhTHRMF+acrc0fDrl99mECgZZ75o6CDLQIrWrl+ym6luOLC6cCBNeRbLsLgg0Cq/k/lCa
GfYTS8pIaFUMKf1myhyLikP34BvNCkiTZJ0a7lx/5B8NTInjOH9NtgcH0y2C2q8NuHf64TgJQ4Oa
3ri4XLAIJcp03aQPizEsM2oFNt/CzFBVJ2NHbNijXqAhzVBuKrs5iVUUzsnWGdORb7g3/OZDY9nr
gizATgYJFOcRdc0LSte2WfrefltxMhP5K//B4QRfS/ERGICllgESWZzh9OrNCDeb8g+PT3yvco86
N/Fd1N5FoZOXlLUzmfeOmBPL4VHUqVWoVMsJwq6CmJH7KHi5QghdE0Rqkta5bmMWx9zPY8xo9F2D
I8P6XR4e467wHRH7rY5XdfTrjw/ipcqpXipr1s2UpZvPSKNQdgA0HMZHzrOlxxP3ln7n8QhD+98j
RXnzM3O3Q+XBSvSoBmH7mWPQ4+rYIasTLndVnoqnaVWOKWeoeeK1Q7raiX9elOlNDetg+GjboyhY
OAx2WtWx56K8ywTWN91MYcd9mwJJxGJ3EVOe5IOBHh7B56AXnCFHuIal9et3VTQn2tma8QMuTl56
iyOcuBEQTeQuptSTBZSXSQHzaxE8ItecDi7i5bwZCq/Hnlzmx1f3uG1gOFxqVLbthJVxpoGeyl76
MaId2M9PYSfDCs+n6oWzDYUAmTam8LhS82Aa0Nep01RA1COzKsrZc6BfMJjVb4N5Lo2qnd0nBo06
Oc5nwpL+5nZ3y2YBRLkVHqzGtkOSKQ/UwoSMRrJSLBLqqmvvZPsP7NelyCLMwymNOyQ5INKWN8hp
xTmZrBXJ0I5YGVuZpEz6lX4pmS0WKS1iPL3812G1d4RCr3HeS8yjMiVawKrebUEwaxJkKkglElRk
G9WIOajTNkdQwcoype6e5DaiihxsNoUJqF/nJ10atHKk+fU9t0KJBxhCoBIcdwciI0o9vJ9CiNDD
mDkMDsjdEAW+QLT1UcwlJy01ZbmHjiio20axcnLbD6R74vfuXestr5fpJMML530/d/Xo6JBZNAc5
woA0nR2JB/l99g8+I30MhmqHmrw0JCbRxajl7fmLwQ9dP0YMFzLEw58j3oDJi7ChpKMHiGFJhz64
lUHpG9+2QQ/L6m7hMoVbQujpBFSSnvOJ+9sniOhJthgoqboez6EqyHajcXFohozqgcsB/qkLvGUu
B3CFZwzyJndyhh5uC9IW3BGkfVehnjcdrpS25da1CJv4UTx+mm91gweWy23myHqxSybzTwiVVSv6
xSJ+MjGCoN8ib0g1z8aHqjZtUniMQTnpcRXEoN5eZVruFiM1hjHPgm5QGmdm/D/d2ikKw8pTbB50
dIocOMJKvrtEnMNKywcJCwqW61sun6kpSEjx0/qKcwSGSq9vNeCnZXjwDvtpo8Lt8glTsWQiOLYm
1PB4lWAPfIOr+zft6PHzIVzd6LIEUe4RxZB2BeXoknE9Fam8kPTO9HOhsxbn28QpJ0MrocfFia1A
JOeGoXY99h6KGvjSXW1jybE6wQFmYs5RqQppNZ+WMPCvHlFWEcLSEv3ZWunvrOSR7KDyvKYC1vqe
auxASl92dPCDYN8bnNi8KIMAnq4inOIC/JdEoyblcKuHBTT7LJz4q8yDL2Wflnnmbe7Ui5Ky4Pp6
JJFdVxXhtWPaJ16zAV/FfQ9iLKebOrKE/Vdbj8czFzTB6LDSDBwk6deDwBRWEn2QQQJI3GSHMnAn
h/VQH/NkuJhMBdO6TTmEavydhpUVHISehIG5SWSdTEe1K7LmV0LFDuM8ZqnpzP2wXZb0C7o7nk+T
AyQbymyy9LEdhyE4LwVxImEpiFmKsFivddwiVhYJ8P2LzsuYc4NPPgnBTwKGmdO/i4tBjYHIJwAt
7zQKx871zN6Hnc9OijJaMbnOhva2BfaEwQfYrxi0m+v0b9ukM8rjpQqOBm081tR4mKMbgwMceuyz
eL9e0iR3h2l6oxgwabt3DKdmJGqS1HOmkJZXg04NfnT6dCMrRn4c0d42iIaj5EA+yVfhrNrKooRF
PgGXvQosrkqE3bj0vH1p1PGDPpU2j2Ld8OqItdOgRa7AfiTHDwljsV/QIIT0Tza9Y+VLhvicK0GD
vasNGVFh6GKZ98KZBRHc3s0bUah3qwM0abseHDD1id8x0by7hW33KnI3C0I6fozeGW8Sgo9ZrQir
zz8EuD8nk87EHvywt5xEmW6W35649cbH3YVyaCjMivXmUKLshKs/Mqgi5WZd5lggzWH/9p5b7/+O
3bhWtPte2RknXN2ieXr34Iv0kGEBOYvvD4KKh7tfx++u3I8MD6p9jIRXRCnWCEJ0vYl73/Ry8G8v
Kcc56bImFFVjYWp2NoObeaRUIBZDVgpmjxk2kK+a4s3w+3PHhz3b6YpGgjng6z7lSkQXxAdaCHvn
Ap5Z9ZEMyGBfRP55Bh5bEeYJaWf2Kw9sOkPBGAYcFDjDH6+1JvWYf7e/vP8ir6++k7iauJ8jMaub
6kFr/OhYCWRxzb23tJ/5q88An99P1dIw8WxTMFlMJCv6jw/p+lmpWk/MWq50xzjEn55Mqxuwfksf
EkdO0IdW4kjKN4ljen8zu7t6SoB8Kh87AldL/5Cjl88XJgCLX/Iq87m0JFzPwmypON8Oz8Ff5Sui
j2ywgWrOSNAEK4/pBDQvKRaT/kHEfK0tDA5GthwYTil03mwYgfKYP+Em8JgPsz9hATsNxSeGLqjJ
ydYNflETNd4cEbhLqNjd2z4Qi8V1upV+sSJTU4V/TYi9RYHpUNcwiwhGlHdfvuOxpdgPF8t7rgtN
yjEHJqN0YKbvubJGtTQm/upKchYVgQ9rYAnTiKhhnL5OHHFvwPjwym0y2Q2JX6vebVOsdV70AWsa
wZR/did85iqWVz8eO0X608288F1lgeGo82GtLvyIWpXt18xbjlfRBVfACAXwFy3nOIU90XFSVTfd
AE9CzuKsmVrkUtV2uJTqHEcbjnvYKDWePlLjBMB3IeVeKcBu1Rz+Por13LV0AxwJMu+cgoIqbPrx
bQ3FRvTPvCAHtahAEbpZPQnv3kpjDCUpA3dEOKLRtl5JbL+facNTiKpe8GrN8D+pR9GZo6GCZC6Q
AZzBOT5vYkTHiDIlNSl6AxvnxNy99Sv0aiBjg/qj0hKPPAiyy52/wLZI+0XF9mojSHIsgBiVwsqJ
E/wG66O3X8KcX64irS3Fwd2ekoihxBcA/ubsH9wB0qf6w6JIOA9su7gNK8uTO6fF3nzb0+hP0R7C
q3161j2upLurPkQ/xOZpZCdZ1ZOWu6+S8XVwEWA1mdqM1EWK+M49RSB5PRIYlGISlPz3wbn4TL/L
050k8E3h8vSm1jsCYk/ldLXAkZAnMV+J3iy0295nRqLVkRWYwymz4yTv8vitXnslVeuhzk89paoF
PYQF95tkkiumJ3S0IfbFi9awU+eIWMN6WyFmLeSg+yF1GMMcQDB0H7tJ8ykyuSPWirPearipof8o
5Cn+Btsn+nJwUE+z0iLEaIx4Vfi1SplCbZooqrurvf+MeSv95fZSLBwl0685RPJgTs1Y7Jk5PY0g
IIEXVErs3r1dz41OxyKDPGwyqSl5229Idt12GoT0oRi0bxH1bXCTXkV+oSQ25iXXXTx75X71z1Z0
5Tjg7qRlfX/MsyBQOuHCq14vpDzsf+3ySGf+yww1JdsnE3bUSgYkEXhhMnyqPNM4BVDUCwCPE/Fr
KvOyxLiJi8pni+r4SktfpUIAS3SKDlSx+YTGjEJoJI80ACReFuNKkcd7F8e9pWbhy/XOzEUEzz1Z
ubjhBUWlUMsyTXFw2Nd8IcSpNP1/vVY6jr+Wk+QC8WXihfTbBUMO1Mr8EDyW8FtBQhmCjFl32EZa
hSmGydV8tCxlEKJ8xV8YK86gm/M1B/77I8+MrCEdXXoeStpvw0u+VIyN19QDHRNWuUcBvRZUNzOH
FP8T5JSsPu6VH2ayzkTqYRuJuwUoaqSlfbK1BW6y8U0hGn2MZf4sdG31MLD/paaXNZbbn2vmPnli
BfJc2j8di8IcUpBHpV4fpI3g2KQeVSCEt4lvF7GoWziR25FHkaTHOjfwWPv0GdW2f6+zEAlk2+MQ
OGuTFAGi9XK1FsKUeF3BfCSR92jg7i1cO1GdUTakUYAUFSgp5lQTBm+hXSb44BOYZHWH06yXN9TP
2UCUZwvW+tq6z1znjKMorB+StNRS4UC+coLhYp/phg47Z27n6cYBaeeEnKjrsSZExglxpbp2MXJl
OJVxa1sGs+KEYmrtpGAwjQWop9S9YdnyE7xiljUACpoFIkXTfxS9zRr08fpEZsa8XoIbTeyWf0dz
L9V02mKokLAq5piNmM9Ep7vYpkH3H623GjwQC2rJadaZlfuEOu2/8fQ6QlmbpBNySK5NzI/6rcJZ
dayy97mXK8ut7UWW/Mr17SFcTYJcJUAYLG43kanfCRcGXYdjbazPV4qoFDuHZGFj1Lc1SXR85Tf1
TFYgFZ4VdAzpr8cPOuCpr4/D9GvsQ6y2/QLhZyRqGaR73aX8FACBisnape22N7AM5mrksDIJRx6r
Ao2Cqm5qCIhNxCkNSVdpLXoThu7e+vUDPiR1V9k5potYaSprMko1bYSIV2eZu5nWP0UuKxxEiKLn
8/064/lG03cjNblBl9k4SjO5cKcFPhi+gPnFz17p225GY98bHnbct/O74UlT9u1Utl3i8dSyOb7+
ZI8uSHh9Iqsd2gXts9UjUBA5Sokbe8ARdVznTuksL1N+yrV8E0Akp3joIoGalIQ8uZoS+8zSX1V1
eC08NthEYah2OadggtQ/1cgOaPnI4ONNJMcmTohaeDotFSe8WcXMpJOBCmPMQt/7o9lisoK4h5+s
lB17sO43QqrI90oxLyMzi6Uv9wW3Jgdd8Wsdu3jujTj63XgFwxp8Ha6SG4PuWo++qsGns6Y1tsEh
9lsnkAPe9FGp5PNR+eOEYyeGzdIPxxgSX44RWCkrrkezRw2R/HfreleOkB6DzDCFVl5VFFY8ETni
ld9ZRAU4I1qLj5TD2y2Tf8IFA7wQFzUR1xauAq9HgM3ZDjnKUV5nOecrFPdVHN98xWCOTb+SZOpW
GV7dbVytu4SYWzq38RkcS9fcpM1YD19UIQCkMJa/yXh3rDGSBkAWDIlMVPQTyMmIdvLASVCiv0SF
BnJMwLFhfGCWpIjgbuKm0bb54P1fdSWQrFSEfPhzhqJjRWMZ7daXL+DgRO6zElJ+Uo8UbdSFzrkM
ImmbgHcvii087dBCRK1MSF9M13EU1ty0VGogUEo1zjpoErTbnauiWSLKyvBLlV/nggiUZJt/ZD9M
4KcM4rmgatXxblON8W7Df7KZGcp9dgtgbz7Ze81sFgng2z5vAJsPcDWndgTQJihwxQy5t3ys7ZTd
ystbJkJrq33S3kPzs2xqAKVixXGZDJV+T23pOtUyuoNksrzZnkWL42T/eO+NeQvkntlhjmnE0c8J
grJyi8zLIwsL8Eing0/4f8TjUtg4QDlhehW00OZn7EbyVIt091tc3ILU15hhlIucT1YdMxwj8DuQ
AJkKg5qrCoUIj6RGsWicJzsm83sSEkf6r1p4TN9ySaPaVKsdgBh3og6Y/1I3EGQAEH8pjpTWtk5l
d1apnaF50tB3oA8CXe+akkPnNIOH1cmQFeMr2qAFFz6uAWgsX8sB0wmjqV6ontXmv4WBp7sxl4tf
LjCWVVCdIMl1JZzgEy6F08Ri6FwuMETX0QF/vHZhXBOfGH1hAuv+kztJA5bX+c6KrpFkhDZLsiQy
EbhJ9enm+e0aTbxXwzJQ7D0ZcUaf6phIbcZlIkW8LZfqK2jQH/sY000HDSPIQrOrfeBZE7H8msaN
HBaMAA0PdEIvVp1jGyxRN+A1igdOLBzAdM79p+XzH3DKfsf5OYFg6KWyhHZRoZ/dFI05j2mSvWVB
I9+0MFXs6f9IVwLDqQmyq0gNxXmVJsYl5+ad3DcvDoMPpO0wML1jUIDmlEjBNF+ZmJYJ/8C6rAuO
pW3TMJSaHEBzIR1NYKVrCONOYBEb7nvNLx0BBFZGADcFdoI9/g172b2JZuegDqYAXlJps3xiwc0B
fozQw6UPnIU8SxJgGUgpZ85MiDLRhfHYUH//hj+5rVVwK6/Bej9ANcs0bB1uEevNmnMZ+iEpl4fF
zVb2RXdpHbYmLK1Wap2VhKYlJj11le0TnrO0SVuGJWkCydro89Lh+6HOpxRL6S5afGY1CM4qHkpw
7I84MbV41QVRpFdDayzmJeOKUZATovkoGpPk0UoJm1hqkmfmXb/6YDMayA9dGPXwCPVktrm6DfFE
7k2/glRGFlSJCimVFD3qDivnQoVH1Y2roUCAoCrVpBZtSJlUVL468vxjl1U8HDDE0w/oj5zytu4I
2MB7yb+n4Cg8Z7XnoDVKO/WcWFE/KN6xp76zt3ovajt15VuojX8ZhNBltaIvdABDOiZ2TgZLkAgT
qiX5BI/9+AaGmFaEii8FMHm5FCP86LbsKhqxZWloU/mTUQYURwREcWIPg8+8q7SCOBykVwM6W2vd
Q0iPYIES1hr5pPtwiL8LPyCFykODt5LG2bo4NqyLp/OAcHzggd9BnswahhDxeWN74GLvPkNZKQs0
IytBxMcsEsUN4n9AYhOHxrxKEiJqkEoAHabOp2bIxuzRGHYjr5NVqErIaTca1a/UI1cz/F6xGEZY
lx+Uis7Tf83EZqF+MM8dcKSLIt3ZRWXgTQptfwFpUhDW5xEI9unnVwRDf4Rd9kO5sHk+nIImeRSo
ma1k0mOr8zmqYbVl5ic6r6euNZytujKbIwWJSO/2KcQXqHtbFDOJO09PhKKN7e1R4kfUAjlbte+6
h9Ji7pz8O94APBoPFXFFvU/RGlnFT86x7/sMJd5LIi8nRd+y+//9KmdLEsigFUGvt5jSl9vmAwOt
kkjmAJMOOcL+QKJQpbvvkQvP4Ozr7pwhw1bsfrOby02SoPoLAdS69/hDRHrZKozsz5uSNr5C4YJD
VA2pF2XeGn2C1z89fNx5JXaO3rJaNggOK7hr/g2Vg4g3FicQldIFcyOyof/DtMDJMjIZmNg0R1Og
8FeL0jpRZcxg93l5atq1oLTjYKTQob5s3q3um5391UQMeyVlNYHsQaJ4P6/KBo9B9LvbleAELRzB
PKby04iVmJRYzRYAUMnRZ10WmvCxG9SH3B7egHC9n2TRTlQMgxL+JRJ7kNy+b9aHjE3DOrjB7AK9
yoG+bcLRWB7E29FL+377cA2m5YLorUreWAjJe7B3NcuNpsTidjTUpbTREmWNLpbZtmOIJjPhmIFj
3vaQInWruc6+CYFFGPul2z3J3v2mKGYSBOxbf0+z9CTrRpU1yUkkF305yftXsjj4gD5GlcospGey
APnQZdIoSEGXne1UCsjB6aGyZHDjs+oE/prozfvQgZFOZmIIosvYerWKAVDhpZWgdCRkHBoiV1t4
nJPhV+FE5asjvCMsAVrqWPgkDZ1HCUiLBgrd/w8pgUBmqW3q6cPBAIKWBJcZ2xTD/Fz5okYqV0P2
bJSKJ9NPxPbjpLJ43LhogBC7IApml0v6uqlRuGmoGBuA8A8EC5nX7K0yElaqImA7rvDm75xVl9mt
1f0h59cIRsw0SOxdlIxhR8DW+pQhrwLTjNijiho7ltw232nykuaOYMoSKSdYFVJ8ItiDkmfzC0HW
u1OdPsDk5QL/JjSsRZrVmw7uNBjjdHf0TIJNrZRIM+I8i4LWB4rkdDGUPlnvh+BXUnSXHj3JkRj3
yt+3brH9h3ZpEtFpRLdDYDpm03pVlHKAiFXggL0fskTFQas+GQuuIpqFVqlvkdwoW9AXGRidePn+
llo0q+oM8AnQcUwWLA2WPREg7VUq6PSNI6Af9zJZbx4/OI2W/O/Q6QYZPodyrEvF3xqO6WhuXgIq
6/LBVNB0ns6/oJSxICUPSOYylM4Rx4CE0hK6EZzLVKV43rrEcyaAMM41P8L4AnxTSTmDUJK02nJt
o1dOj7Gy0Xp2lvv3JMq2MjLYeOE2rjf+KetgQUjilKL5cfz3zJdPgd4f1eWe+GDhy4aNviKiZzlN
XsQdrmPoddneCj2AwpB37a6JnNQJmwvVNpdGlmvuBOAkIz9HmAmTnES70vgIy1FfLvcKxBhodRob
wzmie8k+WD5rclRClbOtNkkXlMLwxvrEDiSLXRqxo8+k6yo+Xlx2r/lNbkmy96lGJbmM/mG1AQxQ
ckfD86UIA4a8GydPmQQuqJHE+KRYG8sbb3UhcYiNxxXdo0LDLWXOYKB0YQB4tOMn642c4kWQVPi9
oAp8dibpM3Y/odMxCD4O9OBFErrziH2mPZctpLusdVJItw4dOMlVJARnon81VFZlNij/i8/dRNIm
B3llr63g55HmUZ+m0EcNCvMVgAE4i9B4+7i59Yym4bEJtPkwZu/0n7I28HToGRXMP/15zw/kKJNN
+iExVtu/0cQlQeu0Q+vI3ONnFEuug7U8VI+EGilX7jUrPZDIydhkH2BGDK5DcdMYDdP7Ltc4sBdm
gdrmgm/rkEPgA/SeXRRQfluaLIlByAl46wca7cK1RKoA7jQeTlsN2HLaWeDLBbZlrVNkF6FQlsnk
uq2x0A5XJPFoMMaJ2qaeIIvJq5oDYN0+Wpx1jy+rqteONK/gEK4iGJIwiLIOjz2Y91kOgfpyDIBk
sYKRHPTvJuiHMg4KU9eYKQKKZHzdKMx4tKiX1sReDV9W5kJtuE9bZqxQj60JK4Op/8R3ybFPlTfr
dmFMPRpKiG3UoIgpVb+vyg2WaNZAdkGlGqc7gFRNttpBQZT23TcYBL2m3oo9oHAMSxh6vaEtfnhd
QcJ1TbLrzxR+TOBS6Wky9MAZG47Bs2xq8AiupazvuJZ1uHMJuavrEogTDCPfCo5CiEUFPzdJlbn2
QgCWf25wQVvKTBiPMsS5wmmC/uEjgTgj3gxvynOpQTQwO1mhc6nfu0u5/WE6bJMr596j7Ujw+3jE
TjrrwZh9w/9vqXjgpyqpqlYyRKSnY29g5S5bcP3gneL4aqBZ1FVccuBXrdwtWDpQ6nLBa8n7+K6j
k0xwXtGbJd3Fqs/qQ6uOhOLE7d/vZn2Rko8P7jPywkEcDdVJftDfTq4bQypOQ2jyIRTUseY6TnFC
f+5xX/i++1EZLPvCDBHOahImfZHKJ2Eu/QGgAXfnMs+ArHCy2ibhhqrTLoazGv1GO999j+esRl2C
areCRw2QMtotabsGuEN3qI7NEYoPBQcFb8L1yz2kCqFScm0rZrap8Hgff03VCn8BjdpiOFh54h2W
KSCdQIZ6hlX/OypGmhfFQoWB14gZp1sRRqXoQf+b7k2EmEqDd3KNd+EJDUeUQgNTGY9+BdahzKRY
JCEnISKQ46/dQ58i9QfdhCoxfmG19jNxNQAdHVmPFZ1ffZusXnjdF4VsGW9X4mdmJkMsqIuPFODB
js/S9KpWH0M6vLYMwXOJ1d6nzFYIN/fIWkNnLRZPFUPhhv3H4I3LXNVxgQMwYQKF2c4/3aosMvHJ
fU+hBQMDjj//tJ3zbzhEKZovh1hXsj4vnZWsN3a8EdO+nDTgszkwyGVRtHD3Cy+izkSh9Wquf/mG
jTlsJ0ywPf94yapFXhqp5vQZnoUtSzaceGVZWgBUZW9n3+wgv1yjw4oYcSPDoPDhdNwtrXAMhEWB
8WUglcyuMYV7UpYIMAduqIkleVevkIBGcQu9+72mSTtx/DV07gAQIApIK6AvWf1cwRURmr29jW1S
5FPCLoL3ygkA6xpyaG7UDQmyrmaop9aHl+fQPkqokJU38Yd+ohRpfTDE48mVJ5TKFwKqh3GemaLt
5g1xVXi1B1wnJAGErcN1zD4LC7/XmDbBANONjwujW4kwo+3NLoCmEXGfdWCCB93KXulz+1yXpCOV
0p5VMn6Gb+k4AIykqmONLcl+4hkQUrEY9QLrCb6zV1Eqg4DAZKyASKRa1Bs2CY+eX4Aen9pnERDj
3RiPvIX+mUavP7hnA/B2P5ddo4+wkhxTa4iXElLiPnbQRJPcZoubB1An4N8wMIf3NjdH/FFfdY4F
vXcgwEAk+gAPtWvP7QfnYmZv1YoHVaG8lPnerjXEgsRhjxZufkzfMazSJE++QiASBmUT9leNsOK7
P2aM7K/7w6QHc+Vg/G7P+Pq6geM9kF/kU05LMDr9uNFnu37aBs43PniHUZP5+rBdcyfoXk+cQocc
JhoD89oQiQHSJlQMyzaXP9QQckgSs5FB3NVTmBs1HvTOUKyIdnvLPdUsrUOSF71PIS1bY+Y9Whj3
/RwCq35nxiOtqoh52lZ+2jzgmAs8RkLS3KOj7YXewCHpYNeQ01nkaHNz9UjA2NhUltbFb19T9STy
csIN99tRbiOhtPkJdXMClvnwH6Eyks1MFh7kSv5403zAo0oxQrpgobyMdZL2jNDco8fygvqVLt7a
tAPEpqsME2ainmDBzZ/TC49S58Br+QA7JP1t45m3g7sWYsft/WMeFjbwujDdWy6U5FxWxOPc3+je
/I4OfOWm+7tbAOqDA6+/kz4a4m3x81+KtHwSIibbFcL2K9Uuh5ERUeb4+jll8k/7jNsHmNeOrosG
Nq+VauEQI/KTnvXoE3WUg+RTtFgMNCN8QeyZJRquTvhWH4+RktR80gp+gmt4DSe8v3LCqhGYNCL8
/ChRUTvnM7sS3r1ro0M8NJpspb/BOJZWLWjKyrU+B7+phD5tQx5W7drxRq5hNKq9Snn0vMIkF9UQ
ixLw1ra3X+l705zSDq3jCHC8j0paAgqWAh/tj7IiXMaMpZJ3Zfm01HqvIPyITyCRrX6QK01ATFU6
nJy+hjiKFrVZQXCgUfyYf4ldwz8YR8NYMJdB+vrOTqmpBWFQSA/Apb3XkmDfr6tpil6xNoyc5QK6
pa+UWn81U9kLSlI+C/4cbzK+t9oxjePuLAYKuZZk+gbMPY1AT1KuRdBy1B67sS9+khTLKdrqYyF4
u45SPEUdotq8vfh5f/APN7DUXpKSrQFWS6cIcamUslnzCWyPZvnWjOb5X8eyyoMCnj1DbfPTrY+p
34nLzCNNefS3mVd9pIFAljzbgXDBqYskNShxQITmn7w9z9TRK/y7tBdGAEo0iZjoJoiw1ISjE7CM
1h7OyJ6iLVvw6fhtFu64cdvK28kGDZTZh/qWYdoaI9bQaYVRpc2eCQ6fyY+99/bpBLtfc2KwyGoT
qV0HZAgY6Wfwe0Jg3N2CnupFfrn/B+bzaIGJK1jnR8rBa08wQIrE+23SU6mVXyQyla9r2wGRpuV9
aCcazWPjKPIkmY9qMoFDalXTr+mgnAAfrMY7lfBL8yfwHsYybjRWV+y3BBiOQtMCGSINGbfdNS8X
M6iiVICV8niRo1DlZ2VEBmB0hQ1ZjFc9JIwb6k7As0F0HfmPx3CUgm/BnmYN1U9YJG9gPQLeurxK
Dtu2R8cpTEKZmCd5B70nV4hi+oPyPkxza9hYw7pZCrWU4DogXWYVbN/m887hXJNVcEOBAfOBB1hj
BDc/CU7JYSkXBSwb2FwqcO/DyvLf2ZktrPonBDF1jpi60eqE5jOmtiyIYSFaMkEH95qVWk9nCDeP
jnYdO9WrWnE3gwat3tKIPr2Efjilq+/UWhRuFzYHL39gbMBKIEwGhu8HB5K2Bkb8kCyxXDj0pnpj
NU/dvq69b1d5pn5H6FQzowhKofoR+fqpPQsqOHByWV1DWuF3o+cNvIKrJL8bC/oBwalBQ/owhiOY
w92VIpfEAlH9wxJTi9xMK3jz6VxaRauZh32LSnJ56HdCL2GE3tGBl/uT6O9AVgN9Oe6Eq5TyLeO3
qdIbk5A4rsCK3xLX3x6CvPRe6ts3XJOX4cPv/+plqdEXN4Ma5sdpJmMOaDsaR49c8XA4D7L4kQg/
Nw9z3m/uB1X+k6cqr4RzQD+51pOoiJFQfDxZhTnLchI4eUjkGvYuIPnZ0PUfaaj1rOB2UCEOPE4B
BMLtqb6EHplUqXk4ll/ns3SYGACl3nEKMP+leLxh9dOM1MUmOop+9kScEaFy4ZIwfrASLmQ4ms0F
NWB4eu+Wrwb37bHz7fTWy7oSArvi8BTHKe+BdwdpZCjKZiSrWpMkRFJWXSPTpn3jcJmiyKe5bbhS
sFSiTpykWBm+X3htzzMLqAipp4zuCdu00FqIt1e7KbjQAuwKWz1fg4s1ZCxICkILoF6yYPrsWOgl
kgyfAPs/3zAROZfPDBwwR/KR9nxe6vIJxl62/nyYARJ6T70VCNhoAIQlpKGeAHiqheJhsrg9H4uR
7KCT/yhVPGQOVMo8yjOsridO0+sexzAD6f+0RsixwZE6B8klxIX5fwHdufkbP4rCDsf2gkdrU19h
kVuMQzosglJmoVXD5U4niC3vV/7PranJ2t3poviBKE+yalJwQ5/TYkW+aaIQ768lfD7uAgsUOVj0
t9UvGNQuGK1y+rl75a77KqfLivogB8a16LpB+xipB6LBDGUNQ8wfGXVMPB7+9QYb2QP9a6aIFoD/
DNalyep5hk2SOEtxEX0JVJjkJdt3Ybx8pLi5OgbjOuloLNHiEOrdAO7q35xifbI/Cekf2H87tJk5
rbSil2Pq3rvMzobUHH3WbU751xN0dhoTTvE4iQWwZz5PNtZnrwd/u4HxGr+zC/C4Zz21G+S/S+5O
L8SDBtPY7P65VPdWPhOZ+sR/wsUwrP8OcSjZXZOyDod+5vpV31/O5EXu6/ivZsK9F4uj7PbosxKU
cXoE6N0igTrbaAiofga8eiZEzB3a69KXHei9C8eV1h3z/FjcyKaA4+moE4t7Drtq+biL0Us/H9hj
T0jsfT5s6TxJhKo3jV603O+PjJtRBM3w5BtEMxM12cCY1JwSOQ4NCh6aVuntXC+bIuTfDNu+/UVF
eTgfKnGNUdoUy0Bd8ja+GGRz3+ye9f+T2GPPnjA7CJtFBOrJrb5UokN1UN7iELMNtSPomlDH+71f
uFFy/LBuPwumFP7/Hmg9OLWBHpXYL72VAi4fwRTrZH9L1wow2d14zekzY9Ezalgnu+9UWouDqboT
/0oXsPWESfDDxOMb1B6dXsXVtm+OHjl3E5enBKpNKcTpQQa37gIMtYyJpaLrsHJiJoYK1GzH/pj4
BKAojRy6C9VdwNpcFrojHPKn+4so96n8Z/bc5DkRzhtKirm8xKBz0PJL+yZooPM3TJfWd8QNeEkS
F0ofuVwSBCiF2+PedDt5WSF+Ck7fGWSYyMZStWY8CynwKAmKd9bazvcpZJO59v87uTjIVszOwlK1
mMW8jN4hFsM0f7F8MOuKf45SWlZC11SpUMccUOJl/pIJx9WEv7QdfdS1y0i7qSVqr8hKGRdkETDl
xSTLPJtfI/xQLeURCiK+h6SRwdYGV6SHuDL2RvrX/YZUxYM+FpF284md3nte/O9QztBigX5Uz/iI
POVi8vXra/8f9vr74ld/YUHofeBGVWShhHCGchBb/BeX/OAtRabqNZ/pOLeGhS2oJx29IJpu3y6m
NjLUy1WpzncXwSedke+Y0Qntyr2QwXv7i4ZeDt12YhxGi0ik2idognKq11MG1W0p5x5IR7zDXEwk
/UAfQqNK1ac/u56vmaF+8oH4KoKrpnmo3aYHsWgq0ApmuwXja0v7oDH9KcKvK6TSB0j55MfPh0L+
GyomVdRH4t00Ijbz0J81/EtYUm9jCblcllw/WnvSg1BtJsFa0cYJb2Iqi80i4KTkKJDdvZic5+9X
cXysOAHb5G6bkQu9MZAhjsENsYA2LFem9tE9j0WEvFGyo4S/l6kwfuUwV1rlHPMUg79/eMMFBnHc
nVaQeYDvXXSQteqjVkCJHDWuuv9rVe3r/g2RSGkwEjpviHB2cX2n2xdUc705ym64dzhiqirMY+D5
AeBYtuV85SPOTZ1jrdwJkDgc656JChndvnRkYhi9/SndD4kQfdiroxse0/KclizrMANAscUumWwl
S2y5u/X7m09QfIf3gAAzzBA7ISGTkNqYRqhjsBvV9z4Fz+rnvB+6lGkDgJXLJAzDNl3GfomYGEwT
V4jF6HafjqDWv7oqkONwztcG3v/+MeONlsRtnGpJq+A5wpaNsDYfo1avm1WmcPSHW9X7JG9DGz94
FvocWaR+7jsaCyuHk02fauJlFDlS8eFigOXGuM9+LvZFFq6KQKNh5fYI2qHRMZW/4V+KerafYOYf
/FHAqPGY6l8+ZAptommV1Q8spIsgAlFm3a3OmMrWxkvdvxAYIE6eNqqJptUJi/WAGeQjkEZmxCzr
BOZ3iiq1YTvcL0PcmCHG6w5NvGGdK2JG3k4aZhTbBIaO59s8M5gN34TzYL0x7OnGTQcUo4ehYiHc
nuS6hAJaxIKLA/Z/1bxuz80PVa81q7qxmfo5UJAyhV0wlJFFeWqUmorAEjpi+7I4vcxML0Tbm2mP
8rNvyR6OTwflKMIdaU4AkyDjAOnX1TN73jla70owCto2P0t3vaeGxVfA60ZjmrqP1/renj3ckKxw
vFOGU4HjBWNxy7xbZVKvsb5k655aJjkKZvQwPnAFEtxJaajSh8EL65OgJ09AYEDL13Pmf0QYNgB+
Q6Dr/u6ux1yB3dfxSVEZqgK4pZbZgHNT9a/uofNnYLAdkK5Qtw67w8LuZIPE6UArI1Q5COvkdykx
5AOfiz5rqPK0HwlzX6mG17q548bXFrWuB6H53f2ljx03iOfDyHuqczd2ttYs8Z7uWwSvP50y8FDu
7/z/2ExG6BDz/io1ics6SM4S5SNxkH3pRGnhW8oBEj5DlKbfvuVMCA8dDUEMZygJj3SQvXZzsng1
mIml7dhZRbq0Dgw6ypgXJOmaGoi5wvoDrYq67aQvlh5P+8El2ANXLhP420784cXLToToeGMug1E6
w7dCb5NNyvu+/GutMi3V0vredzT7w06NJLbubTZTtElFtJWf0Ze0vIj5qsg9qPM6ztdhTzmbxAVp
cbmrF4zr0Xpl7XeWM5k9SRuN3cM8Ky5uL1aMtxfkajXQGgaagB9PXIBlgo2OV9eqSM5H2SyebgYX
o68gdFpM6DvCnjvHt5xkrTkkxacJkl1wsuT+nVD9Rkqxqu8KDxxSebas9oD6bBYI+Z7albZlPdFR
bZegkku6/HH24rSD2G/qVKZcC0TN0+yCYKx2q7qfVq89sQktN/pyqDQxDL+HGUuj/GPdMKLkhleF
CDWiDM1ckmBYyyyXpEv6o5G/oNKX23j+9M01rvTzueG7Irqz5jRUpmFEcgGZkMLzFUcLyYxH1M5/
c8EXVHLaFDsO949SQueVm6UW0HwUJMQXH4CCohoVnUHopAhqR74fsunWligSMdgsXfxD70nuC5Ne
VZszxrVty3xGEKL2wrGE3V7fVkoNG8RkLm72i80NmqdgtzKRRfXjZoYq0I9aDae0+O4cpzJigPRJ
+upWJR8dpO5i2lI91Uv3IvlXjwGoY2p5y2dtSDiCg6lp3aTsKyD77b7W6B4WhL/aSLYNkBk4MDwk
570irjHZtTX3RMMG5vBRT18TN3amDP/UeQePqdJkx7UBtfAdbaM0wBeUUoozjUG+ns6DwDwqrq2H
BudDm6/1RO3jtEftmaiIXljpxb4YSJmwr5O1I5ZNaMDfTb8MvrA/I5mFphqR7QtX2ZLSVob3NcAv
32UdefhsIcXAINJpWsTDFlFFtVc8fRUlVvzgalDWTjSEwI5yJ2a4TbLDs1HlTTBalLU8acnzy8Sw
fCKL2IOVi3eAO/WjrByKVUmK23HmJrponx6JE+06ftjzLijEkX1/2Jtu/7mEccGSHN22XBZF+UtE
mf6UqxBkEzqHpQVbp7+mG7EL5L2G2M30xJ9YhGT+MdJy04USYJ9cdj1zPjzjPgwgIFNXyGO1yH9N
fLadAFGInuW6lD4+laMoz7zalVStecnc/jmWJxT1LN7DfZEBNXov2lt7E3+vwRxdsaVbiey/I1vb
jrVrL8JWTpc3YX1fgFQxqlfZBJCrLOchSNrXcTE2wSW46TrQu+quCPNUWcsMLbYRtgfyAcn/oXW7
jT/G89XlSd3Ut5Hfs+I7Q0Vp0seTFy3uqnkynrvQASBRe4EN42VLr7DS7LJlY+zrjBokfaR3heM/
1R3oud7Xsd8ABlflF48tq11hMiH8INNhiE889mB/48X3G68w95uUfDogOvVdwWyKm6Y7DLUq0r86
W0SGiHzh2ydgU4WiYAa7JCOWVBqQ84NFnjn94Cjj0epCUkuqmO1f1dQefEzNZhnmEoVqEYj3gept
GwpzKY6qChndWWrpAksB+nQP0VdMOGtNxT5d5gkT9BvzN1uCn/5T64uqU0NIVrNgvvvObgUu/G0I
PNJChIH5Gy9wsr017zs1PSVJ2U8/iBtpUTyNdLOFk/8FKk/9ESh+csdnSgJd8caVPo8Q9EERp+n3
/7fyv+WDvXxAa2lfmWxnEA1OzRLiaNRnrjCp5cpj9PYdSiIjT/hur90GEJUMA8uAwZsFE0nQLTGC
adMiYaf4ULIDXuhuMqFGOt72/z4NIuIb3cvI1OmWaii7lXxXfNxoeiG4JpEaHhuVpKkM0hly2ZVM
dR5GD/t7lOGxYVnCxZfT4LjX7JurzJsMNys7jZ49efFAPs5xGXpd5Sb1wU6vR4jSUE6rSZptyaPb
aqsjzKfQvXrRT8r+1nlc9rHI9ghGICoiOiVYjqfKIVHwpe2Y+qTNzIpdyEJovy000g7+dPtpeT82
0xfakyIeCCoqTuGQqiVgv6/Y0pt9FUan0D4ThGimZcZECmAcYNs5nKdUBaQPcxn49JvJnycSc8Sk
DUPv4JmSXSpoxesQLqUitCeGEH0UtIpFIIaCyELCs6LXMdFO1d9DEHRF0OBgv5Oq6eVOCtDg6ufS
qvbvhrWniX3jzvCaCT1SGAOOT+qScHsM+rNirLxvvFu6w64YqJCIx2cOziEYJD2Zj9KjWqOR43A0
YnTdNOjMQTdFmM0RiIDCZRHtgynB5hQQBsV1QqzFeAbBZZlZ8IU32V1p5HCxSQ1CSU+Nw71/0mZH
Z8M5O4WohLOjVw5kXaBsPu3sTERWhJiTPupEXiVzlxibVd2U4f+pcVHnWoRt4zQyxf/37/6P6+u6
OzOjoHwRA3DAKGvDFCpWhPe7i2H5tZGs0l0RwozpMb4p9zcsP3C1/M2yo4cmcDi7rpYlPUynOX1q
KwCRQWsprZYgyNLB2WcFlhn/BDSydud+Ttbt6t5SnYVdoqhP5+1JApU7QwgiYxc/DiYH+fSoqdQ+
dOvc7XWl7FvtfiCDTi4M7gzDM09nM6xUFYATWCPUqFCzAt2sgFNRo/zaSsLApQefCYuzf5ojdWAK
Tmuh7O0pGh0IIHtOqBt2W34qVpAtNsqMQTQjC3Pc/xeK4imU/CJnq2FF03/+oo7CIbPuiUIpIFzv
Q67bZf56rBnhkJVWUdKjd149Xrv4hbI2niAxjwMr1TPKptdPlSMN5+k3yuGMZOIuU0iI5xZiQF/T
8ho8G8AJ3UZgVV+02K4Dkw8c8g36306xW2+JCOD6KXC1eT6IUByX7+dLCxqiG+V2oik03UJicXYg
k0zm0hlCm+U7QidAlLmssgMRC37J335R1JMVrJay2dS4DL9Wkx2NciQeFJXJc90KOcXWfjMLfOLg
itMI00PBefubDl0Oziod/slPict2rM7CbCSMXLbNOszJ0N4FeY2xEk+QR7JRwnmTjyd+WOXKlwE2
dqydJsDUR+BktcPL6zEinPF0YLSW4g7yvPOqejXlRd1yNmBNg/xJlw451eFRMbT7hoAhhoaAVrAg
N4w2KzjjlpbT+GGu/i4WVeeDMdMapk5eb5oX22d2xMHgeoSZZN7+7RNOMroqQkqSTvYsRXMq/73J
oYl92yuurE2wvHhgjANMhl8ePWA1Mnlt/0376Z48hi+/9jBNf/DeO5SY5Mfme2dgWnbbE2nSIMBw
zTDgYnjXFgBkePaCqatdMDUVlTMNp7LAlzU7+WV9/sGz2/FfYN1ecrkCB2ejizTog8OuDzfAPqrn
+NSKq6iPGDFqaAbUWOwJU02OlSET8X8KaNp2+PfUEOaTiYHWlfQwmRzOADIU9A3vAFBRRkvB7V58
dorVFDBdK8J630YZgCFWoYBVQrMrMPpkd5D1CeVDYCCFWQJOGvaNvQffuQ4ydAW3R8iGfXrMh7WS
pyj+4NrriodoRFFxteaJcbFQueh9JqnQwz7ZpT4fjMcmCpX0pdN6dHADoySxdyOhpklGcXRgbxZK
+jFHrx2FiinBhRw6Xu+9c+2GkPQP4idyrtZZOOYPFVURuT4ANvJaRtJ7pqe46V4PgE+eNiuypBN/
93FBCh7fittXeC7+ocyij0RW2kzeZW4PFBTfioBMd0EjBPfzwgUA8OdiSUVqrNxyOCkcynxor2Hy
SKaDavmN4gGXjbJdx/i14Ps3Sr9gtKd4iy21pC/sasUdMbPtBgZQiY/CuHLjdfzo78EMLroclcDO
fpgS7jaNmBfN4k1C37mdAujVmWovXuxxyVajQ/V0Im39Kc7jwdgT/oBkVqL8+j7aYzmPHDxixSCX
lB76ct8yA+E22yzqJEC6gUKtJulOK9JnaH0y6wOhwjTB5d8jsQYJ9g7xFzx5hy2KLfOczK6Uk4Q4
+L3vgImT7dKerPeGV1N2nfk1FYMqylPiXZWCQYR5PNnyyONI6lBwoVXv8xd28nnt8+wmtG7uR+ia
6RUYVoT1v2fXWIbVr9+OhINKjxEDySaEVd+XCdMGTjYWrXGn5oxEFJY4HKaUOK7THOt0lw7jZm80
i53LpuY/8wK3w/DDXO0pW6fcdReyc1hfWRtDGAN2+AzRu5lXDpWAeo8xJiZLx7XJeSMdWHnbPfD5
4rGvtIhkhpvgTwAGpG+GrtjUj3Hnu0o1pjUxAK5/YeDmxe3eURr4SQdj76HsSqpNnR047Z2lxcuA
/CFZPbvdT8LnJcePPKblLJ6egmXRT+bxqtBaNTpzKEshOfikxilWUR2+toLiXmi+Fd5Za9rh/XAz
NxjjAGBUL7mJpeY5Kz+3TaOBkX2wXP9Pitv0W4l9+zsOfpe575zVOHWIQ858+5QD+Lhze046KCOc
tFrqm1qxXWij9ZK9MnPpFct1O2yDg8rbQ2Q/yUwivQC+sgFLrj/9B+ZE3l/SdOIm/1vBLUqV9Vwp
WOHI34Rxt1AtP8C4431v1epH3rGbeyMWg8HCtXc/EWa7C6rIJXT6roZvdW8ie846oHbUWOuLlCB2
X7FazzQnvHTe5i+DlaKrqe6oVBL2W4oCltXxP9pwSnoI7snEDvDAR9S2jTXjbNoxDhFIUVigSxdK
u9ElbetBB9nexJAu49Pb81cfnK7U2HTOMOSju7EoOnWUR5DIsK0GfDTkb38TBteZWwNqZFSR3VFx
wav1Lq5OLoJoEYyg60KN8O2awsl/uB646qV4/4Q18qsQ4JF/J5r+Xqkg/4N8YBfq1folYgE0bJBK
uJhHXF7tkYIMRZLuSrSOqEPuPRjxZFJHga6UeofzR74BYpZX6gS14cCB/CkUOByv0kMHlktjndYW
A7tYEgvgT/KpMklu4IdASin5QEWMkAmmq9zS3V/Bmn2JQRk002MzVw9+XLmzU+wO6WISnhNEU7nZ
Ddb6+GT1h5Rd54EpN8mnqJXoB2q1rY8lvH+C82oTxSNNDkzhyZOGUwhPvHBVYVvR/u4cqle6lSk3
uNXjk2CvpCMd2odTd70oXJKPlGKMpbtqjuqeu7hcL5SM1qLl+cac2VfHI8elqe4FxqanpkR1yfWH
+ZLMzI0A2ff0Hu9foaeK6dbhiSuOsM9nS/SbE9AQM8guozOySJu9XcrHisZpbdFhUeGlpJzMh4Pm
nTv6KI+/4nPuuZSc80et3CVnMH0dNvMguiUyYcX/rrfbOOxPMU/cdvj7yutddV5LuDZCJV5cdIAd
zUsRlTw2OTwnTvCQEg4f8UCvEpRiMyvgQmPHqaoIdLlMaU9nVqL/Ap7UmHG67nEl+Vyb1YJY4x/M
puhjXOUcurbMGlMSl/BeOPx+VcHsYfq7GmHgaVwbb+9tLNsVLZtjL2tYjNAAhkAx4M22sogMxIar
r7ZcG4YaGgpRW7SSQH8Y1S8lzsHg+/xWe4eQACUMNwwte+EFYZ5DfxqOZVy05Z1bCH8GMTHXKZuy
/gELJ+zb+yV/7PX6nGElEiXGLOSJyUd2VETbOAEHyrXmJM0uc3AvdYwKVTH2z4hQ+jQb1XmIVAM5
fWrGNgOkdSh/wNzKRBdxOD76xH4KzF4WQtulZ7nZB7U9LLIByWf9vdIuKwhXIT7rxMWhzD6zBwFS
EvY9I3DSmd06Q3vEw1a5c+DDqVTvVl8PoATjsXRYF/b6dJwCvz/YiPlbPPD7d4PKXOuE/OMmKSqO
O688muqtbh150vipHaqfl0LVzUghrJIkFVJVuD/KCKCANmWDOYE0nJGMprThVTAPt0GaFycLnnbA
Wq0ZZ0nIAY+9k7o2v9+JVg9pb4ayzKOKeC1yWAUo/DFhVwI5GerU7SYBQEmK41sAhApkHVKVjavV
ETsIwhg9hmanxT+NvYcoInkuDYV95Y9xHq0OlKxtmD0G+PKHRGstuo6dpDmFCpkXfr7r98Z0ED+5
yag7Bamc1uedajqFFOtYVOSiO2NlTnBP2poNH5E864DYtfLAqq8ZGrdeU/iU9Ep9HL3ok5dWpoHx
Ff1uYcAwWivZwGGuC7U7uPu+9hLtLRDfDLnJ96u3/qiCNOxow1lS+hR8lnUGqSxNhq7ac3pgPwdE
TAZvZVRc39dYoleFSyLUN/GJIh1s9AHscB4zz6lJfLE1ltQgeOOtxGIV+QabYma01h6SIEbX+Dcw
1z/Lsrbr2fPJGwWVzygkMb/6CeGzU0ONoHR5Rc/tRAuqqPX+WppY5RY7UwFnG8MPMVjA70ur3dgs
9F/FgN3OK7OUiDKGdBgJFSbo6WHc3OTdLDo0+H7LcDZ1df88N9C5L+U/rBg+GCicKVrpfafNtdQ1
cLWizpLiqSryYJmUSOvcCyboZ4exgF2XCsRbmAJ1uaBKjePVvC9rJXtNHjro+gJqFMhZEuF4GLUc
AfXAraINV6BO3WdkpXJZ9TbmJKan384wgksdd7+xEWKtvs3F3gqSS2VxnpN/KuKgZnuKhVKVx9ts
VFtRd0yMr5IMpSTu3KnSmwRZQv1AhBUfPQ8AXx3M1Ed/ccBqjkCcHdY1dOJbWpPoMjorVnSts1Mj
KPz2PJH79AZ5eOWVjmlIRvGS0Q6o4mOIycbR7FHX67q/bkVR3MGxL+Y+T+eSG5gEk+T6B+oDI46H
c/hGC6SAwqYUGYWvOseu8+txtv363bHGJ3IWYIzj6ny9OHrLaU1Ex/2l/IuK3yT7RmRvD0O4UkTQ
nAh1W9YBJreOGXePyZ8nu4flSwioQS9uwcKuJEG3AWyazDo1tUHSQcmJdmwPA96ODCfZyPxPJnp3
1iNyiRHt67/jX+CVgkgBwdM8PKaG2LXL+9mdf+M4byETWn7WHJnKH2H0wKzbDGBFtcuV4omwO8mH
9e1wxGerEUdZdLXTIvqkFHMokeJZNT1jMxb5qneu8s84defL/RtbYb+4FDXAwpeRggWskfWG+x2q
u537IrSG5Ij3ZtAKdHCEhrgS5V6x0Ceitmd+ZzNoYUrSwheJzx9LBrOhw2okvNFiP4UJs2tUOPV3
ginRDAdk7yUnrZDCJEIbAOUI/D7m5QsVYNbF8cEHrNVgsEdaA+/XyM8wz1doTdRL++yliEpcXEXG
akAgMdKiiMhhIb350nNjDIKtQqG+ETr3n6yHtwH1xbfbeVkYgLMN+nCAo1SItOhMmHIF56RvQxuI
hkZGdgo+6ZXtHPv85P7E1Fgc2GeIPq7/Tipdlm0BgImevp4uIwxVwr2wv9lPupPrGi2PfgwIXuUB
5q3CoJZwca5/0YDWDB0GoxfAfZ06UL2qx52cwMRSc96xo+kV++g3OqudkvsCpoPPSH2XOXz5vNhg
htzvjX+IdwxLdOhSzKAckd5sqwJUSasyAvOlt1TOlul7ZSyZLdsgxasfuXloOT4pLclheWNtyrW0
6+1O+5g8ErXTO315CGQW0aR3HR2u6VKDhRPEnEVC5DqwbfnwbPmGxe5uVYMU0Fdx/EtO8OBU66Bw
sKYiVR4eGxlqDdJXYSL85zdb0SlXiTEVmTp0LcIFoipJTUKNMZO63Q/ZycUyMJpXrh6Q6WiDQp08
2GxUB/SVOHyaxGtvIe0nk8cZFUb+UgFupttekbGo375ZT/cZZMpVAhl8/+j8EOm5O62wDlqJB1ew
SRYeQtk4qomxp3SXgL++poVN0T8gFzXyQqF/FAn6+hO6xXmv7vUBEcssV9u/mWJ8KwJDYjCh81G2
s/aEorWyP0JZgfFoWJ3z+fgH0Sj6ic/KLa4gTLRyRWm3eEGe0vBcIPeOWAIBF1dvtGPVxqJQoKEP
f+9kCCySTWm/d53DZ+7iO3ntrbijyj8ZBMcsnBfSixAsVhcpYQMPLp/qn74jnS+NB+aUCUmgDLZh
Q78kc+OWoWkoSZxEd7+KeNazncLEgVmojH57LtdhD//+fGvjU7cJOzQHb+L+b5yuoKkAg2RwXt/8
RraCdSHNumu9V8B3OUvPc8VvbBg7/YFW8G3RpT8NfZajVSBAZd/uQg19Eruv6Nty918H5fKZ+vlS
7Bh8zc99kmUu4rbaqeDx48324Tv5sCo4zFzokY40YnfnyXSox0V+Y2QzfUF7AV74ZVZMnQXMALPM
uGK8WBvhxyU/5mKuJoer+nf12mGpdjdIpZrHUtWrkWwTOjxGrrW52lloOBg8Wj41gH6N9RG+702m
yMonCLvZ2/rwVZFL32p93cWoUJbkzyBMrTfpsGLF+xT3Ahy3zcLGa93UeiBBAzjcSdyYbj1RX4wl
luO0xOBodgSHCQv6YZOrXMH6XvqB/NAPLKgqyNo8ME59+NqVQysBfljstL5QAALVCGEli4zSdDP8
oKqBIpMadiDwN9IB5y4+wfyxu54Gyk43zQKujr3oniZRWfISfPjPmtyBSGWlhNq0wrwFwsU5Urfv
HWahSgj0PfhxlfcxJ+a93kqTYQCon11+jDhUNOfZOgbxMHQw+sTsmnPmcxC1NnxNzJlugzKT3WCq
WjF7NGaxqXZFOO+ug8RZ2qfJfo9CnzhsSlMMEMDNSJ6QcF8RVl2BVAAyVNA+pdQIOq5Kk+eBa71E
ToTXxoIwBDMevgvJ/jCn/iizpQfREpeitvn6maophhZuPv1xZiPV3H4OzHpjx24z13MxQhr4Jele
morG9dyaA2FThiWCHnNF1WSgRR5IAwndVez15e8oFplBxhBJhdMbiiD6tgsEPQ0aREhWmDyyrnoe
Xcc1zJ1yfY7jCr2uV1fbVB8ya5MSeeuR5mGCLN1p/V31syD6CNUCPLfIfeAXjSwl/HoGP5vQ/zjO
YFN0yM0GRcu9IQwJvkN8mRQLWaZs05KSX5hlRn2axV61LlcVRz30gFFLoIC5YB5lqYp8lFgM+XL4
WO5qH7kDVOp0exHGpDtSdlrT+/+7euAVTSgh5hsDQPt/gcNAXAOzzSF624GekSzIuWmoh1Sp35B6
9d7wwabH24fSKLSipbI8aIr/fGyHRoXoKg9RQtJ5k7TMkyoo5VJW9uOCEFAQw/yV14PtwsK6sQhz
uTx5t8Qye0Ykx/d8q3MM4Keobu49y77lcTtGfNlQf0FawJs39+dIUO+Lbd7wGuoXSh8yXXJ/GNCc
wWiKFQ0nYP3cjAcfWCqVZqzHD1Uzi+avYBlZsO/5dG1Ieta+XZKvlnZUxYqXUi88tGnpHRY3YDfb
jaIJ25vhqEVR7y9BTGJbespI3Up2RYMYQVbp/GoH0yl8JfjYUjAk32CBq8+QcWPVUKM36rnapixM
/U2Zlt2ROabNxfkUljDv2zGfPsuDhFmrQAMp82SF+cheR96dlCFcL0gQUxdwT2LrpNFsPNkhzrgc
YbQKcslYf/J3SvROG1YjWTQSD+TDv9540r3Enz3qF6DfDaurx9qRE1ZExJ+oQFJwcsGl8ZgJmCH1
7AkMiy6E5BAXPGxqPF9/o9q8+AI1mKyY4otEdmIoTBH2f0A0dF7DU7+Q3B4F7XxuzFfQ++z5DpI/
/+fgu42gb7Z8wuAGw6wPrQTUt+2eKuNcEyKhcAv0DbCxMrebYvNjyP8/+cM10nBeueVDm0x1JPE2
KTcxrbokljFK81AhATID8BcvI7D86jDRL2TBJTQBSWTPv9xxa47e4bU5U/V0wGonx95FfqzFV8r2
t+e9vwWTHtmAvvma7FVQJt0ux6T2p/4wwrKKM7eeGVmAc7WfinmRI1tGLw9vMPr17rhfay3Ha8se
iimpyWmwwuCxSEif3/+iF9jjvdut/W2VXU73XBj1h9PGb79q0u6uge2Nz1WvWi2CUNY192u3OkzS
peYrEzOBONJSkZG/uyboQzLeCU8W6v8HngKumwGEJuh9A1Tnux/KPYX3OHm3QrhXQaQcpBDCCSGH
DE/YnWLFALdP0aCTXs5GfJSCltX7S6OIjIC/AR0rwlaZW6M6A9n/x9bwZmnCHvCs9nKw1xtTGEwH
S65oDP5AFKxqGPrnm4gY4SbJlOD27YN+z4m6St6TU/gl07/qgmpPYlWwAuj49uWT3M6KgTKhs9A3
a+xIJ4wTIkpJiYi92rmJl/P73E3WxJzgdkrG4LuWKvcRGeAxwWH0hHvxctvcuA9yabYV93w6eL8l
H3pNaKWicRsPeRKb+E3ZZShlotTPMvYAIyxrHFD+uiNphwzk/EedMa+nKt1voRW0u1BU3qP9mU11
sdokdkxg64bVjnlu3xzQf3m5ioxZFNV4t0RvnfyzCAHWYdUbmxefxt7/IVABUq6pGkAwvgc8URy1
Rq5YLAHQQeu61FZHavvsobxnfZ81/wcZ4Y5kDWnqmTvmzyeD9AY7ckgo8fbNmIeaVGehEo/LktWU
5UrWBMi9txDypfIgVOK079FhDlu9KDNb8459LDtaULV99eL0Al49afkOqSS+fI3qTjMdejTUMQiu
m6QC9oFsfizLWW54OJ16WJT25xrziQGayUoU2Q6a0z4LGkEPzUgVzq7+QX9F0Vkizq4XfYajh5+0
9crjSi7ebHCgWZp7R/+qjepjaFaBnl42V2xKvB8M3WUriORAyVgDzdH5Z5YfXWud0FLsx1ENQ06r
HlvyhQ5n+ZnFHbBlXUSpbQsY5ed+i07wKD49KIAv1HZD3ZRCE7IkvQeH6Fljxv4uPCsvo022XOIu
tkmjjKrsHautMdJ/7WYTTxch7dJHnTWepcPxAAXh3VaFdwFjCLQKervbsWiL/TWftuLcBHccIG0E
xmxRfKOS6qj3L8WwQ7ne8KdpRf756QrrIQDYlwCX5DO1zYpJgupT/IOZYjrYbxy74Sk17RlhLYsf
Yb9bK6W5pZRWeHh+0BGQoozp6ZAouZPrrJQLeB95uVy9/ma8PdoWRDVy4Gebu2FiJsD+Rh6KicIt
ABdR1//8/MSD/cKHd98zQ3BUhyBh6IhZtB1iLkx2mM/VS4n7xPx9ayCPKCRN/FtGEjA8YsFQFLYE
zI0QQGqcec7TBZPem9voxtVHrD62jbO96pGVTJCvcBGVIGFUN0ikDfqNI3dHUy0Cesp271lYAwNf
0XL055tv7jjlCviShLQQubJUmq4ftzEzrV2XvuJwHfjc+LGbMOO7zucyvT6mhlss+u2bVyRfJOpt
VMktJGgg7kqcAwpibAPYTQME+qawPmSBwRQlDXqh5tzB8aOdZXf6GKCuzbyOVg7Cn1KvKnhenRnU
zMFi2jEdWq/wcnl8N0WOm2/Bq7suuSeokYDfYaH+bMMONSFNNLRJabB3ji8Mn9sUCuEq+TokTdCn
2dtTpWBP+8JlVySlLGwoB+C0nn5CT75tatoGbUopd1maTcaQrOY5Ay5dZWEAG/oKLaiqwXSFDfly
X2S8dMmtdhZ4Jw3F2Eeo777EKjHulUKF+mvAB2VyVwoGVtwTGkj3ZXDoYDVNjbXSBssRulDLg8GG
RTtORJFzb3GIFvVuso73LlaDVsidPFe31pCkm4IQB9xOSsuN85i0u+cuzz77/rfibvaaS576AIls
C341Tlr7DQUmv99GGhzRxmdBk/sAeS0uNFGGjIoIU8EmdXQ5P59splM+7Oopw5XQirRqO9VPXvwt
ikaBaSpsOli7kyQ2JxM7mOl1OsHx7VPrGQRHGG8I8ZS5PRVNjzX0+8aQR6OILT5oLZZUQR34QYuH
o9l5XYESn27gqhIMQqsav/a80j3eMJihC+nxYcPkNI2Au4xVmwpl9wl4aW8yfsLN/lHn1/JiwG33
qJ2Lg77IIkn3HFf9oLc9lmLed8LcN/20oChR5af/g/li48f2Jxla6fXIQcJU2T0ZBzzzgoZnGjiV
vzG0j9d+I+WGQVNjWuDWAkx62RmkhwNFo1pdR2lOKOE1uhuERM4W3KcTlgG/FrCEa9ugzT41bZju
b5GFRXrACbs+N/LUtZ/JIxwT2jY/J2421JFim4+Np12VdG/FGPSEtbqeFe6aB+NFTBeyeaYqF/r+
7r7sYnf55lHw2CP5cZZduF6NXppubfRzkwfVpKMDniPG2hDj3HO0tfTLTFulf38jvriUx4T/5RuU
P7Ju8cGn692vIxK6qmLVWoSpjyr8ZoH6SnkCy8Uk1RuCx0A0uGnyDd9iDqCdJG/WTeH3UbnHjF58
aq0XLwbzA1RHUYdDxAGjRFnhA7nczgBAK7ZDeIUrDPU71VjgOn153C5pb7A4D9iXpEOfhHI+Icoi
WdjHxGzmG3hTaNzMRQ5420N+O6aKWlL0CZLM4WnClamKNziwFg8UiHnKR+UayEzkW60cwWHCBRsC
HbWn7DAxpGt0CH+bxMqDY/wU0aFNqt+ANyiTnTAD+HnE3dmJXYzZK5c1rHHJ0ZuYGxPiXokTJ8ax
9oUZhuW44KUcFSiYLSguGhBSEN+dIjjp80pg2W66wGWvyFCOcO8ycLy9jhPwEtirkrTL9taHiQwc
Qsh43n1dffkAGuXOtbhMS0fGnpecdX73JXxeEGA+tvAwEERkP9HHmOcKYQpcGvyN2s/3HMQUtQs7
CLLqTI4+FUWbmel5EcDWCovQTJd1ZG+ddTiA5ZO5Xw/b20/ByQpdgkXfOQiDOlvrowrKvSGvp2GJ
WsgKKS7L4DR+iPMzX00T4l/ZUFCHzWlYTAxhYhdr6n1oNsNhhKtx2kS0feGwONdlrKbgf+Gb6h/R
DEz+nxKksPup0oHU+qYklWQPX2gpGzDgo3WeLxXScwRrZr3IVg0gRarfZuyDSRnYut0pF8u/8gVp
YA8sy6dGHePRCT8MIL07ljP3kdGX2FY8J4+m8Ltf8E0xOacopvv/KVkRqY5FJ0qgPOsdkpTQxfB+
zIgRitK+L4DhHpa26wXOcztMstFWjDmzPEFfk+J+FrU+INOWW08cfGrjUQBylye7QYILkFAiUNG0
ygNfGxTYFG6gDDG1hLQ5V8W312Zx3EUblKu+c1olM3kn9giJ2Rv56aZ0R0xxc5FK6GAYoB1pwshK
Ey/WKfc2qculFbNv+HIY/ncik72kL7J4Gng983fso46xfdU/KAtI7A/Mckijgebz6eyXA0g2zJb9
tA/bQP6sOmMq6gC1A+hVlygYGLvCklqeTOzQdIK/pdI/xgDrtF/lc7HtArpouCRaMuwBjfzfTf+F
msy6ZIT8CUfhglAKx+L+xstN8U8XDwM+GMaq9zh9D94Ied0piAzXaL3U2dPJqS73PS5lKg3Wd4eK
nMzdq7ZXCOSIatqkc5UzUQG47Npb5muCmYFoqPY0GrWK3xoJE9vqjnDMFxzd3eFbPXzwzmIYYWz/
1v1CIGBh15V7iXSSJpNHFX4jsPsUA3WAeqPFS+cgZF3AB/THm+gwQR6WXS8Ij7/HFjPs4BOqJxPH
RpFCPl0S9LRu/oVYYTzp+q+KxihZ8a2gA0s7e/W1LqYcbClKalangcbmUBQoqP2fwAPMWXQ99YeT
6qb9Y7LGwSai8wVRjddE5IamVq3QcuL2HFr/5W5lhfo4mKo5aDWmBjEacgI+6AedRGkaH3HA4ybY
K12E8mfQ9/MnmAA4BxvdMvkEaeGjb6CeEccNeyemh/6z85jo7czUYySmudHiwSpG8q5Q9eH3yWNp
6IS7e9S1cNFojgqQOQf02GNSs44ngKe3iwM2+BSQE/Z88QUZuwKVwevMV5luVhLuv0dw/5E+BK7v
I8DTG9JmjwnHNeZwI2WR9H4ndLOQBq+mTR6Ap5BRjzoXDUcu+Em1kj1fkOHPF1JzqNBXneSiL8lS
YHg6nVvofVwtwMkhB8DWCCVXweame4XsTcU5b0TqTnf9XmC+0KBpJLODbHDjb5A/UgrOV9tg7K4a
CnoFaIdTLu/1KfTCBKLgLYBMEkcu9+SRlorpC306sa1X9yHoIhj/1Q5Wq7jpxNOL7EI1Tsq3gM9C
lsGt/5tw0xONQrY6497Zdghb8KZ9XeGSkQxlh70Bh5Pr6DAZNGlKnIpGGfWeLrpAS3KJbMX1BOeM
25XngivuouUfpwaHUqqAzmMnyzmHk7JTKJnK0Gh9YkNQ3HMwW9W1Ccww8jBhH9SkslH8kWQFXTdc
MWPXQ3Ln03nV5xPWQUc83dP75ytFZjXOO3xEsZ76XZrMIbSK10Q2uZQvErMC7fMZjHqSmT2pmWcR
fPDXo5oO70M5UFvKB1b2w1UOpkdI9dvBqq6aNeDC1XK4+ZO/nMqcqxPGp5eDC+UV3oAiMJ6xEkEe
uGXFVO9H0QVZhvJ7KZFJJmpnXPeGUqE6SsOMde44P7YLto0R0eS8QDbCgw0m7vm0RSTJFHzn5MGk
XcVJPLI3E3wE/r7TVh0PgHzU5cUtvFLntejOFgc1M8e2hqpromwM/kUE8Uy0wEwzLTn3I7wUxt4f
bnYf8THcVdnC3CYqm6b5T8PhCy9i50+BwGt39vVJfFBzBExLah8muKmbEdUIR8aFL3KqbAlCR77s
kWJVn3U2JUt7wjffSrxOxfq8ZyGuRueerrDRYAsmeCFPxz3IxrhOVuFJNpMBj2NqblkwaIwRElYi
4N2zdUPo2M776Q9D89Drgzapqsg1Nqo4/taFjSlhjDLUkq2cbfaQRCw6hf3TYea4IUFe1eV+tqXA
lti+Zii3Cq5gyIegA8al/1JG2aZsDJKlR0nVlwZzlA6ThWlDiP0iE6044H/NfKgP86giMiEEeuEB
plG6Z7ZB/k2Smr4aRhOY8vxXCsbF48xkaDJOHSmbB9Ak0F0GYPLuiJiPfcAL/jm6ura0P4HIFKIt
Bx/BlJ8iLGMn8XH8NzXetsKYkeKYU8VQSKM64AShZnAr7j5/vg2EfYJ4rj135VucleraQDDLxgS8
pZWH5o7GK3xYWWsVQryfukpcTaPFJUI8tEqfd3taZLw4gevL/yJtllGPyAjlCwD7KbBu+GR7+eAi
vfO2EfdUZuwrvjOdQiIyCKo14gTkYqcPnI+jw4Yong8CnLHnhi5yVHPiUxn5IKNSj2R4e3XbLydI
qFJiXIW5N1i+RpqpkKD1lTMXx75FArYyPJDsS2a/37Dp08qME1SpwqjGdbdCoeJO36O8fERepKcI
l4PjMJejR1LIO0qiZWyNd8UKceTQDHu8A3a5Yf8MdHUGnF3ighisGBTa17nESmpl9eqmklEUVb22
s1aSzXWiu98ky7I+2E3CVZJ5DmEHDzKjiXlYdjA/shv/zzKA7jESpl0Jc9O8XQt4nUY8Zzl8fnAE
LWSW6miPdWc0K6NTyqWuRwvh57bw8MtN2dQdlYs7Val23OvsPSk7PQQ54T0SAbDy+o7FNTsdpDRO
Zd8BBa0gH+z201OUPMYiSUSw+bURkOhey8cv26IiC7D46GS1dtqITS9BeDKJBfH3gHdRbEGA1Dwz
3yyYMkmu9iBq2LjdygmSaxfncXV8S1DodaWGQ4W/xVDN2skWxov7TkeWRIHRWFjcAziVisDjt7GG
q1G3YLURmWWlnyw3JsRhNPvhu7aCZfc68iuyEaHfEKfnusiCbhxrvtRF9qfJ7fUU6cXqqT5r9cPV
jq7WzaDo4Z2gkJ7U7O3iiRyu0+nDlI6575cExLepgrcy1oITzFGAQvZLYt/psSGhFYJg6j2YJGv9
q40Yiv83e/k3MoWIJyAMHyCwXTEJ0Obb7wSePutydi9EWPaG8mJjDQYOQtEm6c4M/aIalwMs+LJh
HhcAQCMfuX2xahnaURhjnik5rliSp1KJXCzTUt1c2CDDmV6PRlPpaI98+39Jq27gB7TNXVRFobXA
VhwnQtYvWZwE6KcqOYyjH0KcmwlKWKHd9W4UBbDewiL9SwKihsIdiuT+fuYfLPk7Lbm5lGaIFrj6
hz06kPWJHasyKXoGr6tY7+mBSCEcUoA1uyqOu+G5rYF+4QscUsaGnnd/FF8hAztIn0RkaV7BdBze
OJcWdnFmjoZq+gsM+lGpfagUC/1qaIoeMzhpaVhvckZaE4waq8V2E5XaSW7QpOgzbF3pHJ8IC5wx
li8vALYAP9QWChehKWviOfjkXADzOeIxtIzCo2vEKWI6wT3IQGxUlx/BDTtvT6viafne1YvEr6qE
r+9llk5vD1uVry61ErT/s6fSjfaqxT5nU1aOvuFXzY+mEMEP6I79D9APqyc9k6iwrpnzhMxwnKxL
EVdjmz4xr4gYemMi26vQXLNzKJ2of8VKrl9zQa1vzjT7JXFGpfc9S8iPA5ivQY6JwibCkBBLmvpi
ZGY4D8TmPpO0P19xKFPpZEWaLp8ioJDac5v3BVvFzl/eGrN6AUSHbtm4WQD20wqvomY/JhfUZ4ov
sj1EjZKPYhbeqjSP18hD7XT62iBE3hWDmDTUN+mydVW4aoFdS7VenBNs2fsdj6vL1j5TllQfuxrt
HewcHo3wYWgkN6xLXsJo+P9l5pgOnwSZsB3Nt/efawxSeVT2bGtCAurf7lcv9hHDC92zOABkdpDI
MYU/XrSfd0OTd1PUFYFHQCUKloi1WwooiwLnUXwsKvzVWrWzWa1Jz5E0jb4JZzs02cQRkyhIbaeR
EvJZ/blkcRAWdzcw9Kw5vqJyost0s88CWJApjseWZ36enM9xMsaxu2Z5VEa+yupe1PlKIt4c5CB+
8nd9U0p6oOJnyKfad3KOk4pOkIDHvsxBRIq7/bu2gsc76qRrYl5owjsoi5HB5D4F/HecnMR+SY5N
m+ZFRXYY5i3u9tOKCdNj2Ld+CHvC0L92jYoBIYc5njnPtTcDR2yCboEsEvH/rba4dCYjBoHVH0GQ
PI3xt3vdfoP6RDid2vb54MAX1pM79iWgj5gLWdFEleDTjY8Trz0caqr55AgaDmpi4Smy36B2H2hq
Nrx2sjWbAzefjLcVTVEVpCJU0+96hjeJUIzfY60jF80m52Zc+PXRRtJ2ACbe89igt0irAnRvVxig
UmJ03xiZz6RwUDFmof9i3/SRjZNHa/gWE2ZDyrRu3cjlqkxJzjioAu3woeuezNIQI4mckKqfA94I
65ioKjIZSPKDICzpOcl3z9mvl+lirJ+Y1k2aHy3CXQGgrW7j6CgKSWKgIapP2IK0u/hsW8AzfBDh
c6GnAr24Qx2SZ3VExZcvSW/lvZr+FP7eesx58mcMH6XRTyRvsE6+J8681uu8onsKjSwYklUJO9+7
zSNxy76MfNt/qWYXfb1/ZITuEhQQfZYuNY2grHHGnqPub3z9xPYnokCmN4CXop3PBv2DHMEF8OXJ
TL3Q9gc+m2jDIrmxE4CQUtA7isO16KhqykeZlWN+F/ae+sx3g+48cGl/SzHjplHj8MVXvRG8fRUP
YZtFJ9fNy0QTwZOcLjBvThbBQTZD5UVAy3ZpQRgBRi+mhVUa7xKQBcYHmzXIS7hHHR+vPQ2prNG1
VqQMIpTqtXhJ7QBxuF+KrI6hrpyS8auCcYJMw4iYIgpyA/iJ0ump13goRTXwY0HokOB2j5HUccDc
WV7NXYNZt/tLEDekw4zTnvEp5XJ29JwToPTub+qb80O0Qp4NVrzWQbPpn3LTu4E2aBy1OigN4gFd
UWYXptmgcmuJmHQpnf+/Gb1Q86FJKHlJnZev3VwKxDJvIFuaCv3s9xC7cQ2Ha35UdLODfg/TSAbe
4TZaHd26Zpk03vPjbOj/ZFX5P6TQ+4op8XL8U2LR7XFE56TUivtJXRo/zbp0O7LpMhbTF2ypPGer
r3aLm9YEz/bk4duF0oiqbLvRVh7dNgddCQiMq3mqOELoGlpda7RLGHLPhWHxNTFEYILlWV854PfM
lMIz+QLEBxUjYB38vpAngv3PeMD54fcTNa3Jmp465k9IDzAX56gcdfzkxfp+iUySvy+Z5JcTCgAM
mLHUrCZTt527fnry1MEVmdtodz7kcclqImb/xYi3z9ZHZVsrNKIjqZFBiIYG9O1jUbgQhzLZ+YrG
fmArQRH7I0Sgt06wmHaG/9bRd7Jbwz/+geZl+lKPi1NtB9mB5PXUtlBSCDrq2H7UmAA6MVWGyga0
vKPQzfuzdZR+CsS+0h6VaEfbOOqNavuYnvDpct04TExmjqVNEGN3ieRCGn0wD/2ZfXh47wpu9NVt
i9b51TNUke5HGgs+qF+oJxadhbouo0O+AuHYMTAg4CkPBlFGmEoNjczZ9rq0aRRAGNF0fCtgZcN+
Co76s7qjLTmW8N9wBnLusskWkzk0U5BONeO/YxligNFJb15z3iybGT/+WdtyYVcxcOY2fmFZqiTl
k7z3ZkcuzJcCQECdjHrkarZEfJDwlhtckerNM2xGCBuqdAJ3mqWjBzflW9ajJYfxpFDde6dx5Ic+
gave0DIGOkX1MwSnnuwXvRTh4p/a+HuPMFu3gDI8Vw5Ug7VfllpfylROEr+LVsW0m7tJRTq03JR0
A5zbF7Q0B0lhwnrqxdut3KcTxB9EbFIX80pE+TN98UYugz4O9J5h5Zh+K18NuEGmJNv9gJ5Pra/j
at4b2r9lHG4VicXz7Fdy3WBOZjAEh9usgBSnKOy81gywE3qstlb7p9K0eyjER+bWOvnDP+1aFaoO
w2pPWeXQV05qhEpu4EgFxsZks606HlG3jV8/z/i5/4K2zp3f71hyh2vmjiHHXrEE+mIUQt9bqWoP
RpLRRFISpdOGluHdbQj++x+CgAr1q9zhLjC1zJbkWXvrhvP5B4zlWPFs5xeje6wr7nRYTQg9AOhV
txjpJ3zH78T6nzQmuXYFtEeLYsTtnOF3TTZ9e4+UjIg94NRYYuYvZUMcO/bR/LTYcx4iisbs+K4w
O8pDgzRf5WiXUzvXbRJHVeKI/Wt5XLg4xwe6dq1H7ea1UMou4qpAWfRIrg+EWTMm+v/PlFomP7Zd
CJco8+ldMKaWgqXyDwG6KhlhUHott49ilJX2N+I3fyOrSylFGvzbg7flFAOFL9NsDupL9/SofGHi
xym3gIU1neq6WXm8XwE0mpnXN7TkCkWxgjFV1Fq0R7RWnq6k/5+5QrrdoUYvrB1oFLnWSy3kRQw+
DQGCAPe+l/AihVRQ1RXVY7lTo5odSqPE53t5nVtFcC46+3sbmNjzY488a1HRQkvhxVzm3bOa/GzA
RMnwEqvXHd+PF8u6n8GyGtZtE3gHoibO+IEIcLKgjEaEsHiWew9dzEWOKZwsjU2PUhOLM3Ru2k7Q
CgN/1Y6VD7V9No4V24IsnuyYaKkPUBFH2lTCFvFpC9aAg3jzWyPf/Ry+1isM+Es9ULahbRyzf0uF
hvwPNPHOQFLBe90a2IYJ9o8XHm/AF/BV3w9rvNpkGqFN610HOJbudHxWpHa85RIerkKyqZvgJlm7
8y/VpWxRGJcJyNb4eVFuxpNCjoWIAzuxvZOX4qxCfj4vbAkqR96YHB2b6yyMMAve+ci69hAIvgfv
LVJB+FnB3j0kuDCGiss1i1EXpNJCo7AUDqM7sUrvbGjKO0Rya+Huhld5XTzLgjvO7pdsd86Teed3
Y6ney1/HGXTNBCmzaFppqgujOkl9aDLI9r7d9LMXmVTXNL7dOi7naFO2Jc07Y01UVMq7FJI6TBYz
ogtxvRiTn4M+zdThWCqgHbrPuSHpz8OzuA126DZuZ6D6Qq4SyX6oOtco9n/TWhy9pwQ9hi20BZ0M
j7PzWvvjNg8p8aPpFrJ80yKqNWvolJJjeWwhCHwqtBgPrrmYsA7MWPuhPC6bYsUR8SB24PAGF3+X
7PGTIx1RtV6iuIJy35bQ6Zv5rUoaUUoFGqP29AxxQ4Uyu8YVuNcAUrJ/4g11VukxK96FDWl4v/5s
RoHYXOILsIxC8FpN1MwomUIaXSDrrAxEjXA/4zEPAPM6/SIeNLMGnhvj4X5BbJQw5ZIeBADrlDZL
4PrEWpBQZJ2BK8M8UNTew3lE0uEJM++2S44/7FQSeRSMZtfvcBIzOMoXzWh6oLWRraHDxHVmTpGe
aIxoyyM1EbqJgLpBQmdEjwQvqVqbRjmmdFQHeYXzp21mMTr072QFJ8jKKSVUgg9txPH5CYFte6uO
5ZLCqFDF8kXNjS211oWqLdo27sR4WlVZdFvOj1ANmp65pYagcbjMsLezhqutDv/XrIda4ujjBBqF
rNNoXbmQi7hKChxeMMDStNTrGFDv/fH9RT6jov0w3JkLjzTSNSk6QIF58WHrmXKpe4GCRg2nvujA
S7hbjz8uIIupxlAV6X3M0PZJR+qOWM5ZA284CRlCB3mLIeLgTili0HFO9YzAG/1JeyQ2MRlgH8Ik
TVLCcZRi2wNHUpK7xS0l6wEASLtZIXuIK/MTFc7hpGTZS0qdZGK40/gD2UHO6CH/m18gNPDgTHh6
V8m+aKvzWIJZVOruf+NbG2MoP9xLo5MW2UHqN4zX8ZiTQIPRKd2HCGkoXGUSCy7mjDotRVm+AqNi
NfiXgpTCBk2vA5PKHsWMdmtvlsaQBN7kaWMok3HZNNAiCnZF5pVhhwQ35rU0TSmpzyBUd9iu0N/h
QBAV3XTplpKYUXinogdD00MpI53VeKS0ZTlgJyHuN6rfqfXcK/kHC0mgf+JLH6Z2ecsAbheDzN58
rD+Ya+NHcGnD9MCXEaiQtrG/UySFtRx+p0TW42zLphDMmVA57HtWoEp74MtbwwtZYlDw5cHJ878r
StUb7NIG7K9sMzRxZOXrPfLu+oNZ4E0bKIrcwkwuV4dxeOXz2KghdTh/eLvyTEMUPBIYSj3IxfO1
LgLPrjHtmpUHRlOdldtlLia7cjFoeai3FgGAvrGln4RmibwY/irBgesUkdy1DSyYYo7RvSUGTXuO
7sb0BWaJgh9LhLvbDrdaAlqGfD/twtSyFElc9U/FcrRlJVFdYUxQYC4vsY27mk+IdrQRJNRvcW+c
q4XKXDyvJ+YPLyd/qiXziuUW3CQU3aQer6Y6uGHqDS2YmNXvsYOI44E6jn5ptHiaw5csyDdnO9fS
69Xk+XnLT5xQCdgqY4b5VnEaJhc1GKQk3kN9OPXXqhDeSCVOWwmO2UZ68plVTUFHmjSjYCL1abPK
kkEeUO57REYByAXHYKs9uNruuXwX0/nngbs9Igy+Az0/wC8rF0sVQxMYZBgUl02UEhYQtm8/AzBu
EFIurY8WdH8znnIty0482SNRu44QjTmhjwoLDWhDCAAb0tRjiwAjdjBDzKKwjhqoZ6fKroejvIDW
abtEMh2VHcsqBXCUWJvIx0c+N853tQbR2dpLMYy6vVe3hKexer8KDPkeDYiJwkTk+az1Knxdm4bh
ul0mcZmmq6nrxfERBlJ/eFoAIRF5nEo5QL5X3VNjYVRfK3iKpmyEejWrlZjMXpoLvLMm50tfhNgO
HRdIgQqh6flBlI+AAvaqermIzI/yPJTNZHrjhDPaYSRH2HD0ynAgWv5WmZDZpQ/SqED+/SALlrug
n6gcqu6jZWbTh/kxHhkd0MxLf+nHd8MhhTUSVvE53dPk4/OyeWGAh+nyOH8NVwwOaf0TEApBMfCV
+vA3MW6UkPnKdwFQSxro52GP6f4vW0EQWL7bmkOlJZ5uGtYAZUnH/qzadWpZDHeHQHg3wd2T/vnm
BudUVNGNF2rWRaIe9w8F58zDAwMU0JOI4cHIKbU0tRWucVcaYxODWSiNrHfvUfX78PLJf3milNo/
+NT3J+XXcpS3fPszsJah6gSolMujwO1brrEuxHCTDH+EcVH4rdVTkQGoYWEVnTaCzj8wDFaDhW4N
WMXVu1Oz9hUDehZVTe4jZsTWNuUHnNjP2RF/2rt79jSMDf9xwxlxabag1EJYKAHW6TcgCViWtLzZ
z+V/tQBZn6TPMRHX8pnVdqkMaOQlAQlDcBKYUY9aXpf9ZCKN2fuE5ff5tEW6dBLDmN7lmcCDtO0R
IiqexU5T4wL8WfBLQlurVAgOLu00u0gIJpQkgqvCxN8JG9Bhsq7DGITcheE31zfJ1dScqNRBuyEC
vrf64FpwTWzxs6I4OCX+4Zg+iWnLkXLov9wYSWiIj1LihJiUH4HYUKIsYimFxyU0jGQtdHl+zhLC
seZLBMr0uyoZJs771vc8bXjkjK+DuaJfnV0pmRJyXcWml7CGV+nrazwDJRAxnuqL9+OPoQByVD3Y
oNeC6DHUXRvygHELosymJzl1oy/Boi+Msq8sDtjkfYifVnxnR9BzBn0ZveXW9CebvMjbBtV+2OTh
OH+unMIh2cTzwc8n0bkRxxZX+7UQyXon6VfeGpspfCf70b7r81lSb7i2LRS0o1oTR4PSNLJyTO9p
MW92KvADAJYmTe03WMcADa2yPMLgPausQWyOcfnm4tU484c688WFKQtumZF6KJ65EELXDt7CD7Q/
8U0YA4dOcu/+20ZhwgBtkST9sLBnidTfBUy7/Dehh1wwsgmSe3+vxJxFHBNT3IXS99LCEg97z/So
gx+kqtEB90Nrds30MrV09U9iQCLj6YFS6YJ2mchIsNI7948zIG8y4F36LbVYI8sPZP/zpQBTHv1T
YDDKxQtM6WNmH4JLlyarQrFJxOmDzOqAyPnjXVLSgswpBcRYEkgS2LidJlMkPsf3la23TZRMgeiv
zbP77uzlFEjxK+IKzV0P27TLgpHHXGxSqAZ+bx26IFY6gIyO6mQZ92F47m2Z+PI9Am7fSVgnltb7
obpw8iL99dc8i2jZ9slWjT4HDKrOqlhGjjNrVJSSTdZDIXL58Ir4y28xO02dtDbQlPCgVyT98vTW
o6R+a4SulsHTtag+EXy5+xRVeqJdJC11KTnDSEY7eC3CWv7D6Ei1pO3O0AT7NSk19LevmCu/dXcy
Ai9O6+CXbn3U+MkL5bBa/GCwXgQeQbkl6LSIOg7jtFE72iLMkqrF8EaDa8qk13RrVkNa8y1lL76Q
6CoProAB1KGHxxGNYJ8eV2Jrd0Z/xw0Cve0R5j2dl0W5RbdqNf3gK0jdpUFkZysPt28EhS3uqIQB
ygBX+UE9iU5qy9QG+lvwu1zlv4uDZYvDhLozbqORlgBlsKbK1FczUw7+R33IGpDMds90pUyTXChe
wclWpAdz9RVrlRPAUO2GDAhk/qrOXjdVpuF3j7nbZN7j1NGR8fpne5VG4VTg33Qh9UhNwfDuMfNH
qK1GypOt1iF/Hsn8VLolgLFAj2VwTHjPlaV2cODW/sAWjyVR+ffFwQ8W8y6ndrUFvPL1n4CVrQiq
aRtoHWX5Ii1bpsSzKM71WGx8jAKbQQKXGAfD6JCJZ1pATzL/ckoDF00T3SkNtJgkwXdPBmByttbQ
LuMcvdH3KRM6ncrIxcDw/p1pXGFf4XxWQOFcpbpOhliDFk7o1q1eIfT4uB+kGqP5rNUX2tmRzgIt
vXZb5Ws13k5FT7LZXOzQY+0e/ga8StJDWRtzuKVrgCyCTI2+1lLZGMQ0igtjDTXp+jtLxxGAWn1Y
jy8FjCvrM4eWIS+mTnsT4S01R08q+IkvTFX2ERLNj5L0PZFzNc7QL25vGPbsexoxK8hx55XeHxVH
GHxToXcBa2o7vOf0aALxlMb8kbVWZ0XW2jBkKTC1HnKe7u+T/mgtFgHQNevvSkMS0mZeOSjZSSyO
BgGe++SNpe/o9dXgXHBJJieB3IuC6kr4WrtmHbLpY7lzfkSRJZAuD4BAyx2yzhd7401ZioWGOnfc
s4l/mvgjyFPzqvQqMVj0wh6MpzFrkL5iaKhMJbWrSZlM+jOzX2m7boamAYjBwU2X2R9M7lSAdfL9
8qtl4tJ8T8kPWMVxd9/16P1PoG7WjbHKWTPfOCTrIRSWlZ+X1FsQQwpCQrL1dDA1NRpDwJvdmL27
JVEYHTgmsaO05YgpmF8+gbn+DBV4ypfp01v6A8fb2w7sy7gSht5GQs7q0HYs/FhiaIgMfGjJAtLB
EHP3fOqQrfOxz/M6nPQXi0NRI32Gzo4EQHUIYxZ8TTvaXriMKkwb1waZyjrUV+t8HmUa17j20GJW
E/D8Fu8KUEjd1jjD49AA5K81uIB9hhuz2cjmyeHC9sEehEpJL127mAj4mcJHoaIwXsS+ksj3VuKi
zwqPcDlzHBmqMQVl6Mkt74krb0nmwF72X8cLO9IJ+pWrTPhuuIrBr7lqNqMO/qwvEb84D74CDBvw
vd8WnIvvwk4HFdnDNtepSaTHzQoeYJUHSaGQCk5xfBmnLk1y0StYCYY9jmPyoneWxYZjc7zfjHL8
+VGNC9VDtFIav81JBP51aUP+GRHKJKj1SWCEe29vlkao7+9+nD8l8TdvhlvZ+wSlBAxWKnjc4fui
SolVKlOMOti8I7WpyY+4m56HUl92KAyNxsYqWaWbl01VhYw49U615gaJbotpFzpFa6ntV2GFh1KK
5KHlVODG14t2442RxRz7+GZ04ygw2c+lEWgjSSL9udcRnIhI0Qm+bQSsxErRZHTO7DkS1eqhVi+t
bWJrUh+euwumC92Hk9SRUrHv+ONQS799pLuiz9ni/cLimHal8z/pnkLmM3EZQnOfaPp84NiiHoOp
C2nNZVaAY2cUKtq9w/O3P8Mk0ztMPBquzQW1Bga5t4opfQwy2azSwSqv3IOiKoedB6ea9FVpfpq2
GGR6m7Ztq0xoBud9mQ5hMlw1cKXt+1T/tU4sXC0xC97ius5PGggeTO7Rf6BW3Q3LODD29I1o0h2w
4rCftnl9J0YSb0ICyKbF7gTFcCx0Y9r2f9NdhHC2J/DQFlP0avm3tfcKf4R8DNyXquoDnHUCJkBV
xLIzCMwiYCrAl5uwAuZ7WbWw6pa+RU+UM+39Kre9Zi9N0Xabkai8h5pCJlU9nM7Y78ZUna7ipjPz
zYvwi8prYW49/dcY9ewqUFWlVSCt6fF1Uww/eqIa0Ol+JNrO329T8qrGrmBlacJk5YQpjeEHxoI8
pwFfKDNTXwqgtFNVHtNgH/OaJG3qfHfNzh4GCH7lTljj/aiAFbUx5JLEovzhV1b92UDJAAHx44Ta
5vY6eBfoI7hXQgLMLpCw+znr7icX+RqrpFPI/M+Y0fSEkz4QTWOOQC0egBnpDfe/LqG1Vv/NyLLw
JaUlYKenHm51O7FFkQMPGT9j0Cyam6b+5ZIZ6CLKlB9Z4JwRvh0vjxyYc7o4cRLD0AHz7vMV3uRA
/e+qJPgO1awYNDQjMZ16VAoRUYXdLWT3ADp1ksoUQImlpdQw2mu9vX35iW0KV7D4CBw5383NXpeq
PN8BLxSXzaiZKgdvnp8kkcxvzv/HGy5GjhBaOKmIJYxBqZtYDecA5YV5Abs1sdoH58qtHKNSzbLc
jabY0Ae+qY5LVYm8me/Vt/cJ7swE/yDSZ30CIKqqn74opwyyUln0qDZy8FenKpfHVuPORWhiG9eV
oAd+F08zsMMMvDFZVdKkTJCIHIf+rd5meYUiPmnR5OHATI+lRfjVftI0ZMLf9GBP8cjGQaT5Wvsf
1KjgfcOd7DM1ATA0BEPXl/hnnEtpo29R7hETARA0fgaRLKuqHhebMq7na8aU3vv6jVKXL734c83P
YM2IeX38Zc1xKDeDJkQaevF19D0UUsKfCs3uM0PasbYJxS17UByby891+5jMVQFL9fhAqbYQx1xw
GMSWOz21pwt93NECLF4t1yQuVCUnf0+dyGeLjqtKlMvg0Z55/Dpdr3oQqiGalnOEAapaSSX9bFHl
/EusJQU2/MaMiSt5SbqbJid772KZlDI0T9AL30WZFEWDd4SKGM9t35P+FBVixdU648xXLGadPlAZ
juOw8BxI9GmyYik/ddUmxTX07Wo34tIj9f6VJvzechq2kS4SvghySg8XoK2/HrOCAA2GlcWz2z9b
mYLYAXauj5UUvMa+nK1zez+1xl6wXMeTEhDTETv2H/Br7K50CJrrx6XcB3XxCwMMVMMp9oRisbij
h5dkyBtrbZYZEw4P7Rl70mg4k1dLuCXGAILylzjVeCDo4QyWkbgHLLHkZmVMa9+E5tNJGGIwHNWh
nZbqWFJKAtVjOJi7IZX0haWq36uhMpG5d+eTUYXl0Gd9K5M3LoVyh7klylW3BsuiU0QMZ0j3wzvm
2Ust9qunwe6CIZgTsxrWJp0WAYITTspD7nG8j5tatG4mMKSQYje7eF5eekYoqFzhjih6RgHWbPiu
6I/aRky/jTV4hwt4KUoHIGDvDSyl5nh/cuNH/p23e99j/70yhVrzqcq25ygPdwuK6A0vzJvSQIUF
SMuTiEj+HKQZldOE1WkzpnLe/R14iSbvT4UacCvdRMy6gPANVgBt1SCYNKe1xlECLymghQ6+0Irk
zQEVm+UzaE8XZaILawUX9kySVt4BzH9cSaDOLrxf7B3Oy5JSx21421D61Glnfpd5UUn9krWaUAW8
FNwwlBKZ95Ov+e4rHtB/Q08GPUCgi4JffU/H1O0BfWh3j+7EuiIBNsNt0A7l83zDotmsbvN+IEge
xCePWEmTVT+8CfrFX5QisvNvWYCI74XLUM5QOWUc98/illceWGr8ztWN7DV4EwS8cTBcysXatUfX
ZtbssfdHrYjoC8usx+tE1GVT18LBcNR21q6603bN3WtYFr3iB1t1Neqbx3jBJZrOJ0mkXfqxB4HC
/V8fhaDSr/22s4S89AOU1o6Tn8p/V/UAPsccUlwnMaafUBy9Kp73rzFO8CXHHJb42tqB2NQELYAo
ji0AdMyyDic3dhoWBj4EVHoGPkzyPwBKYya4DcyxDPFv8Z2dIZg4zDNxOaT87RQzMvhojPvIIFLG
y4+XALVLiMTSghRzbOi+ZiWGDAaV6v+Hy7AzgrxZJiDkw6XrIsUUENPsMrySwBlhm0iHR9Pu3Q35
Q1ls+X0cgbv1sWLk4Ma2CueKjyPgEmmAmj7CgE0uQibGNFksOi4wJIwLvEIJJcIvveixFCLWzPZT
1QLAF6pmUsBeosAZArwDSuTu/Owtkpj9jurQkL5WfEQwxbGg5eJIQysiYOS3WfDmeoJZc7uhGJ36
YXhjbC+/aBkiNIbYDc/0Tvu1kHc4KFBFq7FS/L2YpNtENi6sR63t4pc6J+Rw0AolfjcNZrnr5Pvi
e64r1EDgLk8Ry3lwT9qNml5dUCie4URW4UJkSh93BiIH0cydpkt213M9zkN2SE2gmgSM/5Teirvj
uAun12PNLbbDO06cxGAVryrCD3540e1qyASmHuBVWqri3W6wuOn+Il+rQm1nGH8jU5TLK5k3LK8F
ADn5UADbDxqcMlP11dYtkDUSZAnxtduh33o7YDB/P79lFxhmAOg6D5qDCM8kfcuHSKuVk5Fwmh14
nhY1mlXYlEsCcbS9dWdhldoNSqJewbGAjaa9/Vy2bytH6nYmXprjXgYYbcjqGbKcBCqBztH4+Wl5
Yd6jZv36En4zLYMWJ/0FbSrOzEVjgTaUWwhPX//xwTmLUFtEYUdpgG/N5cmX02ifr37HOxvPGmyV
LSpSiRKg/FRoWLhyJOceg6+v/yraL2psti52BNYZ4bTl1/6YF7yVNVGdQ+pcdmaO33jVpBvrp7Qf
QiSn0fuuSicskgQa7Xs+ol9sY37CseTHHycyWZK5JE3264JrD1rd0WAmAMYwNpXEaKrqiBzMAcdE
jxTTQe088uNjyAnC3ZrCteoUnCtkHq12kahFJxuS17FbkLE+Weo2lP1h+wXc+aBy0YA9Oq+MivNN
9+FCxlc3h4RlZF9dvfxvgjy+BLSbDbBkCvC3Xd6C5rvDciyNT+jFMpLFgS2Xp4gMjK0qTQqumtO/
8oQikCdgYK8WQmrEe9hqH58K96RR/mV6/zKisS4rQ9H1bQYwACOrg2fuS04SEhtHnmAqE5u2d9Xb
yeoMH5cjfmKjiU3xty+cu7NqecBKcG1yIo0kQFEU2Dy98HNlkHrV3oez0SPaAiSn2016CugNJx64
XFCvbW8DRJ66pl3HMq2wdrHabik7atse2SzJnqYVnFZ0DWdvNjFYIQOtOFyPb3/ACve4cZffaGyz
Z6SpLMICuX1Q9mpj7n5a14qLIHf8KVHejijI9wZu9W12hZedVPAARDnxw6DQx2/HrCfs1RYchpp2
P0buhzigFGNXITzVDW07APP091XAyWDrJtiEFkaiC5UWtKmqlrAWV6WJ4HyGvKu5LjFTcYC2+oPl
XBM0QA+1WG6tZEfQNPRmIkI8v35wh00Nq7dhoMZ9wCVCaYSrlobpmJ+pqKrVJK4+W3Hatlixpi5g
48apRgJbtUJDHYBg6HCicXTiAzQZ/sOSUbvg7EfQaXTwXRnKybi9UTpgwxsae5oO/eAmfUaZSrMc
MzIjN66dHgMShQe4QhCF2FuOUK38/6yfe4wukiJVGrtUn8K1d6miR+Bdgn21jHli+3SHHIyHLwSl
DCvRy5QSQdNxoOkSLp44jyR7BIgBLcStg7TyHqXHcvYOem/0ycnoMLJ/tjU/qFcWYWbLs/fx2ZJl
CfZz79MRFgN3BR0+XOac+ZIS/2+PB1c3O1rviCR7rc17kJg1kqgbym1cfxO8rjE6awgGTYFuUlgb
1TY5yW9tafI5wFrc5b8NNX5w/BYxqEyGd7q/2ek/Wv9hsuIVP5tICEwLyZayvc5R+yMYBLMMKdDK
yc0OO7z/8Z1Q+3RGGE0PhEi5BnZWcdRAoWPBGj85BZUytsMND/2FXxzpNlwX7LA8eo6c5cbB07Z+
zYfajx3KeaG25iS4+TV6/7r6aO2ZqKa4MPFQrciP8ziDF727lnCVlXqBECzg/S6HSF0dmkQc8BV4
tytvC3lD0iEkAsHmk38jTTrDgufiTIv4OzWKo4N4SQc3SD3rDrJUOU0VShT4haWdwMtyxszjN9uT
Z4W3KR7npiG4BzuH2zH0LhNLgvBbBQrqIl7s/ueveyfhoftHoEstQp6H9jjBY86pHbdZ7Eu7MvoS
4wosmMz4LGTyhZiRbWEt4AilTqRyTFDGVW7UKPi8qXjVCVdVsm/x7z3SOKrTROGaCF/XrIR9Dwd+
GwlhgGOApAV3vAQYQQul6muZH8buKb6lbt24dlPGot7q1i+iVLgg6sU7tEHcVKHqJ6VbOuT3HYzQ
g0DeeF0IGGbpFpnCEJ+GAWVcjjT10vr00Tv/l09KphhU1WnEtopK/7M/QPK8m3tDjqDD4GLSNIZP
6vIfniIGr9fysScw3Ynd3dmI5Nl6l41sojoOIN1zOQpSNkxuR2v/BbzGcGrVtDouQxad6Fr5HLy/
0o74gZcrXu3agyeWwH//2gxSBNpk7h064UlOrzBA+qbEbsHF1O/abKcJUKCx7myf99R9w04m/bSs
Lz3+b5SUActMXtG7+uLzcLTZauvt5pgyhxRbqIyUHBg1ANpuVv8naBBGAbBCnEEcWjp38TkfbBTy
Qj3PZVN3KxVYbM5jSlHVi0T5N0WTg7tTAFTEfWXg64NIr5aiKTHx0UbS45JhPHiu/j4i3T8VHo2r
EtGiXxWgFyDVHzLNEGzq6WB4tSaWnUQhgZikgYiBzWsZ+kynIcqF1hc2hxpDZ7k7EvmjPifOMGVh
rXo9/UsJjqpas4NvunV7R4r4Tw9/YVBZjgVGyr1QdM0eQavH3te9xzk5x72xSfnjNIkHNQUwhkfu
tSbic9ls3431ui2ZINJ6u/E0MXRhINYhue5QWyUHB9ZAFFZP+SKRSn7BQ2JoJChBYiV/8tLFB6fl
rH6km+TE0oXkhpCOYil3TS4BvecGI1WBy0jfRvhjDoN1/HTjCYGwLcQGpZhqWpAPAFDUzWaQeskM
LY57IxBoxUEMKQ4o19UPuF6T9lZeQ1HVXuOBtjZhg2MH9dgzi6qU5uoMYlAMomUslrlu/JRySfqD
91wUG1iOu2TPTeLDZLe2V6uk8B5M+gMv7E3db+BcgD5xvRDNuj7yZ8xqNljS4v1hpw7zpuIqGbIs
gdU4TdomegG+oO7y9k8MHajD508hwj7ZKg0TMyNYiklelt/IxzPQYD0ZPDkVeiNq2ar7nD/5a8ZW
7FocggoSP4h35eKUO558usnMI7OhJjcQUxAJkuib2UxfeBdLXcXRRyi6HVBm0pe8MiyLy80DXo+G
5bwqixxoXQGv5rs/4sx4NqCgwEzWwftUhNhOZEZ/yN+0+2Mijpkw0IEE4WcdBaSNNxg4B1rvZJZ+
Dn4lWe5rRQg8qqSrPjX3udMixic7WfkyoWP6FzXSONEbipegaG07u430xbXoORhZKb6C9bG281Cp
hwlr96nyU6q+rnkNGBWqd9x+SZfkg+sRLJrX4wVCWZic+IMA4Ou8Nlr2S+ehk+5ou97eqqZr2jhs
Q32oU8j710frvfY8MNB9E6hhwJutZAlJ7jqzQP/b4vj/qZfXkz4Y6JNu8tJou35CiERTMTi735De
e32AQFokcL3F+8Lx8qh3nyXQHRs0/pvvygmHddK94W2M6+TQNrcg7ukuJWLOwyv9T4urCdXgAh2W
J6iXpa4GQt4Mio6HILdMwsAu3Q4e4gstiD8IBse378p4yUILtA6TvB3HTpCYXby6uHYF5nXZHJZz
P0AOA46lONPx+PaFR2COwjulS9SYoVDPoyEEqk5C0qXPsXchfxKFnvZ/mmgERXdBQRYD2FOFY5w6
GoeOltJ0j2tgeII+u42FKiDgVLmFcuf17RCLqwPgWQJymABu0eb9cNz5IOk00vb0sXOCXnTEkqjX
NsQU9pxikEPLtIqXvpV8C+GUJ9eHSULD7QR71EmKZwjNkpsdah1ekQhqJxr587O9LEqpd+N2eNhf
58h5mjiK39gMUC5uvhj1ngPZzr4W05IJsbswmgzmNXn7NnnJIHBzujbaNbMpqQh3rve0WOL5eWJX
gCUfV0Wtsu/h4nK2CQBk9weLll5NpT6H1QlBxClpxZb9FvEVfX8XyGw1xePo5ZsJ3XLW64agVySa
VvxNRyeoe5W0p9ZKDp0aCTD8acJlBi2/9BXlDkPJiJdDOnZC9xQ8RVbBP+7I6S3rR8RSkTIuJy6q
VMVyoMf2TBoTWaK71EzRjfiJpWrY3rq1nmufpszEGc4LawdUhy6sypCW/nk5wPB92plOJUVaZUsH
i1JwLnIuD6Eu+UoAI/EnSoYjb9eQtpKZzJvACiT34ob0VZkwtDBdonvEv/KBV5eUQpaYT76n22pw
b75hoe4X0ITXysLhuULMVC1hrWvlDZFs9cVJV4pc8q/+ka/EO3EQ1gbcpAorbxA4wEiSPMxh3094
oHTafSxWIxyk2ER/VsmA4atE6lfkDarXsjxFhlFpTNsRflAGhITS2wkS9IiGFW9EY5wSe7RX1RS1
G7WE1evlTcptYbzvokyqb0DXIpdAPGAavlkghgHHvfTlsS/8qK2q7b9Ob7K8kcj5EIGxIULTKSZk
1tcNlyxZ3ViHqGBzQAyVjGiHjQcWWrqZRoVPHEuU2dV5beohleZBPg9q8e6BBogeCUw5nZMAkWTr
l5woIvCaW3rRgESzv+rm/CFwJ3jpPfIQCtXRueLmUX4+9vHKe8DznV/8qZrX7ahKtsZ5C4EWa/Bo
rIVR1PcJ5vbEmL/RV90aWz0Hz4jJRhEUQpN+DpQ64/TuB/vo+UXkyLepKc7zEbpynHV0bijaxcs6
aAC9E52qxRzVxPxJlSmg3BO3O0l1CYp3XNnQQ5ZZEA6DAyLtEMzaajVdFwDk3Q+Ag+dcNdS7Wasl
jgnk/y8EgmR6pNU81iBP5ao06IzMfA3TWQP5V2dhroz3rsdYcq8ipyuwcummZkrEFNT+Ed8fPufC
ODBD1di01FR9w4hXY9F0BR80m0djI7Z5vr6hV/n4cl5haYPOOy75Vd+L4SGk/Ojc42DWxRx6YN6d
lCjx4r0jgNO7zrH6Rr1rUfdqDVAmdEnYd6Ecthp1Vw5pq98nO1+T+bw58V4rxpYacO9DsOv6TPWi
rrjxXXVlzEbaRxuLcsB/WG+pDWDH05RrZ1Ys5aKxOEus9siqS3BlVaqvnuW9GlSV3XcrJI4U8LB/
ijK88ZlUymLOPrbznG5hVtsJA10rFhVoYRuZYhyeD2M9aGlllVscti05RBqfLC9PoAICoUHCXBxV
cs1SjwQq5tDz+EXQX5PthUrtxOVk6rQr7lO9Q6MdYbusF8MTEBwiiavBrebNdTVdBVPHSaRYKb0b
daV3lnLfJB1M+yap4B/lFKUBMiXmNRMyCctd2xRGmDBf8SvP3IscKEz7jToh8DzEV73ktXFA2BAu
cGCulTpXOvLI7AhBRV7UNpNJJq6buE11H71aZ/hT+hDoqYIqwSSubWrXsXKZ7N/GmWjthmwegBqb
IbyJgDh/SW6kAuxWffVh6IW4xOR728nHrkrs0/1mhOuRpHKoO+4jDjNpYJO3yVkrP9+nW0olAVCH
XnPNep93gb3CM/Lh0bnwV0HQq0TklOxSd9+aAK5wHEBmhMPkBHHND4Drm1xz4781d4kI6AjooW/B
Us9kuYkzSLr56fYiK2BheMJ4BsI2gDTgQQIHg18Zajlimar92Roo8JY1OR2zbuyb4Z01wUTDYseD
pt9wSrPQ4GI7iCSr2CLzB+Juq4rEUsJbifIIoEXnzjqDKGxq6r3YPT014Fr8kGvFtuVq3JljCr/t
t65mIfWFYDpeW81BgfMgkijq9kH7ogw9Qv5YpcXK3OEhugXeuIxKoUsC9Lth/XiUU6hSse9z9WUT
scBDUbcdlGbB6xiYKZMHoI+3zGGMOQNnK8URuNaco4DKz9kqghfcNaiTThoK+JEt0fT6Fqo6+dy3
SQ3e6kzqPUr3atakJST1sZtTyMktWlCt2uUNftNpt5b/PISnmvIPzAJxyZMoPD23QWHZwmgyECZf
UiQejPPA+1+T5rg08/JM6AAgRaTUIlUSlOrTmgz5Xm5g0/bOuF4jHEnwx5KHv0LeWcDCujoS/pLD
H0GC4mFNeGDvi3gSQJ5zXTvrFI3zs+QXMzE4C9Kp3WpnRFA31GdhhYELOR5yy32WVqjs9AKoGTbf
1gVknXKJcBUvb5mU0ypt8W1LNZuj0ruk1jOyg1PevhfKqDDXAv8TuPQ5XdAy/BgObDqYblOCfsp0
YeXOXCHEXMXnesqA1+V99JUrLj+VJ4vnq69kMi4ckGI63e7vfQ/8SYza/WEGycdHmSNZvIaPBf/+
b8rvyiZ2PebXq0D2DkTvaDPEZ5DDStZSLJi9AlV+ZxibnsOXZHphRSTBE6EsGSrfYjPorrVYZTin
0Uy0HM0OtDdnqFjQ5xcfLExrcSO6zN8BC9x6EyXNZbdfkw3tVMXvRCbBcYkedvFCi3zJb8U9qcj2
ENnERmjgf1VsDFh4Q9JoDNv4v95KWOoxyXyN6mlg/LSjzRCbXyoMltP03pLhEnbNSmslasAnnCK5
4i+zofI4FGKE4g/kUCj+FNItJskJDZvF5CT227fUoKvBSDEOVpRiKr8C6rPcu6/4BEHapb/3nueS
lMiAROPFmDgsQIeLniz8kgzo8MVi8DHfs/jyvzhFxNTM7RZW1ACQD75XO3p0uGBxyXtsxs7nIlEt
lS+TmJDC8+zgYfC8+1IIFesMd5mNS9Ax5ph4ykHvGP+PCpltA8/HFyZKlwVKMZElgrSaBNzOwWGk
gaXYJDwGbNFF4RDYwRaDFKQKnVsZI58NO65u7sNkmkJzsqajeqQnqfH0xjaibRacd5pG/c/POANr
dh+YKjMMshNK0PoXzLgikj9ANIgfBxBbLOt1j60eYFpY8CRuFGEy/Pb8319sfzSJISqMatXSomro
5NQI0TPNRasTRVZ2HPokXEFM6iaqBUCE5TqWmg6THjHlv5RqAW2wzdu3c/ejIwjntWFR7A27HUOv
20ul+Jb4TtDHVsZfvRGMcZtK4fKCGA056ACMtwkAomOIWjDF4McZ/5K0TRiv+/EoOhyOui4bsn5U
bwRQsELhuZ3i7HoNXbDOkd58tvxQXcJ1ykbLkVU6Xvk7JkgbUZ4iw0lRk83NmYw3GcCW6oZPzD+i
3ofxgzKGz+bWZT519hCl5YIYZnCH6TER+VZkdF5cLRM0VX1Wmg+NubviUZF6ZJJlhYEwcBpevwit
MMUfTZMfsRqZ4UGxZCROiZ1d85eQ5f5YE+UhEsayTtDwuLrpDqpsFoPo6zIZZUgOcem89ZBYzIMb
XXTmvnjbWMPPyya/Xb7LXrh9MLcVDzmK700SVq3DE0z74UKoQvbgOusN8UCamOF0QKdl86DINTEe
JeO32ERKhkavj96zKD+e1NgMk3aieIhrOhHBkv9nBrmbH5phpSk1S/RLtictbZOjNyuiFY+M80qY
DC3oUanSLvzoAmXRniDALPJNsypMaknBr4v/OxRR0kefPM+EoEdyzgwsPcmYKYp85pzzB/l5n2wT
fNenCtN4JbARaW0qJRm/sY8mNhaIXEKHpYYwqXQzseRlfGHud9OaTdEjUqeiXMEO77Aj/LWqd0Ib
5MBgZPBr/9fnLQpGma0FJC4PoUcDOKfZwP68YGrBIwFznOo4Jp1KhoJsMN+kQit94d/d3F99imWN
cOkWeYc+VCO5g/NtuKUvKmhRoksLkviEe5Ab8rI58xgBenqh5WZRmwgDQ830PZ0f+G728lj78SmK
1x95Eevl7IbEoWrH/Ez9Ggi04WNSDIRMKYlLrVIfmyTk7HiEpty9N/oR8djel3ZOqnwUx2HfHkbD
EDdEuGzuFCGXwOjFnvaIXaXMwooz8IE7nw0g5MKRiW+lr5hwtxcEOl3HW0xj30ugSkJmUjyGIG27
/qphwkiz51KTYBmwsQJNsVIuhmstgxOJFcFFSKpeeq7uTIKbNZ7Z2Wnd2ga2mnFfn7/KndLAWUmN
32o6flBCEGeGaUcVyiVlrx4TSeN6lg/+zhuWnetCJbESuUQYNztonmQQZfB9ceKDawxBVV6NJeqZ
g5gHnrWLFbmOCa8pwrCEiDed7D5cAqN06hm/GOyRpFPlnajcHz6kd2we8XX2/aUm4PRK7deBAF+o
+V79z9tOn5pz4EzEg6FJhbdqlbxlD370D1JHoSvLLlUF8Y8jWojwF8WfDXB64uWGaeOP/cLnZDhp
+1Xp3gc5phSNsjpXmWg+rIcsD8KhsZqZayitvfg8jAwzGq6cD6mQWY2GgjQcQY9+cSvaxshavoA7
pj0iIZUgnN6iQR+LGBDlnjBSfC/WSs9ObdNIPh6t+w2qh237CxAdEOJv5LXXlRPuRXLSaehv13lV
Csy3rcvVroBlGC77UeBZ+RtlXO3dUMHJwf9+pk9Rc+1GAotnO1Gqrhnqqsq7T1qrdxIAUX/DaCGi
Wv9PODE3VUporg1S+8X+TuIo9Fx85o+9Ju7Oms+g0hiuvaVkJ74hAOinKD/6JifADeO4W4AR0kzN
8dfSdWSJ92eKMYhWyKyLWVEKaP10/WULa5JiQl85CP6/DzPTcHPI9hbEjYf9biPke9e1jHnw5OCh
muzkR+QD8Ez2nWDp3BQXvk49sDGoh303YU2UzjxuZXzbsoV3MffDHgVcHsxZjQKHpbkfdSgpFFFm
Hl2jFK279ooBlWmrAznmnT0qX3zfLQK++GDYvwflRlXD6FX2E9y+b8iSaUQ4eHGbIdf6x0j69Wyh
18RlcqCTln/pnhAdvHL0qxQyyegc2jD5mecUgKb2myLozzOeyAFX4rAEGLHEgreX/0rMv7Jcwchq
u12FIay8WZNvah/wbtrfRwUOuR2RkAimqFVsEbQNk8/pilpVbrNly483j5f9YP4faTbBtjU6wFNy
51FJ+o/M457qh1r1Ount9ojQx94SR+kn3yKsAQRmQN2RkjX/lF3yx7P53yG8pMM3++JheJ6Y5mYv
8St9QavGU7tuT+9f2PKvLBCTSxIbSKj3eye2a8CiixHrbFJtA+imujS8vP+9UL0XBnC9BWdCzqd8
5TMhHCMpcKRDSVCGpqFjq7Ekq8guFXm8hfWxh6eZOSX+NMzAGS1pimrzbE1Hi7LEneKy+yuvJa8e
9AfNBrR/8HUfxNTwonPteGfte9KHBkTSnNJLGiAqEOeKXDDLH+UnAHjHBHmZZpzf2+Nyo8AQ5deN
lp8e+ATXC4S6H8358t0oNMLcT8OI+8BkiNWo0Nb9XS5jjzzVhZ1OFZfjW7pvNti5F05PWNyd0FuO
geiXpJX1Msc+hagdqoKsbsrNB9psaCGCM3DyoUWx2F9tmO724MSAF4pMd80g0jRHg5SCA4p22uj6
Wc7bcFDguiOCk9KbeQ5e2TthHnUwXC5d9Oc7RTLFWC43CMFvIPRbQyPwz/+l5Adsde/dK9kq8vzK
8siQGeZBBwLOuVHx8xBvdQxGAWkvUS41PdXf3NYpp0/cDp5Y1Wvb/q2yI4V/xJjyZLDDbVR5r9RQ
N0sCxPnoWVnZhHOMaQr1YIRcKrfsNziPhuIzFEDDo28WKNSJFtG3X+MVDOZIdUegsgdr4swMIIkM
MEG6x/ZXm+NThBCzTDScMmijk+gJb/bSkh80g+QVwSKSLMBbs+t33hlB6bjuY4hTYv2hMkPBqh1Y
EMDT6LnrRHrTBlwUFeVd+g+w1Q7kE400kh8FqOCx7Wkd4iMSGqVhcEPf6MARYHPZPpsCwn5SM5sV
cASgxnJLUp/6RKGlhkOGnkUmWuVbDk2gBUQLwJsorbVpGQwiZHG1AozTTSseMEHpM3SAtq7bg5nY
c56pOBViK924ohL18ayNzfwfZYx25JgeSF6wP1Vw8eQw1IliuuH8+4MLMU00l5ovQUKL98yI5Dei
aNN052TZBV1AHpU9qsRv20JfXzdVvDd7mEPV9hKCbyHhxNCDMpT3EhdHBwQIJ6X41LrezkVDzhKO
IxPWFo/BUydpuEBUzj3/5b4YlXcS+mkST6cEL2M1NzxoisfnZbJ1L5pse24cVkA4ip7o5ZCZZ8z6
mHpbo+Oncd/SDE+JOSeRhVSVC3d45ppRBkp+djtqRSKg3QpNY3MtVz1f5ySlnqoo/z87pzap5PDY
z2q0mgJkLAoYyV44Zf6w82tuifEUmdnaXybaTqaATXmWmCqSb4I7mjsc3ozgSoKDKRY65xPXPyNA
G+6Y6dXRJ250fT1I6dNK4P5JfKXS9oSupVk7OsPJheutVq/+3JIrcWolTe435aK4AJnKmZKhHmOh
BcyJs0c9zsAOGdrFp2CtTBBBWC7ndKTsv5D3v9AL3gG+NkvzAMKgTR7TYpSLEm4vzrM10J2OZNHm
D3sjc1pvQfQzjb+VwYr2rnSnN3g9fSKzTIVLDkT5kaTJ0PlQqn6dp4VlbtFxKDixmhh6ktd1lk1G
TpJmDsOPaunrL/pUgOa+NFk0BJ6HVu+BVwrSET7ynjXpwgz1sqQORP0nbqOa/HH5C+sxhPAt5uxe
IxNehc5c6+MNT9kDQ6SKKE7evXXI4ihHXFbyx038HVIA+CaoDlStyKwKNfetA34FjWMpqIcVx3gu
+IAfcrs88293vWsdDQp8QgPSyh0RVE8Jr1jo2DXeDJfm5O17RC7F3U9HyL9ygJn5ZgaB+ftx0Ic9
aMSp60jqTRXaprZZ33eJVwXnWBlBfbFHKgK5szt33nSn9dISXheZDpHKuc7ys1aFvHgMzL+nxPp3
7cT/76Zz1fhRbO1jPy3xe073rsGSzIgKGaTLSlqnwoSFTk8ZfaE2/bsGRmAGQjmzRVkHpNMAj5pK
ETfwkcZIuH/1qJYpxtdVnlXR2qDceIuUc3dc+I8mH8QkZKS6BIeiqWUDN9nGLg2Zw/BZWnWMjpeC
0FqhisSWBDLjKsWUIGjUsBhEP3MRcn6uvpn2wjE4q49h+b+L/lG4QKFy5tYW1Pkm0cqyQdBKOhDQ
RqFUtPUyqUAtjqO2BorfLw+sA8cUGspT1y1YGCc2pifWvDJbXx+Klvwy96xIHh+wW+44uc0ZpezH
pMLSAuyVJ9slNVpa38LMh3spgx8FZ3/Ol7sS/d46+e9sCDnz++6YpggM/tcd+4zMJICL4Df+JkWJ
uKFDFD+Ku6p6ZSFM0ccCxYsQ5B0fwYYu+TYIFvczgXD9IriXAnChD1OHk9YzD5BdbHYRrVTe4V0v
07vt/D+Jrm8VS/lypcToFUsdjH/RtKwANiuRu6uwfybpdp1qqSnPx/6lBp69d9WTXp5ThYdGNla/
5wtky2o/eiUSQvZaWFlkzI84TZSeQMYfgrXUvJ2C4y8SO7TCAMC51FpP/tsbpZ6vyD6sgqtmmOp7
b4bNMUvxRh1Op1adBlsv2vGkq9LhLlzn048OIEAh1BP3ulGGW9Z5FtOb2zAvcQuoJ3bULUyFDfan
qaMz+w55C+M4s3SCQqrFVe/L8uQiaYT7b7IZJ7M66JPP9PSESZE7Fr6GBSVMr6Zr5kHfpJM8FhwO
gks4YmKLx9ZH1NdAXlSFRvWv4oBfmZj4DcPRd4m+tECoCjFoPXC5YmHV914V7oCFDrvRfkNfc1Gv
f8B3NJUkJNx+DNvLGWVnbYM021cK5r8MTJ4xV5qaF0QHd+KXd/ok6Jx0bKjMLGyF+zdC4upy5Yqa
S4QNODN0DErBluoQS558kFAPPn15hkU9Ih6uJ0kN4J8LioBBTplSekwFh7stNaRtSrE21BwqJD0u
6ZWYQH1wacU0w5lNAy/ijWdgdkgxVmAHyczkK7KPBcsWa5Fd9LN2O2J/YEn0AjsdcBmdjI36RrmH
9KsECdTYgQ8taHl1HLD0Sp9hhZE7TUYbSK9g/qqeO4vohcSn2Y99s7Gv/BgIKfEDP8P5cMAPMS6B
rQ41CsUr2XJwGU76cS5XsEqFoNfJ7ddepRfXkYFJio/4bls1mmpt4krQB6FDwStW1n6+oAWW5h+B
rQHN2VA/QjdB9PVbRO5lCpIyBRae751b2E5k1mLMHTKjhnmUFE3vTNznTzSXaiq06Czh5moDsfe1
OAacFFS6LxV9ChpC+0HahVXvlaAoMcjfpbmH81FYyt5lNs6sGxU/PAxaJEcJ+u4dXuYZ+LqV4gxC
4HOqUXUSCdFmnf4zhVdzwDABciWKpeeedqicOK1OGNk8yJF4fkxEpCpG7779C3IFVmQno77t7r2s
nKSVac7uxKpFrHrKQ+3F/Lti2+YaZcHveiiAMYANcUu9myuvKXZarpmdq8Y+VZLvWSfSUhZpUO4h
wQB3/bPch/qcqV48Y4wanfVODmVp2I7ZclLEY2shZvxGw5XhojgouPo4jlff6bqgwaZ7O0UMCkFS
Xk/TJ0Nzuze2e4Vp72ZowszKtCx2dvpTV9oWEbpBefNnr2NYN8kZ1484k8xBYx9k1+efKEuxSbDL
t8DyAZi2rwAlmITx1oM5dfHJLg8yR5ZTz7GExNfM5pxFd9O9M8h2CALtdDFBNUvkYCjna2C6llY3
aY95FL2QS5nhDhb94E2bh1xjYsexZ/AS0f4GZiX6O4ZPKbg89eGxM124QjdTHxRd69EwQ3dT2Kji
QAMZuyTcFKOaz5cL/XQV9251ZrnH7CV1S07ws+csL3fFNFKT+p+gtN/dE8MfRot0cB+g2a2ui2Zo
MVXYZLNrvoZl4ko2W1F6nPVluLtyPajxiix8Ke5E+eyk+o6AViklU/C+C5m0ATaymphSvneU6bB0
9kGcQYXw5X7PosA2ycKTN/hPZQkeWGPZ2TEV/VGa38ZBxRqIN62kGCi2bbMZ2R/n24TPc+i/Q+ya
XNs7/8BZgn5EvEKgrtVsjR7ZtFkS4r0OnqlU9a8+VWnj90VxQ5ve3b6PydtGlhKBLm1u5MaHUO45
ylE+V1MboumonLSPubA7x2AybtRecnOIxSWrxio7RhCYo2n27+ughkVoz7rPzon/n1Xn93Latz2A
TNFTEVGxaLAazzdsydmud3mNvuSo+ZXawqTpKdfHCnNLbg9DhYAyCVbTvCba96I29oH1roDbfe4g
9u0AOkO3lGPdtchFv37xLvg+QRrwf6AwFNxb4fe2feLlvJ5VU9FMNQxDG9n8KfULMzROvu0kTj7L
EadFQiBx0kyWOXq5K0i37I0nLMghWRHw45NcKcO6SF7UOYhPV9BP51hayFrxgY9mONuhV/MdxgDt
JxMJVcKhC0+MPCcNHpv1ShoHvIGIseVaVOI2lto8sc0IBBnvySPnNt2sy9ta2F36HfsBankhsC7q
z6jC4q8IRzfLEz6Y23aTkmJvmW7xbKnzb0Z1LJORYYUneTmt1lYPG9N27LUwaogbJmCt2ZRw+OrB
0JWlIVJq2IYJhnVXfxXMSxVUz4ITEIpC9lqattOCyaLCJUx6sCywySjvVlkj1uD7vhUp7R2hGWuZ
46iq0ix//kS85WmWZU95RYxztCwFWYBVcSZpRB/GJ7hCsdd7YyM4nw89172miwcRdVG9C7f+KerS
pF7rdtpXqXJJXPjMk/HCHq3ukiM39wv8ZF1g8FYnrclhNfRKb0erSmvwBJSMhgOLK/iId2LImADV
pkdpmP1GaCAComxN1UcYUmZXYWFiIzHfVNI4YWYAHpuVaOPB7pdNiOEFqdO/WBdaKh65UcxLdGKP
sehD9B1sFiQvC1QG+e9TnIMCmh0658/IWADNpl4tok1Xu8DFTb8WNrVB08EU6gcvKLNkbJOuurd5
Qi0Em9WcRTx7U241Jo45PFLcIyIC87HT1IlmqIXSvM86/MjB6vNqq/OBNunb5+0Wk9VEIeL5SzFB
NP3dvY7ElPvkdCoTvM/7WHhC7cMp15eH8qWni9jzHOoi/GyE7qApOSMu4nxWXfIovrohkqjYcuU4
x5Iav5RcadkPtbC8BAndkNv7oi20bWw3SmQhZ7RrqiKvj4R46UJBtm5V05wQQeUcblUWKK6NNTmg
WpMZVHjxuNmjhPMJS1K9mk2/xlUH/66bZgBdY+ED6klXSLzOC4j1GZZDXa9Wkq2kLxqJ/SvlA9kn
AiKRL+WwFACXset7XNCcCpOgtyN4WjICiqMPJlorJ8+MM3qTD96eF0pGMdM61sKAXMtqIwCfeABu
Zys3HahmdqYW8D80iOHmO5n4EWdjFnlgmdgr6J6H2cuc9iJzIVX/MadcF7+i9CtAWtgPbRH9MrAm
km3NzjAGasecDRul6Sd6zbDIy943RUb1yHY5tvcMM/muUqCPjvHVLzTRVh5J3Zqt+RLNYtMs2Ex5
a86EQFsH6LllQJh7AO9t0qdptvfqNfJdkrsej5lKgQpfuD339KAv0p3AbY4CtlnDdSu+GM5Bmpz4
LccCvPuMcZ+nf4jTcfvPaPfpNKWwgplY9/6ZTWFN1P+eUricDBG9r2BapSzgoeNaeZVjjjXX9Z3d
JdBZkk5/wykK9Ho4T3y7YqDpMlxt0uSiwb3xpNF/pdDyY+UKhgI8Vp951eeEyVc2bwEJnaeK9Bi2
CpC1Tsc7+5zD1rdsJCJh+7AodN7svjKu3Z8NP4rxyoSxh1QTxsMalliOLpN0nCAZQ1N0j0szhx2P
5IQqw7imzE0TeaXwYf/T21yncKW5i8zCi2c9ri2BXDlp7Fd7YPGEa0NcVzjQC7byKr14Y9EUvpp5
Y7cIm6hAI5+YZCDb2sESeldKvoAlgZR330rudN9VbnDOuC1XmIFdVhOpHDnP8g/KuEf46zJO5YAX
nMmgjItkQB2Q/6Y3qm/CW4QctpiYfA1dJD15+E1ty/1SePyxUQl5cNnx89D8gcKLbR2mtyHf/d2T
jJAH3bIv2MQ1GOMF24IJ9V/5qsbJBR61HmNzOTg0u+HhSq9o+LR+rsbxsL+dtxZEQe6+b4W9801B
DOlW+PkXZg4WeSMesPfHR+ejTC4MndmiWMIhSWyEv5m+KyX8zl3ZPPtWRCXmL3zHnGTS5EkGiEZ3
izzW/UkC4f/WvQii7CYNqe921v4R8/Nw/R5rbldzDHMoUz6kxcEbHrXqZzJ6RmGy7du+JNQR3Tc0
f1gE4fbT90JMoFx+WrX3ki6ecnuTkS/sYUQ8+f+fw8bo7InyfR8yAWkEmBnCk5a5lIay+gSyj592
dD6dxJQ4TfEqNdoKGKP2fwGJb5z/h8n15YuCUe1UFrLMC4GYtdgQMwpGihUJn0qwqxzGI0X/v8df
5XhcBHt9ixAnza95vEpX01TppnG/OgZSHQXoT7BPfGqpOec3BsAq9Bd0newO/osXDgZJ5mTFyIZn
Djr0Ml0FQMakooWZ0XquIjn1bz1EOjRY5ljrJLQGKzjQ84xBKWKvHMkcDaweZZsCmsK/0KoYCJFH
EOR/8/FeSyTL/KA4zp2DiHhefl06mDvLryARzle3j90EM/LLtRgYMtbBPZ4KJLOCz2XKyJ7X8I0i
FwDlceBnKZs2gmCNYORQbA+KdkPMIQOdQlgmLrOWdDlxxHjkQnxxDKafzbxxa2CnE90Q4ju3i7Cu
QcOZ9UuEXeQ/Fr3nqEJ0QmA4ESiYw8ujev3Mh+tCG45lyvnhJhQaHZoNDCnJ9EUpsRdYJPVqTmPW
C0+veQDpDwrHR5+Fbc9m2D3oLbRmoJkBv48ZOLIqpR5J2zX3KtA/SSKEL+QXzm/GXzWcs0h8mEUo
5nvN7TQrSpNed+zCVmQHeQuuM5sDreR25nce6GZE1GN7dVKsS87CAv/FJm0qKI2w+WDqdNSnhsrD
pWe2ti+K6y0wH35cVn54MQ3Vb8qfNmrUQH7i/tZsZd9QY7mzp9KPznX2Hvqerku4sM2dYkWpiDiQ
yXSZVRJsxCJGjh9vEfs9srXKOGdDl0SYRLWh9C6N4KQ/Nz9ykxCeFfk+wIn6a8IykmimoYXC0ue2
R1nn1j5PEA8QybPRKE1kUQ2Hv0SJDNq4DM5/aFx5xQTKSXaPr1OiJXtN+3+Ve9E2HQrHrYKN/iGl
DgbQjctK89IZI8hWVEW6zc8VySrrEChQ0McAn3yq/O+aEum6BpHCVR53VQssaHz6gAd2HZuvKlEk
HIpoMptFZac7PPfLjy3geWuB56dPTKmd9vZdH6jB1M79XSBlvBLb/g3Gue/G4cVX9NCfo6+PlT5I
KxA6yrylL+uvDh2fH5adWYK/S2Ow6OikaUzGWoaqFRq51fUILrd3Gdj7hBMC75XJs2nci46K3cHz
VR+JuEEQA7OfuyAxAbF5+pv7D8exis2bj86bmtS2nraaa2+MGGvp0qZdMdGxcactF0plc7iyxWWC
h4yQnKNL/jbmwkb0qi75PU9wTc6zoXQBGuw/rWBgg/BSbIdH+1uLND7z5kJJv7qZQ1EO5CK1MAqB
3hUdJsrBSVM45HssZeH9Yq9l6rwQsAMM5VHf4nGhXzSDSci6zxZrJdg5U/T0lSd7SZYzD8ijOKt0
LMNEX+TwGoGkDUulJ7vRBPwK6SRErqhfEWWgIlZvTsDZmz7Dc7+6PnqnO+Jo+CXwC6tmdj2TKG9o
tYNFcWuMKQmlyhZuIW1L8YVBnWCJHrpY6CKVH+KgisxlroAFJcIRxdFvD48uZ3SUTjBfeizOnmYu
jtSaGQIAZx1bj42TbbWXlS45RfbQCuT0P5M6PCwyQ5uNr+93jPIplZnOvDr1HCbRhJ6ffURe0F5c
gKkDzZNhpcjz9uQ9bDx9xS4D7b1z1I/TP/V7kDZOhMZlDOfFSaKo0Ie6vGfiEWe40iVDBftiZYKI
fxKjdueaGtcpZeBg3+UDVFwTL+NvtfImwLwyG3O1hPre6vxb6IksFJVzAVzc4hQ74vnsIvnDupvt
L6aRoOcES5fZ9bVZoycvkkUJ4jx2y38la06FSG359E+sf5uvBzHLN2NuicawQb+pl+W386OLBlRZ
MSTyvjaxEPDEBAkQzBdquOGKLeRnfamuBBpY1vUTMBcFhm85B27PiPga17XsVIAr9/Ej5SfjJsgu
U+Frl9vBsL7vwA3ZTvJ2Q/I+cXwiVhZodCpg4zGYXr/3G5P5p6mRzxrzUYkT8l7X7wBIZtKWIj4H
Mzl1hhbZ9x1dsr5hwIsyeoV34bZOBe+UBH9GO/wdEt5ZCQKhT0I7ltliT564U9odTRGdtghyzIRL
LX69hQ6x+soQ/F5WdUfbCb5/ZvH/z14gc4msINqRiHpfr/S6ikziJNIzFKvPCfhtjIal5iFLLMw/
dVe7+H7uJHEkdI7hR38Urkb2ORLEx3rOkPnf9WWRAgj3cMLLVX5+9bamE/RPlOmfV1APUrgoINRy
+MWtMqEJCCGuzUO/ty0RMcl74rejPf2/seyEqDo3sRSjmI6b4D5JKRJ6rrp6TeE1JYSMeDSIY0aC
oC69kQzQ7quEcskNGEDHWsi8ay6AMM8W78R6cayGiex+qQh0C5gS4Wzz23cpw/BXdaRR/mQfFcN2
mi3U4sbf8PoJMv0To9xwB1P+WLtkL95AcLAU7jlPUnFdOnypuOYC/Y1/bwMrYJahJ2px0D4cq/h9
kklMIaIu043kRxsSn+T9C7fK5iyhcwo7A4GjFJY0VHvrY/gy7s77mCTcpf38WsZDlEyWVkfW680c
0uyEoQqH3H5hr5amdy00hWQyPDvSSxgOSQ4ugF1dFck+Z11mMqcfamMLd8m0lC1X2u5yOTAsqOpd
ZJuDaNv/vHiGQG63Ct1CT6HdskVVhG610uKEiZujv0aM4axW6BzhG0/kHChHQrZbNB07DntltYRN
hWbfCfSXaBx9xi+Of6c5oAL+GD6xMQuD52AcFloadGcAtgDQ3n6d9IcHKnelM0dpT2eigSPU/kAx
JVDMzP0OWEAsVi+Ds8dayVHgwW8uwlmvTXSLsX7LTSlR8bczjjBOOgD2u7VbjCcwYEbe3bNFslBb
cBu0w6RLLlfd4/u0KLgGWPAuTDqb1yBkrGLvjsMRmk8WnWcXFusvkCsdUrupyyyMrZ2Iwhg0sFRa
Fuh7jTvBMILxIvNegRluO6BG6PwbdTRvqy9VKDHbyuE3nbnAtWqBF5fh2UQueNnnMwVowfuk0mAr
CF6dsuLmn6UFSdU5+0oySdiA/AAsA2oQGtlhUpHSvFDhQ99xxENCSldz3qwOc9aIFfZ41zpSXBlK
qNZ070UC7abK9IJYTXfEeBYmJn7fFbwDNEQshulljqGBeBKVhq989ga0abI1SwbtZKej1KyVk0KF
CF5ji1QVpbED//C8kuf7rcuwds8n5j7TzB83FrfYFmD49f5JLoFa/BB4D36g/VohO36CgOK8V000
jaawauYzDjIeuXX5U10LimtexXHUKD2HnBapefLM9v34Iskt0OXphtxXhAcNlBlbPV+QT06FZ4JN
H6SYwu3ErzyqGPi2+3J0TrjFooiA9NHW/+q1Urd0gp/lhSDf6xgmKHANkY3HT5YutFev1oSpUBC3
v/ZwQoAujulyWEJyPoZ0BzWLLRNmA2QXhZwqT01ke2JTbt5O8iEexnvgpdqbLbyrpZlGDEPGzasn
OMr8DRyUYqEDxXYefw+j4ugOwktcgIy+TnkEv1ObOn8hj0BQrDmauFLyhYJf2BQ6OTPxUDDDdEdt
vPgNGFN8dV7lOT+8AWRm0lMGptoKksABX/uzqm3Ftx2dOdOFScf7Woyl03dhPjYnWVAK5ymysq3f
7LAeHY9KVneor+XKmECwU9C8kouCNcD6fQ5ecfyr8pAJqHPVkK0pK34GLMquri7QfYz8WGWJ4iIE
gml/PWy/DhekOaCM2EMWCt991h8l3k/PRYRjSglSNQscI+EOHa9EyHDeMFILSuY8kuCCikRa3zh+
WGGCJD0EErUQf0lNr9udMdJ8t9FKq3V9ampRNFS7j691FtElwfPCNaVe4cMk55Z4VUFXONIg5S6K
NQNQUfb7SlwRD7WS9rifz5SISrf4ye49/Uz42D6qWa42US8ef4HCM9cqJtY5dAe1jrcIrCFfkRwP
L1fnv2BV7n5gCavdXw+g9k7pfoYDFIuV0uVKKZVr5+vfdwcShPYnhm2uKZQ+XMcd8+kGHv0taCpC
LPPGE/irVb8twROYjtDmBntseSJl2UVQwbUaf0t9z5gIb4OQIt+2y4icv5cQ8P2Vb62EZ02wOn+F
tvN2W8Kws0vagJYJbYu5Gp6DCMPrOEaT0y+mq1oBd378N4ge1aHxEZUXfyDqKhktdZ9mtImsHVVh
ZPSDvRzaWJixxSfK3N3LI9ZZOqiW84LGJP4BVXmbI/Yr1OC7KJONvLSvBm91Xs2nmfhsnmt29NHO
Fp64YokQADZMVgRo1gN3XIiubbq6TdQXGpN/uhTPtcAsSxXS6gnZ55qn/p5UN+fXh2nxPlPxZQJD
FXPtiMYoxXj5AwguGCsIl66YOuzzPgvBAyo8QSpQZCehjk3q36CQ4poofEFx3GbD3CBCRmlzks+f
3Bh/ldRcs0XF51RQpeexPKOcAXzX/vJXI9m+6LHODKY2JCmd91l6kP9Rl7Fyoizh1BrFD+GMcgs/
LlhUqztdt+ToKy1pYkZeCWzW+C0wP25S++ci91+MSJaoRPDDv3hqnltN6ttYSJuQecVVQmv5jWGh
XxSbjNg969XfvpqUF9MHWgLZRAwrMKPTyBFPrrljLksimrFuqBIR75mZN2VXqE0lmEU9U284azvO
c760DUI607J5EVgwuffNVZjHFz9zBIdGAaAZ7WnUP8rdMMRriymPAedNlmu0ohUGBenYk9q9BBv4
cv75ujI4DrE2poqBQ51i/2gKbYNnu+o3HXqqwgnp+h2cVLk/6izTsQtEK4vDn0juvBqlcintW0eA
f6FDOlY6r+2QxY64n+q+r3Z+jNA2nNDBuJYCr05smfzSPZ0iVfDeXyli/0ywNVO0VPpDWSCYMBfd
sHdAlhSjc0P31hwJMi5PiKYsy196b5oZzW0KceUJ5tiRWSFNbeu8Dmtp0qFxqHIyNaHXPbvuKVWv
xLstofuTt3Asj0D2UEA3EsifYlgmsQ6UdRkhVWvtn/pUqyTV4AvV4f8O+Ln0yHOLywrnaRDZh8Jj
2dbZnuEtz/1oML1oGrxisedabR28xxp1pP7oXmvk1iosCyBfjVZOaJhXHfJTNKxeLTuL42KvK3HG
flZfr7TZ6uMUy3t5DF6/n/hvnc7mmwQ0zW6d2kWk/QNXt5Zcu0tg4CDkrG2SEIyXlUxUwRPfAo8p
gQMmBFCnhsMyn74B099lzH0LSi1dsMWwYdJ8mqELhzl3ANeBNMLmDizD6kP4OXKyLE4bUdEtGVIW
XaUjzyalWMGphkBQhM+3jtp/tFc4C0klPCn2ADFzjeAb3sBTA9MVdrQPDvoSi9Rn4nLlQmttEuEz
IePjRQndfT8Kgbfera++AikKd42W5SPB7NLPGIl945q+Lw11qBxBO9VhTqVgpeJm4ZZCOSX4LETS
Am/fFS9m0k7Oz1emwGUd3MQ7Ubf4IZH8N/g7bys6NsetU8aEnCctmsIWXioV6e073r9Snpw/wtZ2
0cBsBHhiur2cG2NM3pzN9xEXPurGGhEQUrwdeq6JgPm1MvAEQpH4gra56Hy+ITJTsvPLfaU4GdNc
P8KhU0wMkx78+DvnT1fIUcoDau5my/AyKlgUHV694eOa7jD+WEYp+FTwAiWbesX4BR0KdiFxF890
uG2NfVanV3D0w4tjj8yXSKUqHkIfmyiQ/nsiJgq+4ucDaZRLhQK+WSY4Ajiya0etrNufBzF2jZL1
zrrUibmbZQsYRKbzLRziPWIsZaH5gRn+psgMfg4hWFRc5VOxM4gevnxVVEjTCixGZ80+O2Qbfah6
R7NMJvreapRbt68Y2eXNfOf9ydtx+md1+H96UFBDT56crTSdnRsrzxqrRaChM00ArX37l3VWeYJ+
eofNhYjBuLSx3XnUMMFjOpSz8y2npj8+Z4sRu+daozOjBGG9bORbujvJQENKqawTKqX/X3vojMR9
f3jU6KezNfqzPO43oCbSPa0Aak2ninmUMzZdxwJ7S2k59t2cQdNj/s/XR6ZjvVCsnZS20EXoC15x
t5mwp3F+cNowc0Roc7L5o9g8rtpsMZ1cQasX22xSE16VBMbAmGSKR3fQWZoddtSfqWUnwVSLvrE/
TWu8Bog93mbeCNbUwcWpQmFKveUMEA75FuqocrD/9US2id3xRduZ9/WHJOUp9W5FmsJmwhQndJzC
6xT9du2Y30O2fDUd1hMjxd3LaOqqELgEItYZ6DPjUuvKKqL6Z8pg5iAiUUH7w9G99Z7bj5mYDUEu
Z2gNgx20oGIZLzwR4eMNqEsFgOP29cz8fdvBWSb+mYaQff0NIWtKjxYJF7JcsYeFPMyVU8JtlIBh
gIW3bkjqio8hVtLFvEXazwSUqtZ5VXPInpDPAwPMa9UaOFWVWyU8htqJRqZJm0TNVH845KYU1mPX
J3VAt7vJUT2dV8cNCCgEyTXhuDNzYPOA1hhpNWz+WHpkLNTkQBZyejEkR109gtGmvF0jRPREfNYs
efzzJZyFEE9WMqEZTGcAM2bz5fskiFo8xnnzXC2FdNVGz9FOQSEyIeZXx5UMp/Fsw+8geVnjByGT
QIeqPpcXDgtB9sY2WKbRc5Tc+mr8zwpxIXdtRfgJQ9fOYUUDVpd5UULaTFZWCvnG/2DeXj0zIpjk
Oy80JDYbg63l96EZm4Ris1LT+QJ2EbWXLsscnJnFsFGmYkFa72TeR/WxpNKErsNZ9W5POyFjD/cC
xH2ppd2PfgocmTPSUOxdK6atrwYvr5o9MhJHeMqQH+bxQcr5gygGl4O89zKvoY75V3/rPcYjwsCy
UE1oO+yyJpS90EBUGixkEC2j2nY/m+G7Z+0I6aww1uXEt0Hifak6KOXgVJ2SK6iLC67zsNtZqMNm
WCQsg40P4KEZgeejC/td8dRgIepWDnVPEI8KuWHzbZRpBFXxrlczjazi+lK6ErDrmTBMxtv3Ldp1
2L+vl4yN7RkF4TeIccz0st2O8btdNqgDU42tog89r44DVDukznuyAY/gsrssXbyf5jLNcNBj0aIX
JQRhqclmfuJAy5QTHN/ADpgobGrTwBb6SXM8pjq3ntqe7t0DR+QT6lgy7zgkPuP+BE6ugbFO3XC9
p//+7KPVJ3QAjAR37BxsVJM1jHZy387i8uLmCgOsNzbO9cfypDV388YJH0uQbeIJQ1QdYth94pTK
MStaZE2vvY+SQEPbBpILt305S+uzkFqMWdD+PVjgsP/fo3sYlMjRVoACrNgIMuxON6ePszfg0GRM
LjQICiSJ5ndv9lSDHSZjuqe9yrhW9QKRijpsh4DBzwBTqpy4eiB0oGdY6bAsmDzMHpQpgNZHAPoQ
jTTIs/nn1ZxSHaMPGMUwnWm74aFG9rjkup7iemUkjTQt+lR+mj+aep8k9SA5ugEpwXntqFsppOHv
bRqoeACwYDEw0XKxe99pqeBORribqiqjOjPkUBQ+hnxfNfnPrturhJgJB+r1oa44Hm50dm/JLZ4p
AZtoXNbGMT2NYko/e0SLakmqpG+Lwop6vVX/4T2xeLozFOdrORwoPIU3DTnQn+J8LIHl5gxWfscD
qV/MYL7V/rQbq3Oa7qka+aaYdIBEm+eYSNYLf6CZkf1wSNpLgJzvyHV1Affm26Njp6XJPPjElDJ5
D5GEWVr0kx5mHLgSzfF6AHBoNHM5fdbJIH6eDykWP6STDvZkF2yFj2fAdi0sX90isQiTNZKTjGOk
z/cZy8h3fcmen8+yCNGGjlQEkhI2NK/ZO/KrYYVCkHlOAz1LEpPMSNXoDRJTysP9vUJ8dC43ohJC
fwFoNlkulEZ3jZCLzXGpalPcji/c+18MWlN60JGH4HqWWe1v8fwgBGAYlwbFM5+LCCIEELLuup0+
2vRWtDl3siaGluO/wPD4xfmhn955YDpN4xavyEQOi9WkgME3iVlSHPMAOYtVJt5VBvFy6d/b3WrE
WVYdEyIUeNnZLGMR2PJOsuHerJInE007oN0jMDqXC/4CbT6L3irzuDnPmw5UOTJAG0CFWJA8K7w7
35GWpV0pk9b7w0NbSGOVH4AF0Z8sIUSgfCh92yf2tRAe9KWRPb/H4+pQH+Dy66JgHluX7GXl+c6O
8WlE7NDEjOYvM12DekEjEVCESWpZnhK6InTOv7ffpZHTFgIooGiLzl9RxwdQKak6XjC8cD+WZmG/
kdSy64eEkicnRjmSE6rBYVNSHXktv9EEorDJbhWTzNe5i1z0hSmQAv3H2UpsHqnwts3rhM+p4AyA
mcfrEEG4L/wEBDMF3qXEHnN3h4oxEOCfYVVw5nsuqbvjMEKXmpKhzZDkM++85ojQScVM4cSXcFr1
DZDTl9uAsJBh3icohPGocVYG4zVBA3gzha+WNYIetbBiiJN+Pn+/bNnO6Q8cO4pTZSp28tfFFK5D
B2Jxga83sWBz6SWPjS4ib5cFrJ+rsO5cUhykrgiKVIf/fn86NzbERTcLoql2jvU4wXTN999OLAa+
+PtMcFO9CQrR7ZCCccFddCF0j9dARiOXc0JDLpo8700qc6U7whpyOpeOey90vUJR0aqibCvGEemq
VaVYXZB/fgf259KNJp51jvndOAi0g2qoVDK06DMKDpO8s3MroSa0w+xTfN644Ib3iA3LWW2Us/cm
923UZZMooshLWhg3wp16uXxly5kiPpwiABFxmiIZCIjwKbIioROdps77UzZ/x+9l1tVoq3r44qNZ
noi/LMc2tQya7F86pO906nFKra6KBNnjL9lE35bn46Xc95SF17EHjiwXJGO5Pw1H6TyEl3OUr9Ub
TrFs0bV2C4sQLjpLNA+nXg5rEV8yzgMrgcnwol7gdBh+KxSaxcmO+frdTxfdUtiqVwwwEgFrDxlw
YarmE4wiu2IGshWB1KgxOoTd+ZbNJjoWujB3H0Tcl2UsC70MSmYNE8r5CfHEinQtkcbnjztVHS8g
9DYiZofdRRqLp2aYhnD8MurvY+iVgk30mCH2KKcPambfJr9hkSZHnbi5xlqJNBt0TMXCHTJTa2ri
sm5C96U/jexaXkMsHxlMfQ+8HCZRWsHWx+1NQL2PqbYt8ULi0lus8qVeDoz5+FzGt1SA07uMDcjd
R1f7DrWuwzFuuH3Ob3waVfhllC2mQLtFz96QWm/V6eyP83cwdJu2dWjRwf3IQAdg7KnuYgClbfuw
lKeirJm8ZM0MYQDLEJGNf9ka1Naims2PEe1/X7ZG4SYPvI/GpIBOOqSX+CJk2LHCajiAUm87rr28
2sfO7O+1Fch6PfgyJSe46oI59LJPBF/h9T5cagVWu/YZU1O3y5NdFWhgJT3boHgJM28hAhxVAzfa
6Q6Dvak/yuHaPkiYDoGc5EnYrdQdUMMQSfEqKZx0+mxKs9OiVkEy+Y9SUaG8x5gT2+JQgFi4KA8l
VA7ZsbKgyVq1n4n4Ujz1KJkF8xAgfs+yOsiYFFwgNdQTaja3XLQKW0jhXR9LdfJdMfcYjtvKsLKc
NCLbmr8071cU17PLD1d1e2oMVsOtyLEygwdCpAIGgewEkWMUVa2Af79HueDjmhGOvm9gtvLHCd9A
7diBcRI8HIW+ilMGmNx/rnjc5r013ebRUIDOmNJgf328AIZGs2LKlrF4zIdn52sl16BPUvIFtthk
FnvdHLloco4C1tEA8RvwNpyPH9bo3EXZGaOIgl/jAi2hp4CuUajiFisdvztcVQqtqYDHhCO0QNfp
gxdgZAGqZPUB6iA/OX4+2NyqXGhnj9vpFhEQmR08yCR/f43Xx0hkfqsF0rNW3LvnBNsRYKmSZzd8
SJuUpDuOjUiXpiQv8tAXPttEzf3fm0bUsG9tNm6E3UidkaogHuVjDfoNI9DtCWymntDNxxcmv9sD
qKmBVql8cv+6bPO+vZCaWyjua+DduvHZtqiTnwALBKiBt1c8RZwpZpSvo1im7ZgI7/hpnl1/aRWr
ALQUwjQYivn2uAcfmJk4KsGKr97d0ECflMAIYpGXbhPNFFyNxY0I7mIZoo9X5a5cxydUDQFcTBib
e9ib5hm2Zg0sNxG5D5xDVx4jeAl69fWp22pj/OePiIlqD8ubIsKlH0KG+pqgLr8eMtlucCmwWb+C
eYrxKpf6e81eQ9ZR/ALaF2Pju8AwODpjR6kO0qFVh4ESzrFq+sT/+oJqlVLk1Uy7f/qYBKI7QpVD
h0NDCizb8fVNxwV9os+fGUM6kZqeWUaJn+NxGwY19B0wvWMhxGUb1M5AehkZ4tFfeeIUXdZ3eYbP
06AHu6AJrltOI5oNL2CUI4LcmycuN84V01hfbwDJI+rHuRxuP1Hj5hneTqCW571+hKo/yvF2UjAq
RibiKlHcp6IjxCb9NxXR+t4rE/kJ7j39Iba/czK1d5X+gQrc4NCLYGEgcBabLL5E3tX0o/tNwXha
wtW0rx3uAHOJb8bNTSlaTvUfo+aMArmRL13Ap+npMqv3CcmTJTlcnbH5PzF3gciKW5fFQS3PFo9R
sOygH/FtV7YkVpLOU/eUKLS2iEB6Qn1H3WMWG88L8hqynbJ0SlLRofXWGiUoQcqYOyopb8/Oo7xH
pk7yYgLbrNyW6IWnws4FKgznHy+PAtuaVng9kPtnr1UVAAHZQqsUIGpEJAdv0rHCNpKvYOqMJkMv
Kn/x1aFA4S1+YF44vNPhLm/n2NmdAhNaC6/NthCRKX+DLY1yqYpS80nbkHlttTGmOO/yHxzRLwP/
BIiDGQKSBX+alPCd/oRj+BY+kjE7ORZBnB3rm2T+JEjHapNQGwAYPD4sdHT+AS+JWsdA+D96WIGo
Uh3NcKUoDxhFUj0XdRjUBGhRdfbeSYTxzZ9eoKi6dYA+VxtEJJSftQEoCbaxsKUz7aQ4gcePwId6
vrOYLoB9WFv8sY3tX0m6NI1dw6H3K9g+H9DtDJg0u2Z89YEfxXTk7GelTnP+girfHtH9Cgj7Ouat
+KnR0QaLzHR7frhbPzdo8+a9ucGp1buv0DZHndWKbOqT1346LfW3XLkmmVrzCAT3U0Nk8EfKwJXT
r55loIAiUMR42t2aN1/gAmL/8PrGDf6esrlQvWbJiZC1biFHRuXbWVIWFZXFKsz0PY+CElZpiHv3
ofw0IcZMXb69cr4jXPTFQPjtrwK+oxWDfRfuc43BwCuSnt9t2KGvfyFDZIbvRUesnWhgQ6cUt1Q3
bdPn7NKBCnwhewBliISwBTPvK2dIVSOJSq5Pcxtb3r9GZTaatRyFPP+MgS4D/btuDq+WMuuXmijP
vcOwclFGtZ1P60nvvLG4JJB4zN779rWAvInCP7CYjopziYthv3QD0ACBjExUYzAuoQwj5yFGZskC
SBqplrO3upjVa4aDU7rXfpQebOxIG0Q42KA5vFd4Xne+YPeDcEoDCbnN8BdVq2UdO6JKqocguT5A
nnLY5+jy6aznOTITat8DfnCanenNP3dIJ+DA+1jQ9jgunVu4os3nuprl91II+AdN5+AZETOXAjyM
s4bGFiIjeAata8eb3QX+Qon+8B6b+sIM7cNMp6rRmvaZ7vz55jd1VRD+EQQazXhgz2QbJaJuvT/i
li0cJdNDKu7+9OZkiON0ilhkS00s2WatON9PetQlSfc0aI6RXEJkruXGhQ9vK+wixndyUw6RHOj2
0aXry7YySufa0cagbywX1O1Xd9HcqSU6Aeo+6GFq7Xeh8EhkcM/BjX4tEIADiwdUN0SeROd9qX2d
JUpRrL5y9kwpH9xa7vftugafNbs/k/73ZCGhv/68idvwbp69CbzN3vPxNhrJ04QpWnkOGjCYU0JO
rXEXwCvviZtH7+Q3OJrhIB5GyP+nvIp810/MurnFMGt50DNnhKsrdDCTSPg6XyTi3gieiwLaOoST
Wg5KWY4HvwTQNMM15ln9Dn/n2yRQk3gv7Jlpc/fYh/PL0EktnO3SnzCAI2kMvD8NWKIsBja8HI/d
0Q9vno1kF5oVGPRTlRqYhJ1libxT2LHPPnApf/81j5Hacemzi89atilR8vAXkK2wrdCKy33XAo+1
bcbHlh13ZDmyzAiquYdgplFgdFlZjFkjoD27Ni3I9G8aHv5GoNQncUwo/VSjBQTe7x6uN+XfJOF8
4Wz+YYim64Ybdl6EJEFjbfGbBpx4oGlCRY5B2hLkZJWLsYBBQDOI8tQ3S0uu/nOrZs7U6FjER9nf
KUD75Sv4xEppvJmv72hIHhMQhYhdtSgetGb1TplmkXPi5ZRvyYY0iz1HIIiSzcXmm6rUIpcZwENx
YfMS/sbWSxgNncqhHipFNpcAqTFFPrGgqekvUbEjtXOLQmpYH84kEc4F9bDIJxSUKowx2LNHlNA0
8sChuHjnnHXxl3UsagfBWUCLlsJhP0Dkzz37AGPiJQS/cHK1ynYGbzbGkNUHt+96izyUpAYfUYLG
ktym7z/QBgRuZu0RNT4xNeyc6JYvJ0dURH9xnJq9EOd+f91G8R9JrT4Azd9MV33dvApJNGFmeuLV
2K/w3zWMlh/yVSDNU/dU1p7Q3Md1ZBxG5WX4DiKCM3OvIyhTYCghwGc4BaF1G1+D8CGDpyYMc5RO
P8QVLV9O3f3CZ+ltOeZuLG1KwYISGWVkCcjX6Mr7zbD/+36JyYMW5eIBrkpdyDASviy+8ARJySBW
NXL6URJW7G8VMfqRRmMr/aEJaRsWaLaBsWeukBTC8JHrXdvgnL8PK/+yFpxkrU2bI0jTRH17UGKz
ol7rXNXOc9NgArMa7qxiw/OXav+kpEE5KbWxB7QRfzLbomqvJk1UAB4kj/uf6mnMGlUp9U21cgNx
V1M7SHQWY0BbuB/saw0EyCgCNxNNUnFq7Jx0n4+ILQotw2h12B0qAqhbwFXZhwgf8HJEHpEHAe5b
HbLKsNULEKiT7GwNaOmAZv3K5+g3lEkQC4q2GYoZNtlTEpEgTuwTvo43JgIJaBP90QTZB++b9ny1
NR2Og85iHAUUm5i5ZTqChOoA4DJQCNkU2XCDcKQs5ugiBxtDA1ahAHD6eDZnvqOf6jGCQT8dJbaI
40GgcNbVthVrYGGRTgzlTLkpomHYywcb0ZYuomU2BEeK/zMIpWAHJJxD+oGzGhCWf7OCpok2Vasl
rMR3UInUcYHyQgM+JMgzcDiqGzbzOpzOS5OvXpG59yoDTohjvqg3joUHEx1tmxPfnTpa6cYd5sab
D7DBRtQluYuvXusml8CnLSKi/50VAzVoKeLBu4IhNsNcQUJhJxzWz+pnvM+DuHeWBjVAj3/5kp82
kHwry8PSeFEvYm8VzH8fCSINBo/NS0Y5VaZGAmFHqFlic4N3bY45MDdXy8CRskpulk5/cCVGzUnB
tPH2J5PqHrYP/UiRfb6yRJI6gEWiVJ9AFKeX2FGgKdUJ0GXprBmqhbdgoIOMA5mrg6AXv6KIIIDD
4C9nf8qQH+fSXDkRk84jzXI/Acz4CuX/O9Hi983EBYbTllKhPQ+2j3K9GpinpKJYvq3e+M49nYkn
DuSLw9aDBf1GIbd/5Zn7MxCWOA+kCiW7oYXdCuIXfI5WBsd9sDzLDld9HMccLFuotW6pdWl31I/u
lvHLKoEAuZbfUJ28cPlJpdlEM6ONEcTaM086RF9yr2//jKiIQTTKhBVUueOUFiB4MAD9mGH3FG0g
M1txZMsVBRTWWuCr9jQCgx/e2cmdNDIfycGttzl7JUjMyHEy0a63h4hNFM6IagFjE6vzaGPURJS7
M/VV/VmHvT5/1o733qg1g/TNSeqvrmzzSIcDOBPw2kkaSvbf3mMhe6TLRALaTDJUYVdyuPSMyhcv
6k90MP1Cnm/k0wnNq9uuiKgmi3QeX6Vs3dxrcfN8AbcFrOOdlDPj4AjORWOyNf8BcTSHbTN7CfYh
DHaEAq1CqIlXD6Mvxk+jwGsgurNyZU4OZ1EPUbP7a4DncYT5hNa3aNclSVvLjEPm28UJGXu+ybHZ
W7ucAl72vUyUG7g6XOSv6jBz3wXbNCTjju9Q98DJ8ro7h6Jmyw86VyMTQGy8x5qLwsvTOzCtJwk6
OEJOBzd2lBzFJmkadqnhs0cTzoGVVxjKDDZ3SWVH+AD2wEdTHbSTfRsUjBwExonwKHEEGrr5LPHO
mL47YQAHOEsFRHbADLCaqBQJID7L83Tkl+8sB52rFxa9yrJ89hJ8UlWBlwPNa6z0JUyNmwioCt+F
tFTccEohegDGzeyTqdURyN44gcdD1lpvHCOtuBWkOtbNJmaaHbABrq9lRXxxz7LeO8TViHHRFg5V
Oj8oF6k9rLUAaqdmZWACPNsV3r3wYjbhBFLt7gmfZE7uq2FQIz75g7TNBouNtVqJTL4n82ZzhIml
Yvwp08FvhnGjOUJoeR4dUqpngKZBQzt6LDQaieS65rleHdbUfxqlxpDonQvN/RYbRTZOazniVXg1
YrxZ3GuIG1w8oCRwoDwltIObmCkAZkpaWzIdLX60aUc1XGX+Ogjt+XQdjwmEnQtd/YetCv8lXFRa
bABfuZbAdXClabtq/cqJ0YZFIzsiEtOi6TiwNZiWF3TMe8npnsmatKpiQvcS0M+IYhNv3qaqiLYs
3IwyklEYzfFaIZUQlbjklpuAHUGIyBqoBvWP0K1nea0yY341NSM6iT5kU7q+7qRnI8b5ZfW/xgdv
kljJqup94GGVNc0pOdGb8mS8XM4TfgSpPWmyxLS5kYh7ci3Q3VI+XN0n5JbqtHkvaID1ZYbZBN+/
K1gIO6KMR8HiohUj3ADbcgdopS4sYuNlxwn14rw6tXJf3znmQ4kKYa2KCZMKEp1HyVXAl6tD2yAC
sbMsYlkjkilBFTCmok++19fdLwu5eKl4DNSOfbSSq4C5PJUMrUrziA+dJd7BCzsihFfPkllagLca
xOVUiBRTQ/Z4AHqrh8RSAO7A1bP7wBs+A13LfyjixaXcZtZs4ggpASOp1zASBscjPrW12cMkcy/Y
tUQU57sMmRQVIHXX/4YHaWKzzieH4FQGBDhTS9sUQ4Hev/9qkgE4cK2jxRwGvHSt61NxFjxgyrAT
v9lNhUUM3t7CzOJI2dMAf13/FyWL5rmDmsyih4ufoCHn1ECjmochjYoG2yb3C6/8OdCPdDviezg5
56ppgLDaHv8wtP4WUcpBddW7D2QUDLU14rFygPJ83fGqWz95Q/vy7W94dsZJZ2OMP/Sa0MbBd+sG
DUjxG0MpryvfP2es9wHy1HQ4AjXCSNedDrUX1xZJAiHG7eAvKUdq39R6bkq0pIw/4YAIqEzqO9xy
4w701ab58rZpJBD03K1wX6dQvoBjiW7Zvs+XNDXCEgMqnMDxccrT1z6Z3EEeyb/4FI/hhc3ZEUTn
w05iQGGpXDsuFxHx/1MBXYG0Ke0uOXJgvGYg6WZxNR5pUZ0GFz4FvnjjowjoLZB/WB7xdtyaUTcA
/bHsZIt7UTn4L0YwE0PvQ1FHm44T2P8ji8MPIPYkgAaxcc6HjmVGiD037jkXLZaQgx3dQMOy9oPf
AeiPIU4DlSVGFwUX348bg+HhBxPXF1U9vOL7IktPaOc7TurXf04vGXDV/6czfLHg1jBTblyB50eD
aIz291i7w9PyqD8pE1lciwHLB56g4ArH90D5LK7kddyh2CmAN4tBWb/0/ELG0iYylNAwqQqrdhVE
BSU+xbo+6O0V/EiBMPIG2EDI9cOBGETI6fZ7iRe3n0LMuhjlvV54Jbgu99jb6QNsQPx9+419hrJe
VkYsA92QJPx6rUrKwP5eooyiFeAILpehKBHWLS8taKDlg24HH8fZAHQQelbvrjX/JscYu0WA1nEM
vu70Mm9JSchjB5JUcEW+LB6IzqnnmJ7xuYAPKyvwnTkxT4/HLX+muZKRIJ4RNsHRIZAYZHTwqlLz
lpM9B6J97DOE4ZtH0n6vwGMUcDIJ5PLU4Oy/RhYy/HW24ioUmTNbYoVCJ4uoTmJLTC9zF2jyt2xK
rk8d/Fxvv7X2+Dq0AV2kLP6IAUWcXvPUHPJB4GD1IszZ5LKIFHpsC/kEn9TBSwRP6ybhgIOS2KyR
p3LPX6+Xq0YQVHkUYVLSazgOSCNqPbie1FoeUfL/qc5ijqN9321PqQmB7BCIDeCXliPvqN1m4Dho
vBopt5Eo9QgZZhBy1piL4uBpDbHsjN3y2zlKtYM1wrlY+/+N30nrXL/qoyfVHTQWXy9k/U0PRSkI
lsAWjrWE6aTcoDbbJdz0mhcN1aZNUS5yxG2Of3WpD2L3p27LuCSnw7y3Napm1nMcHIMwh57mnCL8
ECiMHzNp+hA/mFcV5ijmj6Od9sbE35CAPL5LHDYraNFYpL38zohCXOMVcqcCeHW2sO+pn/2LvhCN
O6/YLVMt/VXvojLt59pynT4yiLDcsA6gFEc+5YFiZEvG35STOBKdMV647+wU/ZXTNFtFD7I/d3/8
YE720F9PekCCCI3mhykkgjycT5teOKdn3i/xczKKQ8irgF1+hF+b+ZmrkZRCJSLaigB2sM3idDQO
3HfML8P7nfLQlEZ0UXy/ykRxms69+INxd7jYZbnTmU+sOVRtD5bIcqytKGP2JDn6nkfvoxu3K6h+
v9W4BcKG/6i1SBoToWW4URB3ASrcB9Q78RX0r1P8UvFNq7fkcqTTDmuWz9MbZINChDLgSMN4UPtF
jZg3m+SiBur+NuwmBN6f0TjNrXNxfZR7/P27nXqUIHuUDi+opoyykRC6Q/Dy81LagtTmXrpXNvWd
GgqWIVQBGGZtLlpms6iTawu3AeBgWRMmTtw1BBHtT7CEm25XFXZN8QnFle9CqaZVziGwKMv9tcf1
oviuWXVQnJeTiHeZedMRSjxT2ZTpAI5KpUjUHKhVdBld4hXv9DvhIEUYdbogRJZuq9ngTZsx3rch
lWKLgEyor0z9kt9X7MnLditE36x/iel5gwE533bz/yKmMEIB2aFfYQiczZW5Ruot17ZqdV8390+q
vfFLXFEmZvZPh4Q8giDte75p6hkxe0hAFzTxGcdvGv2l7T+4u5H9MkSPqa3fz57opMWmFWDjQkzU
p9s3BO/P/dQroJLQuFPkVXH6eAcKFXAFclIX3s6EHeRl0uKgLaycUiupOcmZ95G45cWwRAWnImTW
4Merucf25l7AfQT44pplvZFNer7nhzLftRzslJxspPswYMIzvFAukLe47DJntJAwxvfY6gkaYIXt
iA37jjw6M/eiW4CLc8qgdgmAAlkl/A3wY9BGe7nySFyZyRVLil+b6WAj6CjgaEGSXoXi3JEFdlbE
goqos02nh7Djgn7maYIvS0TgNtmSI70uFiN3L+1ZHMKeowltEbwTOa5DeKpGEuJgEuLIj41Jp+tB
Ts4DhQDulETGNMUDnWyIapvnnybuwUyVLpuiUQlmrOYIFwt+UTUAPTH9EmayHdqRJijUcZ2jZPhT
NKI3UeAqFgSppnkLe1axtxk2YzVEDxv36NRsE3j25NaygEJWdghn0e2FInS+6PWGZSN0cL8/hO6q
K07J70XEPbYprjRTTBidwsMZKOO/wW6V+DiGfDVfbEnjkdtIi9P1dDjOG25VotCDQdfl+bkHJjzx
oHxtd3czgK7mtj34UTGOtRmiacPQOTJuY5zAcC78jDjKOtShzPB2eqq++yQLJH3GwwnIwkHzaWPP
y1Po0sk+ajF8jJz6sJFgmOWuL29Ej1paRTFcMprAzc3E6UrV81qjVAVKPphSE4OUSexQ02VZE8t4
fMqyplUEkkucYmrF6SZcbuwlzEtGh7o1td+PBmNxnDnaI7XJX6NqYP5vAqSEbUwUglg5O6qEzMj6
LqgrPN2GUNt3EhJtX+adykZ9Q6t7csrHfuWbIBeoXnfF7B6EzPrvN33fmK+b7ArO1Y/qI1kbcUXF
3nDRjQHL7QKSSin0rUcAMKMWmAUyUh1jDZBPzayG2mXm211I/VfZTsAhSy5XZGwvUv2O2q+KFl6r
LgLGx7wNJc3dstdLH0kUVMiUfSdjGvdf8R8XpJfxhCNN+QrivX6bC8RXuMM5gHt2rJ9Q77fI9Gy+
FCldNepCheRKiMcC+CXgfEAwW/ekq8qZMQZeX0C3I3p547ZtK9uUdcQ6ThPFXwGX5Cq8hmSS3RUc
FWQsqkylyI1lji0XwnI8vsKgs2GsbAI6CHT+HAIhjvUH6rSOP6LmT3JHM1nX6bsfiCdz3MdCEuX6
xWuKGwKeZvm2Jae4Qv3SNjKPOL+GK6qAxgSr+uZk9LT+sx89dkZRxJuu6bnctDJGlkCfbKK1x7Qp
LVyiWAFH8XA7JoW/md6tu2X9oUTMba6wOeT0n7QMtxQovy1qwmZKxPpX/nPlgsZ4SFcKzQqWPg/3
2reoELoQlnulpZX/0WzXrlekOFD+QfZSaJVffTzTP0Ht5Mfw8mXUvF/zf8UGZGbASnFGuyT6rdl/
h/itC1N783d/TubMNRw4WzuIP3t3qd/EuFsWe/WKbzj2Ln1Oh8hLq1xORFyuRON/4yU1HPbXe/tZ
re217029cA4HRkEHg2AmoaZTegltTf/3g+rAUJ11K8dSKZdsNohrIGDcLDc4aGRKqkbgtbmbodKX
SW1XqLbaNdLZnMyWJmxOHB06za6GtVhBgX3i1FozrEEC/E1PxvV/tLpyw6n89Lln85lUfa5eZlYv
rUmdsWIbnueGOae03OK+8vBuYWK3vOlks/UEK/RfIzj2SW+KYN2w9sHApTDs/hV5QaMZ+yXbMx9E
nkmkywn9Em++y71NHQpucz50oMuvWLJx1hp3xRAC0CUiOi+jp+0Nrv4v8McVKwl0nAdeAt448+iA
ZqRqzDJItpJxKG06sdq17+OECJojacxxqdRjnbKKb16DJPZ9zxOMorGiddfujfsBMcoY20V1n6vA
SU0H7XGJB5P2yYq1JZf0LTBk+r95LMy0HHvrGkalTYDs3VD4tDZVLwWVSbOsTPjiX/CgcuAZbf5Z
543ksLHlnlHnXUeGIj5CrK27Ua1tJX3d1Dtwpc0GN5DKlUtqit5epk60rodzcQAinM4itb5Ynf0k
ss1m26Xxcyhz9h3mIgd+fW24buBu7UzRiu9yzDmk4V1KCbX30OiCGlZaPxjX8I15w62MryRurNXk
5M6+le7SThbBsX+57hXzgeHzYkWLSz89cQmlzepXqw5iCjcx6fL0+qD7sFGx5bFWNc4SR7Q1AQDH
LUF8FdGa5fwo1EK3ONNu3ks//2Do2+JqsIHYrL8rbVSfz98TxO5KQgv1cn6Q3AHltiMtwQGxrqfL
lY8bF0aSJkPtinlRbekH2cDBkTd4UvuaPDQg0iI07PIHIyI/lA9D+ZjejgAaNxcpJJ5tPLORu8C5
RRiknyyT7ZdpUbCsMR02Tg5xQ1po7nZyiOD5d5EJllNlGK8VN+Ig8dh0FlzIAR/hOVdqLRbXJDww
AS6v0tpw8HQ/7hye9QzEtb3MGmjk10yL8H3zbpelLjJHR2/i1ARUr/RbgYmyHJOF6+ByEYkIXYJc
YK/ZF4EU9JS7PhGEZgd7zZOJt3zHJNIbmb1xkZYU410viaCoIoPMaahR4efNkTU/6YaXYAxMvlxP
gibpkHJJ0VQJxrWr1+DSMiEoacUSZX4dm7ZGg8ZM9Jd/UQXQjTy/6okZ+/RLuMU9fgCGCxwTjyZq
L4kmarxYUfOQ7wSMVceiREAIpCBcOdSU7bZZP7P9e5uO7I21IfD4yDFA5o7er+AsPRJVYAFzIHtN
faL1rToFC/rTH0dLeDKJUhNpkZjt2xyQMdA8QOHa4vAZrqn8rTgqRP5P/xo19V8s8v4gy9quQBJz
7g6Gpq0zSC4NnClLnt9b1Czx2nn4INkiYHxfpbL132KBpozw2vHTBrtL7kbHotRKBXgAbXtuON6q
eYHtrUjk7ViQPHPTrMxFXV/irj5jw7sG8Ohl5XPMaAsR9CfUzTgbZVF6nF0XXDGGWrbvqCatst6l
ElKShhzcc6RjeXYWbvLD4cwyplfHRqAlmbxXxHpdSy/VPi7/8TcKQXtCjJ/8nMmUo2fQ3G5htmgZ
J4/pEOeHmsm6Cb+ajkfjxpLF2hPp6cVHiIeO9SDg4azKolC/1ICduxBP+2sOk/Cg4XQ4dbA0NLbw
MK3w8cR5kmtTsmkalh9QfBr/cHR45ZMoaxZZgeRN6TmQ+RpLbBeMS9458pMIn9atSEtmq9SwCaPa
qHumHAr1ZSoOyoFNlZAeqK5I0mETwm4zCnow1zNtW1T3beAAjN+uW3CuQGwgMwuaWInfoDAhaPKm
p8Y5Ea3BeX5As41XAk90cIxtJDepOWXY5lrZoQp67aheLYby7ZjZfSmF4u7kjXutT1tdQrFA8Af+
Y3T0k1n/+DgJJagd0BhZSRc5XRuBMKAGbEKjaZAQL1pzpuxrfSxviBNRr6x50dAlPrr3smzrUser
y1mm7X9r4TqmpV8Ramusyunsmb+iK3eN9Hr+DyhvRpJ+J6gobHJ9UPXy9IhSy8m74UAw8bXSZQZs
jL05IA9iLCR6hzZMVPTPCYcOghF9c7tv8pfOs4QAQSSOb58ZvSJ1174yD2yXgmIzWMHqii4lW5Ix
J5s0ExXzB+2DslQcZ0E4K4gn7vjpWdT8d2CT1uEXXw4VQepQp23AxykZXlYLH97xzUBclztKD/iF
IMm5G5+nQl7+RqbtpbeQ+Bghr23xmCNmKGk3E+AAEuTheI/J9f+UM0KzapdGUb/n8g6/IcPsnWMY
7ck1MEXug1flpTHldKH566cv8QIVhCJIsOMpC21cJZQ3TvQMYAk9S74U3kBa1ljfhVuL/CoUSYjo
n5t0Lm4EWbXgtGguB+ZGXux7jEGZILDQmEE1k3HXugJuNUqXgOW/XQjLLcQ6he853wMGXgKehO6n
D0r2Gd+ufIywjHqZollq7BB2/bhkET28MP2iDxlkWxeD0zL3GCbT8EpP8aFh3bgpiKg4K16OxjU0
RVAijr2ro4q0doMl8MHV8VZaxfbwzelofudpmY1kDRzC951Z9JAR0j2qsswRLUOShfimgx/rApK+
gzw7eKHsN4kyAbnuFZpBuF77Nvv2lnYvumg5i7GRI2WGT+0uBuCyrfGSLHXy8cucwlO2Qn0H9/RW
TzZM9DBFlrgL+Gi/PxqL7qBXgYiIrjhQO9haLWmy4juczx1dapvoQ+nwMQOmFUyx/U1gzia5Lqle
KaKIqiU6nAR9reTl7PqXkIrDy5eEWT7O3KkjUoa/B1f6KLvxIMup9Jug7x/Q6u2J5124FjnJR6Kd
iPq8WZ25r6r/ZuSqLaGAUwmy7NXj5vtP4yWERwEODQYpNDL/Lwlhrp5snW5Z1LVOxuDNxZOFfSQp
vgzWpT91fmU7x8fnlw8731HCK9DVnPNekbiqSJQI386Us9iEiNz4EP+5fFZ00Yu8b02Z4ohmycrK
VU59q+7gIQMNo+6nL75s7kfwftBBrAXvIJTYgCHQ3jvxn5NcPyJam2LVkIPlPa1WWnMbaNWEEkEF
mDWcW6c0jw0nppid9dS08JJ3ZwYxBdvz5WC86ZRndoQTtNbRoRN1A21DFPGsdodRUUS64Qcauosj
kTLYsfOSifYdJqXlobG0srcQ4TImpmDz7VfuNrcrGVdrZBNzmdH+ls620Z9OISaaWIQ2DmyPlFBH
AWOOiTaHSqc1p+gan1/IkJmWOIUzIwDj8ezKXZh+CAyCRAtx8nttmhBjZo7R6xeTDGH23eUO1iF4
VwpXGMC2+OyiN1XgTj6+3ZKpeefBaY6Kt5yDr3CwxfPOvRH6whKM6Z8psqGroDIdJgHpzkiFBK9l
la1LG90GmcJ0+TrhxxaLEUzU6pI8k3q6SX66+bCEtMAsnwZu0EZtx01I+up8v4Apqpbf3o0+C3JB
FEBZbPohceVkCVmv1wv4tuoKB4TmPzVHa4bk9TuF5Ytq9+S5loJLVArgL1mPQcPKt4QhAydyC/87
FgD3E6DMlvkKdkxj+LVub9taH/Clc2BoEguaYTGhi9KQQiqTrtL5irirdG5wVIxpmG9AaYhXCr2P
/bGbihBPRFk4/gBXMDhzp2kEb51LpbG6CE3V3HKaVcIzbX27zyWjolerYeR//55+iIpj0sIZP2NQ
ZXg4cZJopy8Pvxh7Hfq5oRd6iWNnEkGrJCvH6JgoUd4AG9GvQdl4N2xxOSs7BpmXZuxIABJjr33B
Ad8BtTtU5qAmMJJWnOa7fZqmXqs9dHzcr7kPoejaTYX7ObirmCf1PpBwyvHIsvxh/daSVKhsHBnW
S2T7j+t7Fv84fRpjfotWyYBU8xeebbwrhkD5GswOF8k5vkoewTgHQzAPBfchFqte/9VzaQbzGCs2
NVluZsN/gK1yobRroKq6ezLNpoIm2/XH0GbcBWux5EKtApj8LjONpBrxFonpPkrTi7cpvGEYp8WM
06u6SAITmvhYduCNQobFKf/n8WP/+35iM+zGU7O81DVXCLXeCD3RCG9VDhhoMmsEvRdjydHuZhUD
DE39oD1scoigmUg9PG2jMX81FAGODqNwCkVn24t/8D1BXDTxWXpnhaFI/Jpr4e8jQdOUVUWP2hOW
iwB/XhF9X+Qj8EQRAsi/dAsMyEjm3m6Zgj17JRfqAswUncfWot2WdvHivS+s/6WKO8r9oG7noFxc
gxcNBenetsnAftr5e7JR6NswJQyNhe+LjGOh2RVzP/+LnXj5PFBWZoI/8wQLM40GhtdQnATpNMq5
F9xHF5s5a25sV3D6nkxqRksR+6/OHWJPl2IIGJSp0y0I8Z42SlpwVSw3QO+8X3CPIlLljN6tf805
0GVLX+wq9junyLRU/odyd5BQDPkE2VgSclTMqO3jMaYEMwoZg7X+fQVoasSlcqfR/KMX3WfeStoU
awOuqAodKaaQEakPHTsz9F8sv4AKix7q/0HeLBvLz8cEEWnf4/a+bFdgVpQPKALtvkJArg/bBIto
OxluC6q/qZGr4EVxyht5yOEjmtFbfV5T5rhFpb3dhk6AnMZZN/EwqYvTt2X1gPSI8YgaDNGynYxX
1WepklflIjpRNh3oVeT/DvBM2j6WGfrF09Vo4z7CcUKozhmhpWSQGM6lCq39SosXIcLtJnBhFR5M
dHFz+++HIRpm6UVx7Ga2glUTC74Ejg8UN11kkEb86HBE/LzyEVvbhwTfGmcVDNd5p7lXjiB62t7A
j0hU8XMvjsOPf5EHPmS5ccoJ+yelLhWXMonF4eVgTI4xW1I/d/NqmcMYiT4CMLWsSOEzbbyK2NtW
IbqIwc8bv9oMgV3AZueLId0HDhBkfrdZpQn5JBLk/FOL8X8Vs3anVIutWcettDW2HIgFj/+rTXvz
9XX31feRMLZu9PLt5QMHRryTjTaJfEVDHDcSS4WHMFZk1wpVCg5CgzFlBXRt88HLmkG1My69lfx3
aZq3Gl1vTXbYlUfXb6mXH+GUjzqr+YV6XAMbtapEK/rCk9YqP9eJaMPTfYLYQ3nfsHkZp6ezk0Hg
tk/XqhXRa4VE1yQ5IHT9ZXiyHd018RkhukKIg8Vqp2bo2DX0T1AStaDLHopM8rlXm/TyOghLIRx7
seqwhSlxVdefJQRjar0aT08CcHSFuGIXljmV9Ch71k6wPnbH4mRmcZpjQhs36t7qepqWh6AhdemV
C8fKC6D23IFdxJKNwsqFouSdrcKX24z6N+Pu1SC1Rbidcs5PC6GONlTbK1JKnqWJ+FtSTOLGozQB
57wWkE+DRirBJ9VJ4hQhr48qa7aZM84keSXmoxOz4OF+oYl2l864eOOmzzVWmNEjhRrhhewLwx4/
1DARtnap6YQYMLsDu3UL6xktiEx5drgbhaONJy4aQht1iLe1LbpxMNPA2xxyaUwXgDUvbYq6y0nJ
+HLqifH4mNqOlWutc3JEErhaO64u+9xTkh3xKv9Uu1WJIW5wM7oWTY+Py6CZp+R0reZ9U8kmiVSo
A9bmn7bbCOB/z5K5H/gurpYNAae9oZyGXJbBHiJqpX+gte+JAf8UjQpWI7Y3GBum3VaRDg3q8d9I
9BUwJBj0oX3wkWpAWD9TBx3W0ELogA9+U0XAtJQHyvzD1kQJczHtMA7227YPknGqr4f3FFMEd0Ki
LhdeBaPNbZ6FwmFkixpt6AZVUSlqYYhbOLtaWzG6BDvUGa7iX2d/9dRaT2JUlZucNyP6nXLkeZm7
qpSuhZqnDStw0JYhVSV7neKUJOamVEgB8xtSbrX5LPHp6g22hN/vzpPo4yzayE6Wl6qPeK8uco80
E5Ub1CBRv7vXR2ch/+CrVCMuI+3wTgrAnjfAexFOxd0HgyS4M1WuDMFjLn7TDw2Gzx5plUxJzp0n
MNo7xHLlJxCGCjNjlBYVxZWhOHpn9irA7jE9XxVKiDqkOnA7hZt9bUDJ+LiIOWsQOesyW5z4JEmo
i17pWqtzcNG5ZP2wiC6Ssplb3NFSfTlSHOvAHaHzzibYZkdaazfGT/TEB/2cu5WrXcLQLJGQz6WP
bDR023/oseX1hKLB4E3Z1TIu1E7qRwY5bXRnfp9xkX4bXTu3WAMQ4eGILGgB/qhLNqww02Y/rmy5
0HX5rJ/2wr2k3o3wYduDsAe3csvJHJZYuTII8vlxv6XuZAbIccZrHCRK4Qvjemuo/EzOPuzfMkud
ui/sBUAe2jRijTNKyHwNPz9wqo7DAqZ1LeHJYvBH7MSKanpP1kTRybNcES7Ex9stC9iNAWoZ0FAa
sSlT+fvyklIkj/0tzp5QeFHQpWT6rMya6xGr6tJt+AfGpn83MyIBZPwgZRPN9mZKweOMslCD6LkV
wEy9Y1dwC/h+1RC/+18Zdwaa73KMGYod1v9lI13EaWisODIvrYKxrcSO27D8OzthZEMMjmUxLo7v
B4j7Uw7Q61kszGYJKw+FyNKHS7W31JkV01JQAm+PIm+YINKStX95yHLS409HD8eRrJc/dzOJ12rE
MSzT8061XtsHVJEcctwLQKw0HW5VI/UOAZ5XkbD0Ilv90L5jMwDjpRnQHucqnFqeZMJxHTlMu6Er
zv71FZpGHaKLkIDIFaGiednxRMd/ooZDW+8kXPIiVmd52meLMJkM8nz/1n0Qu/SQSZm2P72qV1VH
gLkAExD6tGxnludbDSsQHKv0LxzyBFqBFqJ4/nN5q7TFkLLm6BQZ18Z8uoMygYwMNaliccnelW8L
pMia46E+VS7LRcbhyB4/7O4fAMjmLrNFg2jIF9Vxfa7v+LWoC8UoESn5fxFKWlLmJUUS64/gLJkC
GFGSAbzLhZl+HUE5H7cA+60hPi4Ez0QTDoTzV0AGH79W5/rZ7susZWPsvepQzd8bTpXa6KZWvF/a
2LuGHaIsXuhBwZ4nSjn7oDPjtSI+lAvMUZCf8gbczxMQTWAwBvIwAyLfBJ9JxbH9Y+EhX5xgyl8O
cnY2qikgXrYhP7HDtZHScNeLMGSCJjZa4v1ceJTSGQQzGI9N6yklumse9MxqKkpIRYf9mOry9fHK
lSrRYJLjJ+uAKf9f1DPeOE7gStZCWdscbcl5F02Dqf/vVzLo2dQKdFFU4btTUhPyPau8e0s8SZL9
OWowFmy4QOQ2ksid/5zvFf6Zh4gx5PNLzHrli1Q2BEOrJvoX/m35khnCDkF1xsKjYx9aGNviCjoD
IBr/RRnM4HZgAmXq7yY7cLtHoasKN+/z/0vwEm79drvS3LBu7yqQc2KhcwGBQ1UAJA26kapwLcnw
9da6dHNrNt0g/4+eFbv96qBmTbfsNrS1g7dGqXHEPCByJ9eh5tIjAQoROO5ZJtDWKP371ZZgEtW/
m2zMreizTEDhMyVttsei7Z72JkBVemxWRYEWjGefcSU48hdgipg5O8MKesCNKJLZiSq3xeQKJD41
xHLC3I5P14JDtsxFrxWMiL1ToImx4TcOUYNhtq+CdIr8c85m14uFu2jEOURFDzF3BlV0JYxVeRlp
bXncy8fLBE7a9rDgv4UxLaOyJpVA7eLUfGlLclO0TUfpy8BypV0VV2qaypda6vEotmCt7HEjXOu3
HsULdFcmDEuP7TdJTga9grRcS+jy3tYbEkNGZIVifCAWn0VAswl4yG8TKeUgoVoIXZu3JY+HAgm7
Ht4MiJjfNGdDA/0fyk5TcslQPHTKxapYUfWqpvFlBkQDVgVp1d1EXfVma/vURD/z5h0dvk69mtsH
tIidaOg4XFaofU6k5GYqfQvzt3IeCFxpHbuc/CvBfgYT5TgG4BpcPLJiYMk3qDax2ehB3jzrV8U0
QUSlYWjdL+MDSs2kDf6af1gKvE8NVjyjNHV11Y43OTgUDMS1WIpjKNqKF2vYxx0HW29W5ztCusR5
TPruylZy6nNk+mKhfk43Xp7HAmgZy4lqx0bejLlSRdq1foaCq9m6+OBF+z+ZWkHYK+AUW0kZWw29
mbW1LZ6kAg9o9cAqYMDEdcgAqjId+vLAAdUF1OOpxIOEaPeeWEatuu+GX9SrIXrM3ZhJAGB6aZ6+
rKW6qHd4VACzmyWNsJG0NqVFgi5mQ+IJT//T1/mUG9VmGmxoOw6hh/RW0iRezqCjZIdeISPXpHqO
SegaJLTZacUg2di28RDI5djei5IRVDTQZ1Jhc1zJTqQ3+8GTCZxh5lvuDtSM/rTJrnBLhQpkuh7o
HwhnQ1rRFmGvqGat48a/efBAaBoLdqhQJjQB+/PrYrRNOypEFixuuQCh2ZC3OTFt26Nd90ksnMNT
Onny8XDp/seiLuaCQM+kiEEAikwdOhaB6csSh+cIgimv916HXDyrOC0+q/XXZ9Vh8jmNwrVhVlLf
qbZFDwV4V46VvLYrhnKnekI3SnQ2a02aH+lkKQ61IKa0+7P4ylPIFmcPrwvuIgHahTEkx9+NRKi3
fwj6dWATJR3eHmISyRmkoaaEknRfoDAW0vfRwp5mB3/8Qh+nvvD7P5syNRM57MRNgMCEW+H0lEQA
LAD+kPKKbEnlIUon9nX+IY6oqpsM8OglOTVDNhkqmoVQi02fuw0btEoax8tTTYCA/PBHB9G04aSZ
Q9abep9Vjw5GmJ56/HVw/GaTdgcDCRHsHi71tYLXVOOqzW8uiR3+yB0d1aNzPveG8A1ZwPEDEFcc
LNhuvX0qIBw63v2VhclnXa4wmzLdqs3iBRIew6NYzGLEWuCP5mK+3Z0lLUA8yRR9ycpkq5HpOXLW
HXiIMiAVGofVTIFO2mgU/EcUJ2YtOp57xeotFcI1sdsHgUXREN95/jFhiaW5INoLdcU/zrj/pgB2
4pmh/oweUAcoBuYVIZ9rdHlcgv7cC/u3s6jkRx7j3871NttSb3ylVcW33vtqnF8xydd6a54BIKYc
cG3xcT0p2Dz+qSO05w/L1rKHFaYwWv0FAWzO2cARIeeZ3y/ll5//VIBKgqeoenyW/XdG652wkR5q
F5MGTVHjvBn/48Q4KMFL0S1c0sV2MZ6fiWJT55tNahIsXMD8/OwhaY8YiM4Tor/Be2qy+s60uuIm
4YwHo5pP68H+6/N8nl43tGj1rvBrE64AlSETsDFJ9pfZ7NZCXlRm5ptuJNvj2y5AZodv/C9EBIbT
0tZb+7X6/uNj+KCuDApnJDBkG0XPVvVwI7BtbrL1/hCj7o5WDTTiGRup6IHIrUdkLwG2szNIKXa2
WtExxFpGz1Q2+atAPRJEEAtmD/3efOr7N/tRmEGT7d1ebkvNkcU+kS7l1GbzaSqLfb4eUGTRPZ5G
oJMSOtSQtKlKP+5r9ZLrxZvBxJV4nObVAFa2NaP7678U9Wg6U+Z7rDQ21F3Je/FAtbRTSGb1/UTD
5qi8RWn5ag4sP/qP0Vvr2CF3w+4GrYanNYnEE6A0IvRSwows7jldNoDm1d/RRpQYuSAF0VxKWWHT
wfUmdSAWFWVw+eueX1PbnGiSDIjoCzG+H23rXaNHRSL8WhU/V9W7W0WqJAOwol82lWLySpI9TtWU
9RGcA+DN/VOEn0NkOpT4AVh90LsJapC43PnLiwFWrc05pVeifCTYniBZLq/RGibvwA/p2hmd8l9V
2K4ryJ2Vn8SPmhJn5jxJSQBBX5Ik7uHrnOrVBH0Cc45H+FMIupeFLVM0TNH+hVMq1bGBV5xAUoz8
H1F9xBsyeyMtPw1ptV7m9EF3Yhb2oZbxFQf8c/wre8WsSqfquQH5AUuKNazirKaX5Be/ZyHBXepj
G/Q1RHX+Kb2f6nw+K1pJ2NMO1a5NQYzVxbpt8jMB7hThRreRJYmx0nwll6mQY3jqnVqOifj4I6iv
emhspIEmR9ZocuvAmX5kZ6aIFh1P387b8jUKHhBSiqxPE0vSp1SxCiBPDcUoQGsZmAsa2mCE+Fqs
KuTgTdMjeLNU8QhHOhlM7Wfm6RBI/54K5vBPO0d2xPneev+Fid/kaZYwIR6OF+6kKQSCbwBYV99w
goFpZiQARrdgifGZQsl0lW31V+j6N00CEpx2Gjya/rdGbRImK6FM6J5qIW1PrairqxoR8ddvy0Rc
C3pul1DNBse1/AG7PRFqNaD6lO34jM+JXxK7ENtUOh/4sL+BK0h25clsZP4NbL2JJL5ZnweFv006
DvVjMjmUy/wx6rAM5vbBp6rT90iPRcx3Za5IQNw0EnHKN9YsV9Rsxn/BAJCK1or9s0iuSzOJE4Vg
btrdQQSFLuoGWOx7M1WNkhEiPuH/uYYXZ8Qy7V7CJWpEcBmpiCz8KbjIuhDXGTMv8BpPxwKR9aak
Snj40vEhQEWmNPlaxKqQoItK+4KvR+YWIN27oTSqty0TqZS12Uhpmhf1FX3nB7woGwVpc+8Lgd/D
O1ejE9qDeJ3k6fospnM4/SkU8qm1331uPBK0Pn1K0jZIvnrqc4WoCJCEIc+mBp5UDeKXTX3ZJYBi
/Z+x8hvvaKhbngyn5prg0CBmHbDKH0ITz+Vvj/RFPLFh70iSbIUAZ9jML3u5wDK7H1TknB5qg3TU
1xbMqa9KkHBVnMPkXUQpMqNeQPGcGAbD9TyITTQGFJbayj8H679tpiKne0Y8ffhvYYki5FTC9cAy
wzhB2RLaiPmp4VqgASUHoaH7cPARjHblKw3BnB/ILJ//Dpuu6o0//zWs4vWc/y1PyRk002c8R+2g
w6GSPPWj1GULpKjXjOxr3Oi8MJyxlW8ZK40nOKnKJrEIJPHlBBAeCsixoMEarM+jSAkHN8ZHl0Dm
Zu6vgi34+x3xxULpYQZpsvI73pl8p4/OvRS0quCsActWaADhjBRlP+f8hPu4/+WZMpqD2++s+2H+
PaajZ1LH/CwWDRTsgntOt3nIaJFG/eMFa5nEpwxpCD8sI/ZOHIzO4Ryg1ChSfPgj+sHYsewEQMz/
7Ed7foyQP15dhUqZOyYtUO3sZQiODzN9wltBwsB8yU9zgdPuQzbVoMDSBgVgdxXmuYymBzWycsyJ
GWcQEpOLeYcJUfdxb1GiJpqunOuWQWP7xzMVSHsYLpi0x0RKKd27bn3feRb6QS6WuT4gkrBixITY
FhkZ0VyKTYRoK7JpLXUpY3vvt6H8dPny8Ejx25xOmvFIRkV3IYSQkOi1IoAuO85q2jxN0hoYwKzA
1XVIBXlPChe7pLVpVbYL4pvIE7IJ5+6zH7lyfxbuDXMly2Hodcac3HvL6BRa3MRBU9+jUBdE/Zeo
XilP6bHpGJvRq7aEgJRiFSuGPYLO9pZTWL/jzwQnJDzuuFdbrGVJ4Q+ZRThDkuWDTYTYZjaObj+W
s1v+BZ7ZAwVyKI3Q6O0Nqkd/sAqluJDxUAC0bDhSUxSkxzDYcOYKatBO1pYSyXXOTTr2hyZOHV2H
DKDCUMZUu9kIUSxAH6CNyThK+dNSdLOHigqwAL6XPTl3eq/zK0WVAO7W8Ty4t8pnbQl2S8LrxAXz
OYcU0bZUTKaBY3VhjA6vB+2Jxsei/rRB1BevD4znVIkSdsgIGPvA07PDy88/sXAP/q2oIn3wPTxM
NY6X0cAqsB8a0Xf/wb1mEGgAlKnkiiwfKlG8+2nN6ZxtN2mxPFX0pvAipUKjHopd+NU8xo/WOF/E
/fONRbemOdkNzA3SuTWA4SlgphufnJDzLJ7SaEGjYQ0Kb/f1veG7EheRWaEn5HeIv3ix1CO9IcuA
s/mmfd0N4W3o3Gqc7QBhDG9gJ3syVbPapzBNa6QPzWq+LBRVMGdz8mQXHJ/Z7rxPDqlhOlx59aOL
rm7tmBa1EdDO64P16KwJ7RvOwv9syijFPWM+duWHDkZ8F5sbr3w7pMHnvDXM//agdpnUoN5gd3/J
tRwpkxktP1sIb1vKN3e1KRRDQECEjmVJB7h0TBWGXznfIB/4mrbqBuTDe3hXkVRuI83XEiBLFrVK
Ya3Y/xVpb7bf6jHU5h5bzqU86iZNbLM5F22gX3jUtGHQMK4tByTOyxEzy73QOqqLL8yqFj81e7v/
P6o6+3aMgjcCINotkfusNmDjAX2jLqhVqzaTFvP/aQEDAAudirsurPe2DdTdJn7+oO7g/VmTBj0Z
jvD4yXnw79VWvkKogaOZ11Al4iQtsbdCHY5kXhhVuhrcaVpCSX9dufIlmUPym79PIpQgmlNgQZUr
PY5DunWirOERO0clW2z7ZJcdfmgrjwNwM3XveLfdvhsFzdKfXjFHnsyvYpsPkwcpTuN8nZvT+ix4
vurVoLxySU+6YZ53cqxAgn4cUEWJw9UbiyEc5QiiPWnK/FRdZ3NvGeJXYDcn17b2ZjKWaaTJeJXf
ITQYOFCl2xPgvGf6qdncuJZGEktkIirzVjhuqb5nrM13PokdG6jgpQS2CCtIM7YIxqj3iIGVG4z8
0UFmWBCnH7fdaeZdNdf+Vnk6LnKXUqgIhLKaDHII92kqa0JzV1IdZWt2jvytAuq+NGKNyIBzrgwx
xUWeHMhjf6pYBVNL85dYoJLMmB7xkt10HvUg0J3T6IfgDeRstKszrxPo+PTgvHEs5V1STW4SCu0T
wmN22HG3Srkcaa8zcNcJK9J6zvFu00JV/eA3yChB1vhXfvdfk9YhJuRxMk4fTLl9jpvVqA9J/w0v
eVpp0PVUlxewY7476B8JgNkKJVFVwyXllzEGDc+1X7+qT75r/O5fnhjyDUOpukrojw7Ys+OBOnss
/p2//WDCDnA+89PlfsHkrFm49R57JY8k5TIN6pOuWod/Ot5qs0XaSBpkbl8b1zl8XjdynvOo6jD+
t8hh3VZnCJM/f0XFfXh6HeJn0VBcm/bRdIZcVGR2MMUqIM/cZMXEP+cAt6lIcvSLvjSHf/2lj6+X
rKm6TMAxa5mL9nICDHqlBFz6lFfKXcK1DK4hX5zbIvibncIpUvBydZr4epxCRhSnhF4d3sXT7FrH
DH1IPnusCO9hmNlZsPQ8e++SSox9/wWtx9D562c8t9yyE921vcPA5LJohPH3slpd0womFVs02OK9
sOM9m5gbtB7VBEEpFp8xnfWPHhvGgogHinKUPCuD7SqHwxcLJELqapoEw86x6k/Wza2Mgmxli8rk
F13RRCJApwqjM1dj4JRaX1ziKCvZMXgfD8EZWMNUSTlG/quC7aOkmGgL0G+Mno2zZKt1IwoF+VW9
98CGw33rvvQn18WivybDdxvaKpn4wJMBUP8Ty2JECF9rOZoswYwtfpStZvK/oK3zrt4tR3XBmPs0
ISTZ+WBSECm3UPBxzOoMxOHNUcodEdGo9fb/Gn87eT0LoXoI2H4l+VOhngfJrcnEHOmxVpKM5GLO
xJWJmPQhKtdfeMwN8/apc1wDDyKLGnz5jV7f5H4P8yQ0zXnB2FD8q1FiUy738U4JsC6Zt5laSora
o0iMc8jEyLMWm+hXaY1i1OhZmhAeiC5PgfzLcQmvDM7bw88XK6PGbYu+if+a5V5jgrMm9TjYGdsp
S0i9HsR+TGDUV7004Egprbh/wUJAIzaKlOTg5fDMAuhgFSqXbc/y4GunOLQMFggoI84WdBDRECly
ps4yh+Pvk+MJoS3H72nsBhnJ95QUaQwXrkphVwUsIZ7LKY4U8MSFKwYIRwQqIcH1W/oBwkEaGYqj
vBUiFOg9OlPbfv5oVQE2b2HngXhpvn2M3qLZQDa4U+fHYTHtQM2nDXyICcXYuJQmS+kzvPNc5y1u
7Z1aA4cWhRyORf0YBd3zkXSVePuRod0Ba0PrHTwhih3yNDklQ5wripGE46dkzrdHtaLofue1Ee68
ookTvc6PHuhSUMvAcWPMlZ3VN2odXcqMu1NG2t7uI0D54wQxwOhUi1+5t/6HYDBK0JZ8mOLwCPVd
B7YpoQg/7U+qo6MlO3EcR8QgJsOusZJrITiIKd0LyxBQvZ/p98D0LL+rqC5ga5hzftZFMqZhed/7
MpaQtTCLGN03Z+dWUJxk/zoV28MzkhVQ3IG3FunHPsfrF0rBdnFo+2i8jTVOVBwXNU4yD84tl49A
VsMIIXaVpfO7Db8pYo5Zpz+lhxF9JCIeGGnpdaDIQDSa0uCEvZAbOo322O317PXcOCr1h9J97yiC
U5rihH3MPRA29rutzHZGYqFvxmofk7HbWlX+vpGIlyXg5nqNWDdE4G7xy5IFnD7LSjzQBfunGNKC
3sIIzerkgEuuUqyMN6blpXhTyJ4YIpoKO98t7A3ONJoYEN771svGOMq7JSU1SKZKqzYeSLgqEfiU
WlqUbxNkP8zYJpR7YnibKXTQ94+6wNogwPrW71udXm9UEH97cXS3/WEekzoMG4OqD0K2ShUQAU4J
X5eC7jLsbv9xHH0O0GWniOF3zKOwu2YHMMGZnz0FzKan0mA+UecoPUIOajOddvQ2irXnFpU8LQwL
iTjrmjPgAnJ5g6hnBVG5ln/F6MhYKI6mc9LiQGQbOtpNsDeN3091jch3iDec7sIh9x6ki8XuYS8P
v7/dmNYRhfy2WxHPbLAtK9saaUXCDL5aINu1YrAS1pbu9K3nqE4GaE1dQhGc1RCHyHqLsZdneFZD
L7CUYSlBQ9472usAdco3d8nfmQ/i3KMg/pNLgb+dSLgPpveqLlgmJ7hfRvsGfWryGouapouJCwq7
XwWtBceIrsa1XFfYSAvrgsKI8frDgExRAAwx0L+c94JZR82amhNYgXYjSiYWdGGdVdiB6Zw1YkOv
UsNqI4qjVu3CUP5grO+VSTKShKXv5RAjIp4x0WkMauw5YhoUwlOw6ooETodK8XzLnyQPRn3Owu3w
GUe4SgJtWCo0TCHd9Wn4CEa+nOUASU75l0yYVTyF7v4jdoKMVFwhNz04AwuWc90d0aP7Q1sTWMDk
Qd5lZ8Fg2OGz4l2/UsxneGLX4rRjojdMbsW33g9JKCzVSqp/mQsm/sfiuZA2BQc1gzHziWZGjIf4
v/YKtkN56gGrZWfZ0CrMd/NyopWdm/um46IbZCdflRuDYgeie8WJpRm0f2e7/vGp4P2aJXVDMdAS
j/Nz57F4TrFcy31DBvRhDJLeF5XtKULj8fRzluUzMsCyf7L4856rV6nXye/hrpYdnk8N9Q12Uc9R
5HT8nqzCPOXFjLdlRuUDuPbxd6I+/NCAOEDl8QZOp+LzxvO9A+La6/qbxcpIk5q7rUqU3UMK8nmg
cbctfhA0xsj0cdH8jyYAC1bF/Xu7TLnPUqsctq9XkQ4uhNseumB6onLkO0XIT2v7b/Q72OAV0uHl
bAot3H0NZ+fxK5jvL9kVyRSy6kSuYglCjX55gdnQy04b5VxFw0JLErc9zf+PZDNX4fUSeDeWWMWu
optwainpgBgHN9Ap3FatXq22rjW6Dt5KiLQV6pEGtSCE381QuwLHwu3j9dPITNgm1SepEqmF8oRL
0ryUKtqE3rEitK6v8wKi3z5tjvXhaW2GKRizid4fdgXi9edW+kQQ58O3sCXIeiaUYOYFyRmEqbGH
jjDKTqoJaVMU1dge5G1hdRQ7QXMjr+lAkGoUaUkXMQtQ6HcB86hegqGO6pbwjdpnb4lp/ao29z7M
EsEO4VzyhpOAW+wiR9FTNxI1LXFlaP1TTwYYaBPeFrrl7qHdIK4nMjyKl0qgQt0oxoFvWm4PF0JU
7Hauxp5qTCRD7SUVzcB0coABz+Xtt4VJyIbBxjA+AoJmhEn8789aMQM4kc5SO7h1fzte82Gmo08E
ecl44ntrutZDTkQVa5AmEc4eLzcIlLWNWJY2xlGqijsUhNr0zd51lZdrJOQuEN6j3us7NMUJ6iG9
hxkfOHsWVrHBW+WSXx5ARapyIOTnHqVJeodvE+ZaeN0z6NhMmML40Mn6SzgTaqDsyiER1p20Mr+D
pLD0J6a4mg8tnWWKkrrR8phzVKP0MYex2GKxyfGBD8dHl+OPBxeX41itBKAKL5KzmWt1rmFtX7jF
Pw5qSSRf1mEvXdHxynqn1NHaNBOFo4aJj+OyTK+1IaWdDpXeSEow1FezxZ9qie+GaMhP6V4qXUWB
MHsAeT51/9Xgqj4ZpkEKshBN0mlV+Vii7EAz9oDKH4Vp2tfnZSD4meI3JKJKRsBfw0Tte8YUiSLd
paaurC1iSwJSc4h3kCowaWPEkEGPsurPQ0WOO/i5VQVRGiowb8XruC9GD4UZ1XeDOE572fHvq+lk
pcXIFyXOnqMWW+M2J5weQRlcXcZVDRVAwXdSQ9M8fli0dvUw93Ng9AEupmmhtGWXiHFaxKnxpAat
W7p8h4i7xtEQtgj1teExRiIfBBItu9aqTZDSwI8PNNYZPbb5PrDx9krVuNGhRt89q7P5BoiHnwFr
5pC2I47Xtaf26vtVVF61crSdVxQEf9zX+NpfmOG+GmXkpYflbdpu+H/JOIEP6jLOnEihxWPc5D3f
pudRDPG/d1bACIsTZN8T9v/hMiPIEloeDg7khmhxkBts6tOnUWtfkPL0j+PI+Ac1Gn137f5XAgpL
YihH8wxZLIEVWUQYFs0KDny8sQ1Ta+Wyr5t4i4QdyGIxApAGnzz+/p/xRQDvoAM1DoL8dr20yL9C
PZhBYvtrRnglE21I2rc1bIhi5noF2B6Ult7Vnh5haoKLQPteb8YuUggbPprvJJwrO8IuGkMhS51z
Zrrjc3b4UqKhkC+AjIiopyg3rl6NKUCO3ZfZDGyIJKliBq76yrOCgG/s4xaPFxt8/CuJ00a3kB7O
YuBnCKmch1pFFiHUaYsA5Oh0+QRrrOVqWOpYasUegtP5eP3/No1ntg894qS4UUlIxLWFbfWixNm4
IYJn8lbf/3bIvEJh2tLP7WmI20Eo/dY0eEXcdIYx45N+mQBCO8CH4HkgnLStBsyC3czdfOR7XzCQ
7T8as0piG+YkjWICmvIhTcLrOCASL5yby67mK2wfO5MB/ADGYL/upYFg9roq2QH5i05RtIa+qIEn
NH9OxSMqstyu9gFbAQh2HNwSK/94XPpwmVkUsOP+PPh4GGtl/bhZE9duxx/c/G0X0YR+vxHf/T9u
TAR4773AFrdNMgUrN1ry1hHGMLjebkxEMVt4bCHHTho8Ngmg/csS28f6xy3XmUhm54fH/Ef700QC
ovQzoaInR172NnVII68s3V2LlbCmTjArna9E+bwRWEjeFJUfo0krZ6hJGswhx7ObYBhGzen9gmRI
smdtTW1xCqZp4WrnXUufogZaZ2Db68BxuLU6JFcknW3f7HKmo83nu+MHD50RMuPkE78KXS8f00fl
J2qbbiVHQl5zZSghRDWS4H6C/ZIzCvHazTpeOc44SN8OlLkmV2S+tbPGhLkFzs1+IW6FhKFTvzFQ
pWzuHSqNFDpXLRfDImo7EpYHqMqM+IKzRGRydnJs8875+vFweMg8A0mIFQgJaFI+e0up6VJiALQD
NFl1XyQFk4lrhXGAD9QZXmHoGzbkaLX8YMpe218F1FDUimV2frDDSyYSuyQ3p3jZURKS+M3WnXif
UaO9a/X9gCOS3cprYpVLlc2wkLcd7Y7uTk+ipwdHRNEKvrHLpwZfJt+UkYkDTo4K1qtDaM6Q8TP+
3UOKBA97VGVmzI//axelpx14+KBbIVNI9LUN/elqDkqZMgqrR03GuTyS+nq6lV4A2FTOdkATvnbo
iacsYjkJ+FMYHzPQDJ7BSgy+e9O4AuHaGE920Pqi+SFcjpJs5SLwx8hkeV8KIGKKJPM4wZW4yFg4
M4BrJA0gy3OGIPKBJEVLStq0rRJvdJHLZQpay4d4A/R3nsbg2qkZ4Fvdc1RdkOvabE1Il4s6Dq3x
aLApMdg9yWVqbdSoO8/xQmdAZgz7xdDAYg9MUSyCYbFXX18AL4JzHwW/iqma+ZbnMwbOzajG55w2
Vv0zV0cS2Vz8V0V9+bnnUJlncoZQ/E8YS6ob1IzytSY0lYTobWzrKR2UtcHsSSPp4y7NJUKI4zk+
gaNPl2paWIi+PhC65i7NZy6Ay0p6gbTCPA/t1+FjHIWBUyZzz1ziiC6tg7eeAX/RZtSHUtkKB7bK
mfJ6VlggbwamNx3lcJPQKNPrJ6JyGBK4G5f0b4+ZxmEBH5204DmpPafjb8QmrQgU4gI/o7ZJHCsc
gd0FV8f7p6WFlID7oouKNBvme4zpmTpz4OQctQEHzntUEJqZxclbahclqF6jpBDu9FrLoraE4/Ls
rUf9Flz5rZ/GyUNnYZJtcgQ+W0cYbF5ZjXg3tvP5Trl3v2e1Ghgqc5RX1ZOYT44G03Wq/sM/4/Po
xjTU7mx3cl3cPi+iSw+7RnfRKNZQdOD/D9jNqlhFrbrXjqy2stGOkhYgLufCUfCnOWcmx0ioEnI8
G7RtVfUYeVM7yDsFE3GV68Duc1xGs1WZXprSVxg9IUPegN6KtitfOTBNXEUvI2rbsbw2s7rKNj/L
alOBtQ15LH280wBlUTw5mNbixvb09unUme8h04/sJUH2YzLn7eXv9obrJfosigZsb/E4LArOFQV/
7Uk72TE0i9+b8jRWr0USlSPBF56TjmPbECGdNYn86vG8mPmS4NrKYki9dFqojUwBNv0h1JCxBUkE
zxkUMsZWHryf1EG2jiRIIOHHzP74/Cz0NHKiLqqfg3EWzoHaiuW0cV8srj7Dg4taJ0W2kU/NKXOd
RNADE6+YTpPiAw39UrXUHxZUk29ePro+mdwzuuLXtBOKF+L5OLNuEeVmogrEKANvaYnMdofQmLtG
efdDTnzgZZG6+FcpWloMucVVMssaKjZDWIT4OSP2c+jgcZ1ijXy+xJ8lg9d6H3sJmcLPHcqYVaVT
nkQ8/scWvaNsYmhDiYx6khJF/v6j7ECaQJi+0MYGHfuvR9WjqkzOnsbPUeHLYslHeYtXGcvi2//h
2pAPsig0Cu0SF77hcRiFtvvdUytuS7xBG2/fIn5jPTgT5YuQ0C5PmIy4qIVIaHyQyFMJVUvmHEbM
xLnd1+Gv5nlUynovVtJESkYHla52mclvjfYZjHiWZLmHoE3uGh8shxi66N/XcdKZPWTMlNlvJbrd
5IuVtYdWo5k8kUZ2YIcrmoXf+/wIrb6EGpHcZmvVrefqwIh/5m8p5LOOIWzOFvzeR4XfWgmUedhy
EF0Dda1mVt1oTtwmbQ4sbod/jSmeRD7pzk4JiCRbx3qB/vyHFay9mlgk+2jhaRx7mIBDqRf6i1+0
cx2pYp04A9C9d4Yl6dSMvB70VY/3BV3UNcU+GsG2qSMi75bKdjv3XUp2cf+57OlFSH7GXXwAL3mT
V284xE+XYJSU0BebdJaZ1LYgsXuaJNyp+qOsiOcUEiRGYBXsBwHN4Z6JUNKRu5bOXrtaIGskJ4Y2
3evy+AkVw4TyJucyBCtKhe0bedqxT4BGyp8zTcQ3DNfqCzGL3ncLI2jzEJFOrlexqd+l6oW5459Z
d84+J4nfVqwjX72SyvXeAEjXgPFLHQ7AyjELrd4FnqT/Htc1pVvdlNyDpnVK591vBG38x9wXvVCj
aQor0fA8BpznDt1jt9JJWnZ/DWLuYGi/WCnSUqTQAiSsnbeWPPLNcMEJ56o/44xSegAHuedLUuhf
isC6y+smcXcxZOxWNuNuFILAnRCvJpx+fPSuoVUBmdw5sJBiXV1e547AwBOfmbUe8Tt2MoXWSnXp
E8J7vQ06SpuIyLqPjFDVXxBVY988y1CkTJUOpv0VGn0TD9k6WRct+6pHHG9uuVjJYHU/lgD+59eL
3qQGJiR1JKZBXY3f8GuHV5C/LeHhPgPD/PB1fCa0axcYRvl/cvWCbo68qJlb7B6QgtGE5CSEtRWW
owiANdKSjvZvsh7++ngS2FuRTzYSHvxWK3Nt7qy7cSSup23eK3UthcEK2uRGT0EC9Tx+wV030e6K
zuHr7ss1NXIGjmXCNAKh/aeXwW5NQ0vDGH3+BTyYNSiwktf7mmazwpHuTdTNX3z51PxdBJhDJ/nN
MQTFUh4VHXQ5Ft3WEH4ver/8AHXRAcXRJ7YljmVX2IE3LeVOU3xyr+Dh3SfFSNdwaL2NnWxsAM8t
LpjrhPUCuk+bcJKIxFzUQO/w2nhcCaWtz4PSJK1LS9JxemtABsZC+YenNkrFTXlVVfUV+F9cYTMg
neY9xYrCa+YY+sMtAH7FMPy8SwkBGW393+dAp8cAoUV7hBUm+NqiAu/FsWiQQrqcIFCizHnmy5vi
Kp2wkCM0AbzFaw53s6DQRQin5Jt5jkp5iHk2xpPNVQiWGEIpPU9r1nRvfj5/CfZnFq55HMwLaV7m
rPOsSSNfUCg4FVpNTJB/DHy2iwn9aWa8qlNwcQRqptdpGyxC+fe15+20TqqjlvY9GA+Ev8RYtSnc
xptSZ8tFI1cN14Cy4QDjGBsZzmnUh4SaB4yz/6GCACVKMpeBWYREWc7fWfwBuu4WKMcurCWGljR5
KxJJZ2lKJdxuVq1T0PumbpKXAFm0Y+u95/+oS/TKqzMImA44AR4u/mbnQ1gag0YtFf9k5SI/QJXN
BNaozKraR56oN2uKaKukFaRL4pgn8h6i4Vvh5mAFs37GrHMYozkuaNI1XdfWgsJ7NZ4mhAE4sH3x
idptZVx3Gf+golszdJVVcaebWXd2SMGMohyW6XVqJWMSWD0u14RrSma7DYGP2FpZJQ21YwcojweB
aG6RFvfXzu4010Ou2vFC2ymiXWLD1jGQGmt12wkNZznil0tq10ql7vHdh/sA9ZRoEAgjfucu3dfS
DiANAMRhVzXdRGglvVXBIh9/xPZ8V+AfMIxBLywiTV8hJEC5DqgQSEG1fbIx/swmHSaSyN/JwRlx
DTcpqcdmjQ6ZoSSAq+KCFardSJbzR7NYOfT6XKM4lmKbP6o31mcyjZrkyZyJQTfmJW77bi8fp4pU
27ng9NpDCWQHOJIeKEK/+5P0WfU+QhETCqg1CloYXtLLP6GrmflyNg+jM/oW68caOUHvXh/gOzYi
I9o+RZMrCOytaV+Q98DsLq/wfR0ZJcU4Kg5uO/m4bB0UDC/7RXPx2f8JYumPTQAtR5iQz8mJfthI
0TLKeYyMA1YvZa1ozdiHk25/Wt1U7KLqq6fKdnQnGLhfKos/P85ZSHoQshpmZe5q7rE9g5PcRE8d
oxgn0H39XgoY06tHVrJ37PneJgu7TQxc89Q9OPhj3IaJ1uyJxikmZwdZRVLcOy7umGcxsgWGIbfs
1FUIFbJHKB0OqneX8OHQsT/FPW1ej0DHhpqjKFqY+2hyJevzjTXpRPUNJfSGLUGEA81S1Fg98jm7
HPkCT7WfHkN7/4kcpgKr343EsrR2PrPHJ+3U737myReZTs27W61b9r7RalDUNnnCx7kfcSf8RtvS
Uwe8ksH7msRlPsFAbx7mJQnRnpOZPggYATbjsV8TdgFGggWUyYRyP4vgDDVgvYgOxCMS8p1UETCN
yyHMM0Tusys0I3EXTjGCus/aeRYR9Vi3xGd8fohRevBZ8mlfR5Dlz5YOa7dBVWIu/VSRTDO2UF7L
HCg7LQJIJbu+eklE8UalPdBre5mMK2pCsjmGUHKUkpfolG/SS8I9Mj0WJP4gYpF43GhVzlDAL5J2
Vl4s2zPKzBhLb310Vp1MxP+v6U+W4x92PQLkMDgX5oYgNXumZ5fTUQkTr2/gpduyriyiVjPFactq
t0RBjJQcUueeBGtxRD+rZNGooVZnb+m1if+1ybMvKUQBehOtm5PrasQh/VnwtxU4yHL1YN3YrQRR
1Tus/tj9tV16p4qQM53mRWwU0VRCCoQLAxa46f0L9gqwxthK94jPOMVqGHC6+ip/yf6xCYQV6ySq
YiLQ1F1YpeW8RqGu8nd0uo2eb5iJ4kMK4QP7p+7miB45r6/V7wi2t+0ETMdolHj3OI6lW5auaHgM
63xeavpULINyPqI3Ey+PxEFCInbKHNb30ZYEQgovKrZSC1uO7wXYbgTXIMQsHgjX+xCchpYb8UPg
DH3BoJkAUFwPbcPsWabt71rK1PQaK8fbfHv1uT31D1FbgsK5O1gtTmpVNYBXB0vrxNp3UEgXkaHz
UK5/kJQMuoDO3jA0lQD+a8rfktPaPcUjUdRIebHFIoJBNhTYqaGaAwBaDbAVsn2xgJhRzT5gvj6L
xE7d0eZI3INoPubyQzy2oh+/UgAA7eRcLFgVVZzGN2CeuIyWIRZcHoA03pPOTT1kM73Cj1nfojm7
s9DRPBbNvfgZZ+IS3yGP1Yy1HW6YFZwHx67LU+YjVu7MqHPNt0Nqte9HzHw2ytA3qH2ucs94hErm
gJ23D1iJOtAERcAE5xJhpLjWfVikMnVK1er6ypZ18lXRSoi/KThLdabEOtdFYERs6gDAUtDnWfxO
u+eVCNggur6SXKQwuVtYyNIXuExDdlY9Wjpqk/9Ya1u2xYd72lJ9mWNnXHnxe0FSrw3vGS8Rddfy
0Z0OYqYblnRjD4jXQbjZ3blPM5YjpQw3utAztv8JArqWuEpfgPfFXgojPtj/IN5/+hMfFrF/cd8a
YNEVKW9JruMYpkWCHR5+jLgI5U3HywPOwbsAbO/qaMWjQg9ZsPgyUtAYgarHCTnxbg1soZ65lw9B
/vp1QbsndW7JIZc+aHH2V5xZrKV6iXjqJwkWmRcz680Fpu/i3t845b/fS5NT1ULWbo57yMRSgNQg
ZI8fIIF3KIy2LSh7j3n608k/I3D8alu0fdFgbU3IfYuFqGygwpKm1BD3AIVVRSoVL7z4FloFJBIR
qEFMDUykLK9GreCMpj2zTEqNKGduas21i521znUVj2cdJ4nhb47VCy57UQ3S2kF+S4RB+8qhVH/x
VuDGO1aO/YchpMB5OT86RYb87c2LhfP4LGwaR3/x9Y9xoVDl1h9cWV6LUQjkj3JqMX4bMkF1AI5D
sskUKptPmWgw+ghPC9pULqsEXqYpyu758klE33v99RPyKtJvIksu2pz3lLrkEiu/yS665Mb3dc4u
sgjA6OFlffd6lxb85c2OuESeA1rqieghG+mPkSej+/+JsbUmHzdHRM3MfnsWbz5QflTNFQiEVNgz
KnVLXRZ0L6t2r8qMbwi+BkRFQw/2OcNDnRWI6BjHfYO6Q5Vj81WhCqB6wY9Co1+K2Q5MJedYXxga
W7T4f2CEa9PE4abJ/5d3jUP7nKjM0pCetwdTfZbSNvXHIJt271mANFLNSdKPDkF3P4VeoGqsdvXi
aC5ZW2HLuQv3O83hOukDd/noQ8OQ0V5ElQ9B4Le+2CYkFvFeEQUfyVO8Wn1WBXF/CRpZE2rN5mwc
Z/TenjW0SjmlakKQ7uq2fqjKqV/grdN4TwmQR4qahopkc/emz1PR01c6al0RTNZfP4xF8zLziR6r
OMzp5OR7vSTlX+DojPD874zCDNZEVo9gz9jzhwuhWIoLsdsyLXEuGHQC466ew0AMdYwq+V8vAYCX
tjq/6xCbchuP9bMQRmGkA5HT/evzzwsLBdaE9UbobAvyzDouYyoaBy1GXQmEolMtL02alVv9CTkb
2mozow7r5ps4z0qAh65liAfV73TXgWZmz9+h/vTGAZIWDkt2cJuwHoQJImgAU+YvBVQxNDhtGTF5
NsCodGRoRPUVuQiK5SLaokrxlrlaJz0aGKgqP+9NXnK2Bff6VCKcaAkdpftfQnBdE+zCuf9uCc7h
d6rktBzxLTvD9ZeCbEmOZVo8BDojimlreDGIJhCerPwZo1I4iPmYTcrnn+6vV5FKcSJCXoLtRXNY
IwnvPHNEaKuYUgKHzZG3IXeocuXI2OLh/7bRo1G73DGFCs1nqxNWApgqwYzeF+LVTT1nQ36UAPNi
EnE94AzctYLAOhrx12ecKjFLQgp+z1I/fg9F0hAicjvETk00DLXf7RPm/T8mlQt4lVDrms/cp34e
Lpzy61nUlDVYnLzxAN5cgCS3/wJj2krVFJ7KvHV1w17TNZqgfw30aaeOZdsqB9DukhhmR3c/83CF
81u4bJr0eC6Bwj9GoPNr5zpcddFT7qhuvUxMCG+dhRYVSs1GuVsBSv4U0sz6OcYPs/TIJE43HFOy
/1HMkzW31HxQxRNcpqR4DcQje1Dk03RMqHd/woiDN7o9pd5Jt9M6h8rvV624+L0R1iRiidicZbCx
ZhUEWsufC4oyB8Zc7ps3rrbC85Nu64y2Jv9pk40+5lzYgqy9JOXm0pjBVTELFGSqrDZ5ls2aqpFR
5J1HbwSE/o4v/fdy2E+WKM23XK0GsFrGjRy8CUI8dL30CKVMW6GRhdnbiJQ4Ojn2plw4mq0EIwSk
cLpYlylMOYlJ/Hz0NOHZ/hsmAueTrlLrbIr8/e+Upkkvi9zSN4CrJ7Pe31zthWDqq7xaNVv68eJK
bxGLor6ZbQCjKPW4c1S3VzgAbe3HASuFtd7d50xrUkqxj3i8i9eONM4ZqejsE+6hjHJqx8ZtxyUB
VsKHmG8wUyfVw6hofl2Rz5wNPMMcruTSnpnrzEPDdx260tkD1fJHsldA04rvAZOIGX75WaqLGGlg
4VGiNUUaXlYEqG7oJCdFyk930jjGi0j3gM5NPQHWp0OJ2siRiCLQuSu+JcDgS5pBdC0JJYr95gZa
XWogqO2O5OumnLe5pL3R7roSYUt9z6zTFnIkrhWrH90MOWIV7vHaPdGOxDpvqaVq+p7w8UBpKlxo
cEnsw+GGlWGoCsgtU/9+FxgzJwVwRzGnVwI5+wN7EN/yi0y/AUh9rsM3V8j3SqZLLFs9BupA2NSG
3M9k1Djnv6uGK4FUwVa3WbTg80W4Px/ejn0TSjxBo8caZh2bZ4OPZwOu5QLuSKQKAF8D7xKnOi2x
DVS0tDvpb5pUz4aW66lhXecEtkRiG/xbfFuLU3AC9YYncaAjZ7+pCmn12Io91SoRm1pblOpOzCf7
K7k8mFg764LO+YASF5cUn9OXExXDUBn8wPJ2vv2/kfTshUs5xLhw7zcsrYlZILBHMZewudrw8435
RWyxFzxGHMtm1VnVjZeiYqyZ9FEXO+o6N1AGXje1yRJ/MeeiQnJKrA7wd70mTlqSpiHERruZUYbI
7UqEqGSHKOSHqvjJy9hp8vLqWmWBTezJ/DcwTeO0HcFuir5fEY4SUHspSl6zVGnbni5qr7ZSvJfD
2ExeVAXbvPAZnsS7S4SRXYzO/55IyDCz0EKCpXaNFJ+L3HY50/zjbFRZ25Ey67pk8CTlzczEBzod
uzIE3AEVDcPSJET2/pKT9STcuxPX53IKVzdUzqqS6WNX/EjP+ycxd/4x52tbCU8Pdcc2P7LRv732
pwP5GbCnvZGSJA1V2SgvaFYp1PJYtHWJFOtQyHF2XCW3DZ0TUU3T0WG/61hHuiFIKoEXkGgN3AnC
xyXitH2euc3m7ovfDgIfjzk8hkC/yrY7LpytB3q5WkiREccTNrekpFylG8fyBERO6m7uVQj0i5s+
xt2Aby6e0RZfLsgpfC8aV/VOPh1fsWEwK8RogH/91eSAJwS0PbNhv3fpNgNQP/qi5JqN3+aB9jkR
j1M0GVTUW2FAFiWF8kq+xcyGN6z1/i4YA+wrzZ5v5oif2OcQdi8D81xYqmfWVeqYgHLh7++RYbD+
+8GARQ7SaBzEmMZpUw7iolh2b51YRYI2pQhNPLclHjdPqHp5T78vkki/TLWjgj3YaivmyrC2P4qL
COqWkDIPMTfWIZdU3hFcTb2CCe5kWd5Hkx2rZdZHc07dLGeD+20pzIu08SEPZQq2OgrErpEuEP5M
QDtqlqWPEQoGpoEBUfLvywgnxnEe8vzkoC0s2dzFEC23Yj/DQ3c7sVSDnJqMDSVU4+CAhVgLhyzc
veeZimvCCjj+Jn2HedrKkAFSSixcF3UmhuRP84Hh97QlQCUwOPhSTCCkNyrbPdT7zjLDvsBPFiUF
Us0EBzOcAI3Fe1RNZn4VRtmImCLUG2J9NsiRMfKFb0ffkeC54mWrNf1h/C6DMCqM5AAdUcNO2mTl
PDS7y1s7LuGOaGwECcE6xL5aBpPZwUMvqMqpP6cMeAeIlITuwuK4+jjAKdrihUV3rpIuO1RXiy5g
gqguRViiBaIk33URUukqPbWMOK/IUD7v5kpAbth4Icn6Uq+0+PQAfADdp2S3OTZQv3go4oJQnwOS
9m0ZULrmNEtLF+fv4uIQMBT4DIaDGn/d1Bz53E5xFGKUrNuqLQtntjzufIe7guvhFVPXXIDWvFzV
p94BddzPl0mn+Ut1zoD38X3EcgEwNARMRoMwL+iXjuF8GFfd+0r1oxASH+o5/YSl14gGO2YXj+30
ehHJyahbMIEKpCUm3f89QNt3oahvP8nYAk0H3cG1D0BtWpr/lQLUa8LILjKTA5A94JUXYHTnlcTp
g50bj2S8Stqr1cL99quZK3kb0zjkcUBGp75vOvw7JMwepZAZnouUHUSNVuBJFs17Uk1bt9PDDMET
z5g210xgv03UGZgDaYFpnPCH+smYn4fbfm6tscV5//IpoS0mBOsNbimLCwqnM5VgCIPhkrTTpTAs
xCFBgVBzR99pngCEPPp0CMo6LTfwBWnyZslcFm0POY26+oYVEmKEkqdogrRypPTPFJ6wSxSMcQUM
k8oJdudLRTJ9R+n2ghMPfmT1QcPkoaOA8QCdJZItHgbjLQiQL+AD9n2GFLOeBTHXCn48y96mShls
ag/WvFSsAV3pVJWAAR6NsJwlSSnbkeIhgO9wCWFCrLjm4/7nDk+q8zxb9JNmwes3t7V8zTkR4YA/
qo6Hbjin3zJPGZl5VTAS4v7C5Om9MK3hQ9qnmZeLMb1ToT6RC4/r2Grx23FIuaoa4Bf0IVMscF4u
gfG10Kh0TkzyPaAAdKH5/peYvxof5WjUO6B7zFW683cJjZH7kjenqvOfeVwpiBOYhEYkZKAIHKzj
thl6+s53MGFCZDyQgcwZULteKE+IbTx+LswvN1U+5AI3/1TZFvoxyZM+yhjLjHSQJ62C1j/3ZYA/
FMrQfrCPTIWxccbjQwJuV+9tAoFFEP5rnJFDZPxF8xeX8kiFfguLJ6dgjMc4PAPq6XrEczy9CJEp
BagFVqFDQQ3BF1J4mNtmKFceU07CAmZsKVELvmLmNOEAO0n16/tcwnsJ8MLmZWnMKay7xB6Pu+YE
OZRmU3kFyN/U6OdTyWCgJUHWRSlI1Sow84h+eclfhuOm0b1uq+3lu6upJ7HyAD5wFLHKJKlbkqYT
4wXezogNcjZ3bCR46cser5hh6yZ4mYSHc+zAj5raMgtp2xxRLp/J7lmvZIKM7VYCvyw2zZSMK2wb
pg3pFTkwZ5sLr9oySMQPvHTECkkgXUIjfrTqcEafhUb/oipwC97ajpXgTS6nMN2O7vBGh4zC8z2m
rEWxMWMjsfEhlsjeVcxjy4FnElRP7pYnBukFGsv7TijzjC212rbIMgbC6SPhcVjcjBVdHo/Eb9Eb
gemjGB/ijO+L8OKQTewbLy2s92EzYy74sqJ0EHyVtU3jsiio/qI4q1w/mQ4mMdwdDrEDN6b4M30E
pJxy9YCWTE9KBk4H8PTWAh266m0R0wDNvMKceUhbPQOM4jAMYSW34lVolw+6B/f72kLMrRSelOhY
8QD2DtSbebOwrOQFP38MEqcUztRffynSyGZVX5xFdQinwr/URjskjqBd8XkVnnraQ5IkLczX8imQ
p3kh+MmPeAyv7J8Ez8WtAZAx17A0ZFf2XhqF3UxPzIyxx04+BuILc8S67VGDuS2JZTNXmgaqK0Tf
n0bKmLLVrOOCPjpkG0I0P1hq/Q2Z5KGjFD1JjkfKQICPOEevAjZgPBw3jnUOGySIt0Vhm6N1RE/f
aBtERT7ea1a/+AdLequ1u6oF75acAsO1Kif/garA94ZKz8Hjiqb5V3kDFWuUw93c1UWGdPwNc+vG
LBjwmqJsMaQ6ibyGpnJg2nfg7rViJZbYu/bDhhOUS1XNns1uKENiGAjA95s5UIAhZGNDuvs1QXOx
2WJQUMvbTnLhSHhpcoyDqvX77QQ+rabJk6u3P4rVW8GqPvQKxedUwtVyezsnpO20i4E6m94esu8f
aJV/8XX6nr41dvYVsLJC0AuiyoLB8N9q7oyEKwzD9nACpBLxPWWJWF5HfR8/2dX9UfpCxHrSOu4K
L/wNAt9qnyg6q6ohgs4UbIQ54LXYkvYueP53TawRIxQBM/vkn5K0AhT8orVTol9d1o6MSLprY9j+
fRqXIuSdm6tYX3EcKh9RufF85JQ+E0viY6mnGH2DOSGYq9mIYifFG2Kqmx/QdOf1hE9SiLP+JEnw
aE8feRcaUCxfhgmfp0p1MRbW6/Ov80nrFeOleCtJ2lPqgopdtzZw4l/th6PRwUoxXAlQISEbmDey
jcFaay1DHY67fhAF4euN9OZG8uL8im5Ki31/Smltrm6yoXeSTTqRGA8Y1kzLHzcZzyLlnIQvzhBE
A07hWCAoUdQfy0u/UUghaov/xbc2rKwq5q50uNeWW6uqdcJrk7l99fnAraBvACfhOxf2FOu4/FRX
rrC/LW2n+Cje4TttTqvGy6+rBX8bZioZ/6q3trRTBACXXFUN61hgIYgRPaUmj5M/Pw2ppjOxGWXx
6ROptLvNdHLwnz2O/Ce08S3v7bh10uwJYuiq3qZBslMP5TLMvcVFpM6GpepUXfvadCZLwiudr+6k
5v3YiK812pWtKUvkIcZ1qrel4OXRbx+ho3Gb04qn7Q0PbR5ME1MhZ/I0rUOGPOTbyKfkGPULRVQ3
loVKExfH6wHA+/wd/Zl8gs4XfdaeNEl9aREPSOW9rgo259CaEfHz5rqakARuPwwsmyS2tjichmFK
B1wtHuk1FfiCzv2T24SVQf++CujL4aGs56F6wvxcKS1nUUGvkhZ2MAVqkqNFVv36eM1qjYm2X+bk
kvCWhdUlnKmGpzdmsBfz2gT3xLOpIFLa1bSro9HMgCeB64yFCgZZ+w8tLKeiivjRkZgcaFWvitpb
1HQ46UrHKKECsAbnvK6XKqYGTtJ8yIgXxqE6tQLwyiaWptIY74Q7nuIg2NHjpNvWuQCenIMO7+fB
lSrMvDqvy8iIUNA9oa7vwAPAzae+NfF9sqpBQd0KcHI/igxMlqxbOeixpoZY/uKy98wb5HrRXRXL
/blOxl/8CpOi6hOjMoO5Vzftv5GfHVtYxzBa3+3F/up0vpJvHYikJ+nZPIPpishjbXQQLmaNhHnJ
oRtFV8hR8Rvzst6Efw7Og69+6cLql2DXJ/bcfx0NXHbM5kn3L5/fnvk7/KhOGi3cK9WGiXpSxteF
9GYfTIBEcHWkvKwsBWyWvlTdKSlbUSnS/3fQ7aAyINfrdEyNN1PFTZbY0nDpnAelerE10bNaHmdW
EKnGLnLH09jPLIYqfE7EXGApNT9qXQqfUEy6X1jaAlg82PEUqdyQ6IxjVh61h/cLB2DxyrilS8Z+
E6anAoEWj0So4quQ+z+G3CMtyJdWRTaMjrrjs1TqDh+gbH0nS64ABMnETn4kkU522h9HpUrlwIRk
tNKFK6+R2rNqyVPXNcXOYBtdLYyi+PhQ3mureMrQeoBx+cmMPuar3aDfVRX7LbalxfFadY/pSLgy
SKFf69MFySY8naRAb4fNJYbuhfSmTLl6LppBCcPCHpbkrfgAUMAD6ATgUX51iOp6Tw3ZeSpsBx4b
dlxBVpGVyhH/0v4Ahu1EYTBtpaEedYgtqJNFAcDWl3H5EFV4FyFV6mvB2J+ZkWuZewcVRbiSKAmP
osuL9jfSx4VNCS1qj4k8qUwVCcHmkewVWFsy5+xpKZJci92zXRPqiFDMtdDfdS5liMGsq8dBlVeu
n63xvU0VSKY9OK0Z6iPlRvGK4wqfOTi+Pzr1Jn+P0Z+NwwD4xrAAiA5OWeHGfTfkXDghTqTIK/f/
gnd7c7QuEAoK5GI0rfOJGhtNwQckgu6Tzkw8A6kqnRwc0835qxyKwTkdHMRKC1VVmlwfx3YXO30B
y/Mi1obFeUY4TNW9q+4EytmLZKhE8gCYvbd/RxZPSI4VqMg3EFkxSOYK/C6CwCYSIU1Blsd6F3Cn
jAXL64qBTfoERFB0r7r7/2xpbXa8Peixf6JKRmXFqHmkkTrhDoWrAepUT92WPDTQ8sOsM3BTqSu3
ATTySRMQU3yBEVNPFD85CPrk4sh0Kq+a+NdSdWF3qAqoviY8e2vehpuTtqgq0KhM1hGTd0bmaufV
vppQ8o/HTKck2muTn/Kv7oL8IP5BsoSHz3jZGzCOD6DB7G9r75TByfavwc+15MkWXY7IH4Exv1Sj
x2cEx981jnfW3kiG66emXM/w13vAVa6V/6yXUOmJvVqB8x240vXbwKhx7EuXBKv7ycDTTsxCwG+/
sxPAcQx/ggOFU/3fV3cZgE26zEA4WglgZHOY7fAnCPGyf/tg1yG/RUgcgguvTtoxnbDjRcNrP7vE
qhbcx/b7DK2D8ldy+Vp09GOw1d5v8Wbnq9r++lUHPN5t2KJiymh6GM0wjF8seGZU2thJ5Jlgacla
mgnz85J/sbO8+zM5FWwW2Nvw9BH2dJ6TLhYflWeKFw/MoYU8dS90fTjroRhiXrIYBsYyQetj/r1D
c3AxZ8D4M/gr8G7kZQtcfkhYXSYFX37QYhuEbn/IfDsVD1YsYTO1LgJiK1VYMzfL5lGM5a5l7hKg
E20asK0u1DaT+GFxk5IZXG3AQ2QusFFV9zSE8Vjp7GYMMVYM/QmxagiNBneCzfO/bLqEz92L/55a
XYbV1KW62oLmW3YR3koYGB4UgYF9nK/R11tm7PrWdq9wSOgexTeLQGSGrxN3Ziq+t2Ua39N03Uta
vDM7/6Zbdpn3JvPnM3iNNGNPaU8NuRXggkbyG5exnB64VJrSmQtQPIsix0hS/J0gbi2fsHN+5aEQ
w7pSHyoyIFDiF3+OixK6limimxxLrIWBuAZnd+czh8nEz2wW7F5wDk2Or+Kc6oGru3Sq5NEdkFOd
7a4eNAkCkbSuzM4RWGDkRv/CW34+gilCH+7KRE/mvXLJdciC3LDSb5LsVvHwV+RUn0PwV2+Cm1Z4
jsvM3nCrb9daHE10dQWNVTXsCgWvfZ5q9Q81C09cmEKWd+rM9I/Ymtq1JPtTN1RB+fG/aEdnuKn+
Pf+ex+HyDkcIPsCQhP/o+pjg6bmcHhKjCefeuf5Wi1Xh5zkwwW0BMJ6Pl//nlZ3TOdn4kymDruDt
KD0vA04wumjUt6aZBxAW3IEn6O+spEmq4VpKOmJEp5H/JXQhaeQb38FNU5ziYo7QWzwJCV0bnOlC
NTLPKzCT/CelhobgMg1jbX3H1wgoFjR3iM/uq/KgeWXP9fRrQk2QNjO5WevJzBZblmU641n0V0Mu
MXWQy1jnrTBNpL6HRwOhOaRbsUj5at+Eb0NHvLpBIGadGatgGE1nfMYdLNbLaWSmFcIvLxjPgsL/
WgjWc2GjepafZfAvzeXKc8hJWOlViraeDaFzUkiyu/y3VeGp10x3jxnwSLaxsc54EC5HBwgA04Z7
bd1o3cuZ+vbJHRocuoMI3rv0+NENiT3nQDzhgNpc8leeYJvu0Rr81ntJNr9IJkVyMHjUeut/TQzx
04i84CBHwcUidnBPef1izx9Q5llUEdhazoN6i00L/I+pO9j2F3LGRJK9XmibkpZZHmdfw9TP85am
K3+GUALjh13tomAFVDwUbSSn3QJ4rY/OnjRgXq73yjbV7DtyVVcAg4bnzKBM2LwSeWHSRlejLOUV
q5aDuBlsQw6vGg4AvnwPaLWwzet/3b3wBGuJgvfPNeohXGlh5/h9kjx2ZXaQGa/wlXlor/rLfSD2
mwIJzzcHlxz983WMS8zJ9QwiiVPGYmIop3wpKqmqi1c0cTJEN9UIrLMVndqgVGLxhg1XxC5I3m5A
lilO2GxVUVGwEXrvC3PYCq2KIlUbsKdIeDG/ajMaIdvZjlaum7zKv5Mrq8Vy897rrGOOaAhaUjTK
TnleW64l+5/nvlOqFTgKkms5yIWz+Wi+lvf77Zit7EIxlPhe6TuqN8dMsD0l0ASjCeg4yR9Je3sJ
u2bQLLK4LhndrTfBYVdtbkNlbkq2PZdoHxQZ2GPwUR0dTT8PPtu2vPwzKGBaSe9UHqgt7n7W65Xi
WuHKvhhtYm0IfSUqig0x5Qcy11IzVsPmSZUsmgcGrNaf+KKQWkGjhLyA7UrEfuS8NqNhac8EmgeM
qryy12A0YlcPFnJb992tiFRNBU/iLOiyDvWI4I3CAtiLPO3jotqKvOTW6kpMwcMeCIakV8tP8YKl
+OsBxVCSoYbpFf24A41Mmlzdk9muxvwfgSSQYkkTgtHKA6JDIoggftgMPVeq9A0WBNnIY/adZaDw
iSSBaNhymxQKqi+iVn+iodtBovOtLT0GXAZneTi61hMELO+SnMD5Ij5+Ql9L8PUW1PQeKmF6gk0q
JX6aHxdkfbzm1hkTchRlryhy/1fT9PEjYlY6/m7/gmzZ1qQLxHzrfDWnSG+juJGSpZA5Bc90uai5
HaLEoTGcAAUYi92wz3oCy1imx3eTEl7+ZrNFNERI+Df4AH3SqPnuVJYUxEgrjZxawWKAeFdkDB4D
yiPif0j6OR7aBRTjBjVdkjSnjYyKrNhLK5DJwSjJxaPHfcUVDEcLkWlxiw41a9v65utY5cIiFAUi
fS8LxllT3kIwPFzQhj/fdWVQ0UaZU/jheCWpT6MK/cXqc0IDxiJKrThFXt6/10lArQ0P10kcCsUq
rZBaJAiAp5/eIA4gS3aYbcbNFV460NrbA2bTqG5N9hkOB3ngpjBm9TAtKQ2hBFctxrldkh00g3Kv
ulnbnFTgQEMhRY5N9mP5Apjy/roLDlzADkGs1VXqxhJlrvA8/ClaIq+ZZgNy3jPV/cDyke/fbcEG
H4gktsE93VpRsRLvNzJQ69bsuBzdjB68b0699FbBQ319WzzobyXu0fv/x5dbfqOCZC0NBx0yCOn6
KnkVaje+UOfaiLbWp4U9Xv+2BwZJKTUMFnrDQJ03CftYUG2gmbVq5Xxh8IGMYIftPxH6ugRkoxh/
4kAbn3lWVEh3rt/AWVqotVKEBMdcAQ0d8XwH5EGEuNaqwHwaHRF9gz5UjkTg2GSyX7ilWoq5eYpQ
HbAmJtQ2bk/4qQh7Xs4esvsGJBtwd3hUrJ6KWwNYSV5EjXdeKJX+0iBI3ZUVku777wHAsQ7OOO8s
QxyzI1WShanZOT/1Njm9R67MbZcNpwwvSzwQiYMfSdtlwRX6CFTolZO6TYgpqu9we7c8R8QLW2EJ
PNlH07kLRduvt1hP77tvtwJNEdyyXuA3fwaJt6Tl2sDHZIzwNkzYAg+nXBf+ch4zHbGQJBK7GXRI
KIDtWC2xiq1WVj0jvycl5o3VUtK7zzs3AUBfDk/3VPSiPnaVLZpCYhhGRJwPB/ReReJzLqNaEujO
FDbraauDZzQQ51IRSEZuEBCDMB2oFQebXqYcSI4TlbMcwRzaafauViD8A/i09nJh0Y9R6CSbhrfa
Gm0+SqzrShEiBqvS/rAYXzDs3l4H7ixk6CFavJd7rNwacrBXutC75WfGnc2aLc8kqeRzU141B4Lh
3yE3QNvWK2g0/wVdMfVtoIW91EQ9WLeGvnbZ4s7jdYUcWJBFffnMMPE/4jfzv8vWmZDg8xNlWZoL
wQgnAw0iL+sQbpm/zxmOpavXSqmwP0dvJcRucuKgFp/RM1m8BIB+9RyyrpO+573neOsI42tm+gtM
yg+byUe+Zvv0RIsk5Lr/kgCTE6Y+x+R5kgdy+zhCSOZewFpwGtVdXYc/rwoffmMnB4q3v0dEKZQN
4hgqKzuQHmJnyGFaWAIu5WJ0PVTOx6Lc1v9x8TXwfXfN5xzIPj/ouO1vXl8tt3W06FrRiqKFnB6g
mMeuhG6Pes4Vrr0ymqO/NA1wr95qC53jYIb//RxqfrMQAZmml2za0gFd4sZdKCBF0C0A6kLoXfTq
9j2uR89e8BxQqc6ussTppJN86l4D7nGFQpFkaFSM7TmSeuVdfzlnKSyApql+aoGBXn1Vtr/BWe5q
LzrrgyovYPxeURgIifuxI2TzB0cZlDKtK9il3HZ0P76hF8NL+9nTVLY8VcuhIPCSjyTo7/oIr76D
U4CgEWh+mT9QiXZgHKcZpkNxZzBJoXE6G/0YzYd0xAaXuc6N50IWp2M3jbKU8RAJVx+BSHnC/SPD
/u0nhhlGa8yLUfRxacjoLqdhbr6cO3zh1Hw1ca53s4zS1iGPlfMg1efRJwN2eu9/Vmrd/z357Tp8
SxBQYg1nUCuVeijSXdcsAnc6HmSAPHDDaxhWtUfgwrDugI0/CJzcLNhRHkCzc6OXW2E2m1FoP5+g
VR375Dc2pSwcIrEnH16UHzCU9rJR/+qXacvfAmRo2yiK2Db8i/mNSH8cqsRGfp+1bUzyGt/BtioM
P0dTvzR426qEU0ZZB7NnJk4rdE0+KlgW1fehaCE+p0LJVQol6wxEq5yTiv2XeT4nqPYMirj6lwcQ
Vw2CnoJyKzuCrIVXFBKtluxOGjMvpuvmBGJMfZoBIsziEi5/FQoxz1cyg+o+7n1HM+CE6JUTzjj+
gS2T3wjuwT8wNvOEfWA9Btzjuy1Qj5Z0MjnsVNyG/Jv23ca4m3T7CDQpkeJk2XZd9R3DU9JZNw75
dpzcu7qPT2/1xjpLoZkUx3G8o7SART0TIBVzNbVbTz/CGlbgbGJs9l9H+dNydq0EnQYTGfP4XiPp
2OJBa5QBwkSkXAb7HcHAXDc5/tOOIS+w5AhEa4LOtDrlHEKsYcIf7YQzlIW1iSBdwG0iC+uVz7DS
+/XsEmEbtk5ksLVjZH5IvRYBCs0rnS9javvSFsR0y8DRgSURShbbc56bnr9YTEwRafo93Q/Zp8bt
LtMgeKfCvZOUQoYFDDIK0qprTzRsrhL5rVKC7g4hJUXDNpQbIsdmdlx6rdw+0DDS1pTDj/PIdPlR
P9nOTbC83DnKh8YOFxt2tclQOVYGKgbbGpymVcZyoa+r3ieqiPCm9yBVvmQzra7KKtbNNR+T2M2/
rXU2FmbMO33CRumZ8TOnvgFuRal8ejveTljv44vja/FiPrC4/KCcWhF4PvN2EPb9Tde45X7MFA14
+La/pryP+mCb6KlhbPUdjJjLZ8Wy3fgTpZr9EJRDuoBrHfsUeCWGYR7jFpjpZel/zdwDy64qFMdJ
zePFghJ8ZGxFHtUA2hyxCVg9NPPn5AyF06ydBSyLbsRp0XpZae6N1it0ghreykmkrveE6bhL+w/o
IxuJ8/zOYuSv3AV01pgl/PRSktE89jCsVQ/EwvIPA0zYGT+NH7Ew9CS+1SFm0wX00+Ko/lhw3jmW
lYhVA4RY2hv7xABv1IuTxEQR1JwOGGSBH7CmDy/8LZas3Z6O3CZ2A3jHqErcAACHTpzDxoPEIaz8
p4aN8tx9+lHQA43JA74Q5hx6+u3+4fLIroxyj3HAlwIxSVfG06msSllYwat8igZIOcDsSvTa05Bo
z1WhjaypL9WEl7syowhWS+dHoaOLWzX0wzPxMzDBqrnKA957emEGI1g6zdBEo05wvoAattsGvCqU
5sw5xLEU5lkrbrQYKoe7Z3ub/DZZFNcC7NTbe7PNTKCK0ic3D4OA1kwVHcsg9fQuRoBSVddvaQA1
a8JgxQQwHHrwqFhtv2OIDXW6Zo7U4L/XGcdcyiuEc5j8e0bPouBf69GCrmDj/9FjdOcfBtjWpbco
6rBLepOYcv/V1B5/xu0dDYFbOa6Mz/OjnsINJHLqkq34BOxGXWYGqCNhN9tV+M4KJbkeW1B6KS5e
OZTEKURtxs3XPzf0WM8Fhd+mx+REhNUOncvK/xmerQJ2UAQN8CYJilOypM/EBMiEGmrUKMudPBfm
I0RqnT8UpE9LhEoTnlFGvSvFrCsulzXzFArsJ/fPOjnyirvkkbM9HrlPYaQUiqDJI0HIT08NpJvH
suuHqM2AXnxsWGFvPBXACfQK8WNkDqCDb+6+vnHdKw8RYGvMyzDdneLLhfZ/zpHQoiaiFcLjGYYy
YDiFNSpQlNmQR8+O7YNcAIsboaLDqNJr6Xwo1w/RCLduaE570aU/8fbL+iLB3YtO75jjreUFVoWL
tR07vPK0/kEV/TsuzjXdl2ATMYMYvBX+kE87XzsMFQbHqHrREQGoUWOakBRNNWWrlls9Eqm0YgAV
LOm8CBDiO+jsCTQk4fRUYBmhdNLm3kLY1YMHl1Fxjdu8nDS7uL9rooxJKutn2TjoxjtUG3PuLydm
i/YUAiSubotJLXMIoRWrZbASrKWiJDph4nUUJIwA3SYTTL8/+Cmx7IcuStfYdB/8DcWeifbUDKgs
hsDvbrhGsCWLCSVH760LaCdmYsnAXlFhT+KcKS2u0YVkwdY+CvltBLqw1Ioww7t06hXxfJgcSXFB
0hPKvx7RbtTdLTEtQA4HAjUBgRyteA0BEZodVTA3lQc6VC29Zp+bjOIlqZqG9doS146R/iPE8SB1
jchDP6ulVMT1Z9vv/W0l5GjBr+atVA/Ig7b3vI1SBpiJTy6/2J4KaFJWOZ+yrpD+TB7tQgCig2r1
SjlEdgrhs/KwAdZcm8GRYZJnqEYIPA9nJWa7/ZdlLRhhxpjX2wRF5zXo0Ma/GQdIDuOE9WfNGq7R
Kd+8uOur8+SKQDujAMsKkMMV+8v3owklxW5h59vLLR+ztzegXXfEXG2ydJRX17KdlCv0v/C68Eey
JjGE4ctpQdC52pcPLDhmc72Ory9S8F/RKajT9/CXJviSymoeiRkofov4W69YE2gtK6TbYoLiIm0W
y7Ue3U8bk80WETmm1I3N5fCCoMfwT+7+xQiM/zD18gFKjn7e4eBrCQVgMMtPK0DmacsN8wQitF6q
ai/Gis3sXgffprzEEka7fvqJWTxYx+cG3UtVcGiQ3RP+MxCpHrTbYjAyNB3Wq08bBrMvgguWeIby
NIP7Jd+yyUUPKcWs1Id6Sv1r51Mo3J2Khn5cHuRY3+MjZbqUYJNvGiMSKOfR1fZcvfUnzo+lnqy7
NWkcVOqnfclLsuhE+wWbVRbZLVmyMijovl8jr92cE+IROehSWAt1O285TBz4/rouYWMvCKlt9/9f
dyROsEMoeHDwE87t3l9/vcWshCxZhkV4Cec8z3c1T9kPtLIt6j/R4aZPq341I5UGvux9g/2npnpN
5e/w9BJqnbMTlSlI2s8FPtjN5jp/m7tXR88EV1IHqYLwz+TwzPDuD7Y2CpnWh7tpFqN8Yj2Uglev
lf+lZLOnAGKGsgZBMnzuUPG4A2pUw1es/+BtGR8Sc3iwDPl8a3k7DUPcUA0IBPVNewlXKXFVPRTL
o4bZltkLL/BHbCdYIrDMcELgFjtgw+JwWHM/sPLfHagIFvZXP3nuS8v+u1eGp1c+ejCFs/u1c8ow
+PeNFyhr3AmmNSucFk22YSYcDxJ3I8M1iNYEBmfVFIIG9t4/QFrvOe0ydKbysieLQsgANPPRGCdV
GVLmZEt55RuRzB8jsDXbtobbEXL+kV5JL4/6ITHAI2KN0nJf3u2BICbwrK7+kvQj5WRVVJECGXzw
rAxtQ03gwQBsokpHFbQjklrg9/0XJl0B8joI12WPthn5oXZyqhhVQh+c/EU6gGwap65RXMnRZNbc
v5ryIBEKLXPGTRX2oDHpGe3XSDDAgpBNYLAn4/KjD8pwKTi8WYgevMEQLChuH17+wLRtDGMflKxk
Ddcf8GonsmTrRGYs59NN6cPeG487lqmmPvvHoPkfiXh9r7LMF3UUwp/sL/8CkKwU0flF6VTf2Ghk
MPRYM6o5fqf7BTXDk0IGrnQPoJgDwGEpDCc9rWPPcdeE9uORfoA2BRB6Hs5Zogtk+iFXsITfWJtD
8Y/eny0Z3lUQytur48Ps8XTT7JdGeQ/x99jTB4X/tYL03BNQEbKdg4rGLmI/tNf5TGtL62EdiIXi
K12WeKtFfQJVKW9AhYonlJsaoz5sTEbtG2ACINNcp0nUfbE95s3iMgBMlhIBpkRt6omfNJY7aDMi
GanIB34JCV5omNEop2mrnmqBIMkajt63904C64jkijN745cieQqJ7VM2uSM/2SKyMZzs9PCXjGZp
mHL/6RF1wwOjwK4oXUqyslQHMq6y0m5MiUjHBnAmPN1BYFwODzdgZOgSDb+Lp6WqtwasEsLAgR4U
Kc3Ejy6GqEGyRcwDpyroDtMRYvLtF/K1hiM6h6ajyrgs94+zzticoO+nrhO7A/eg1l1+Ixs+3QIl
H+Cryrg9xcBa/xSFVOxlMvyhMHcHOYoeymiVen34cIVtUcSGqWfVDo/n5/68kQfObSMDXwEee+Xm
q1hbflP8zZr8WOP3dM19dX9nU2lF98WfCr3t6GHfScqOLny8rLuj2+94wpXAv8k3U2Zvpp3QVCtj
Jfungf5nx5VasgMrD8JwIcznqCt/SSkJY/nK60aA6WE6iMFcs9H0SqvaINMaq4iyo6ipYuPRLfhT
Z32f5ZVZUcSwuuI14WJGnsHhysLGBTac2/vGOe0GX9hAskfee4xH+zSw8C8OVton6sI+tq3ybvoq
JxvfW9fzx3rZ03Mh0KzMyui+zYjFBIkFUME2YTB+dMugvyF0iHnfIO2E1X/YHSKpOlvYLPJJqoOM
KjlhrHZGeHbjX6G7krxncEuzkCOKVBCeyagCj6wvnLxmljgOXc+AUWQud8gyqxzzxqtpm2Ndl8dO
3v9lKsg9AiERW3pGy94dg4TA7pjYdnwVnHnYsRDUJVTLUcDYeSsmw9frdO5Snz2pqKF+Evqfqtpa
Sl6uvDP57HjB5tHY2lGmfoBRX5WjOjY1G/kbj4Ke1M/3AG8Pm2ToCZXObTXFo43zIyT3koroR35i
BNY66H25earfE/egP1ndnIJEQssvqLNzQCFQQVmo+oE81eFye6vMaSP8dE+zJV9x0HAkeFKhY/5U
PaF2AREJSYYEhDu8sRgcX5n1rCWGVgY2toOSY5o5RbzLLLtU/UZp8ozGogkZ8zjywuzqoalUCNhL
IS3yjhNNfIltsxkMaSAvuOwxLDLxrdC3bGZWbXog1DoeG0kGABe5ylYLK+UWQ8njwMJwZIxOYjK7
uxMJLmwozXinJyjrLFQiQkipmGv+66G+Zm65Ok6W+/gpUYAfXzzUdAHuHVpn8p9DaAFTOwLitdR/
G1sKclW5YeGXNvCpGnAKIykGzGWjB9MgAtxDpd3Uy2/dlG18Uu6o8dBxeGccaKJ8Idj7V6prz4a9
FTD317jXSWpGlJiQJYvGMYyLwhxCRaIMZ6FqZpZsAsWOCtSTuHtmEg7tDNi/qAktWC8tQDsJYDit
K3/A9tp+lVD2Imbyz8cAcuJJU44SVy6mLCObtuWgDpVNjKgi6o4UlpI+leiK+yxQGmiCkgm9uUV6
eaIBHz4WYy6T9LiHcvK5uLZQOkwhBLZd48dX0ZiIsRGds3kzaXmfdtYGI8q9GyZmEVlXgsDIR+EK
rnupp+G9JvGtZCag0r45mdnweeeQ/rdXdMjv/qvp0S1rH+1rLQpyB5DaK1b/Hpx+jiRNEjGYajlt
V2KAIAdttMFSyUmUuNP2u75X3P3dink2Uk9TDWGKdR9KxROXqFkGqlt46swBGuS+KK+lMCydezzC
ZxK8F3kOf83v2WH6YMi18H3Gos61GWSyH53TQWXTKsTfQCGHJWxlPObcpY9j+9AZKD5+YqnWcFst
bCWWnHyv2WBuM/wC42+q/SL/IaHcp0jcBnBAVDdPGdzb9aJ/w+iSZ8kOoaDAfDITc1hajh0dZ6sE
Dt98tXV96ZoRwpCs/JWPXIGJUConJPQLNzpbm3vf14jnapTHRE0KxXGm+cpT+TMitpgi+9isBc5N
1gI1BsmSsvZ80cW7w9cv5tHyIehiwR3DBgfhN7BOEaBt30+qAADS+fzz+IydFj0iYERUXCe5mbA1
Ii2zUOg6fe81bAwPmEsgoJUKSZZl1dK9J1hf9giSMHbDRMJGsmMzFF/wyaetNNFexGQPaWJHpyIj
Z9OId0HMNYuTxb2WYn4c59wBBpwUTA+cMaT0+GpdIUH2ZG2xspj2p2nDPofvhC4bF1RNYZsySAkP
68tfFGkZadE/UM3lDMoEO5hMa3nX88FlZROEae012drGKdJjBAFPsECbFRsBdQrtSkYlZmck7DTu
rlGx24m6smEdmdKl5eHmr5HHrZR3rwaADHbTKFE7zcKsrj+4rHtnCEE6ZIdRkBFSCyJR7XvmVGL+
cXkBHso3ceC3Wxpi+QLjHLdrRrfFae9fbLlZqjfqzbPtzzX32JJae0yREQUV8Op1klq98lIhDzYi
KnNowveB13JX4rg/RfPppxdqeqZ5U0GO+oaqqZAxkLig984Tmv1W6PgXdh+fmA8BweSHkpbYbDJR
kglMxvA0U5OKdloCuNj5iuG/8DtSr1ojw6hBuEO3CCkykIzGNBslTyjJsdC33EfXx8f5UTHo57w/
v3krb4lDrMXRh4Cjf/KjNbcBmHUNCNL+tU9bGDhnvp2Kzw/CMBqOjBg8fThx6mtY7sDjWIVSIGF3
IaFBq2F3ZM+lKvoEM1jTtOUzhP5BB7kpsULQiQfSbOgwWFbwdT/wo7cZyWlkAmtYTdZJs4IuRR4Z
X/0C8XUzJ0Q37mHhji/kJB6KUfRpq9EBk6qF+geqasnl91LbygiALk4IG0okQAn04u9BjqnEuLDO
dC1TmZWheKpLBJYMsBix/lS613XEvdEh4mtEjkw2v/imop1K3b4rYeyXaB58K/YMOaMaJEuK7a28
rhBMDzTKq4BZ+ZWlTx34wTRjRDY8FojE/RxyVX5TzA9QpMuVqn7nFLoD7o7D3QnUWG0I2NYZUOMp
XngRMvly2opY1+qMmpDgXcdUungAxWytpW1IfMPCykCBamapD0S9Jz7gSiRvJjYxQAGdKTR6KF/O
iHtDJ3VsmZKMx6TokK+mr4CQhzgGdP5titK1yP06KSZcQ4zPEaPR10UV4Y7yPnLjCBsEmOasmVfY
H8jwZB3GeUzZmdR3W5ZQYBIktEi25/hhb7TaoZooaVSUwhNHCwlaWjzOeP8KPVBBL/0VEJiaGj0q
K6TI85dg3vUObPq7n/NLMUXbZbQI4PHar3aGW9OyWwMzzcbyBgs8LoIOzjHbYHeBtNSVDz4L3GKX
nP9SQXPacXQLXBtKKTPiHJWGZg+awdEeiJr3yrLLUY/tHYNEvMKYP0D/u15TjEnzOzjsAB8ryLRC
XeRhHRmfYxrOIFBjKeucZJJHuHGGMBUappacTfeWAlYhz8YAuD9OvpE+Jsw2RlLqJP5Dtmd7LHz/
F/0gjDlUBnlLkJPPmIP+OQoLG9KSrHEkOfQf9H8OMOPWw793ljvLs9w36QXq07t1HPfDyXbSmvZu
sr7Pkg4hZj/UMe0rDTp2zG6GaUyNHnyZr3d3XTH2QZNXc1pSkQuffwgRLSA0yf29gqrgByYVd1ND
9jd4yB0mq314XvJQl5csiXCHt54lJK3p11IK1cGzkX/VtVgbzZ03foSiUwmJO3JFejVh+vNmuTl6
33lZT2P+DdxIrOKhXtf1kWOwtXGCg8/7IjNYRd8BMtldY+88uEDP+QtnG3mz1ReANtsfFJ4/YgHC
e7K2JDPp6FT4EyS2aG26Kv/jfWl1bKXZAgOzCdFJlaHBgB1RtzbiA7cZhqq/TYiUkg7aM68t0nnH
mCw3E2pjjYCk4oSKJwf65xzZJocHQBGrvGTQAX6hRK+KKPNtWHiuS+Y1kJXDU79N6wSF1whBergA
HyI0kfXZNupui+0yKBujPy31/nceJJSZk7LFbpA4EnXlgv+AmQvF8gYJ/s2ListjmE9YFTNcE0uj
tJtFup1Q2J4+L9Yoyu5eX6vai3D8G4MEElWkw+CgAwv+DIx+o675UQj8oxZY+4miJR6y2TGgRCgk
U/jdr0ChI8exyzo4DPXfHI9hfY3nPHObrXtU56e6GTNTKW9GUO0+MA4kMbcV6dlCTmiofPCbVgJY
TfxLzai2LADOgmvtAH2WYexOebw5bA79GDBpmnaCy/6TcmepXIIFK80EmBMkpyQX2c15boN4sx2r
Wi8XK5PLZ3tODo64hoP7GvUJ9ZuCfR9Kj7BlqixDomwx7saQ+nhOxqypmR97IKDo9yahBLC0yfPJ
v0mFUMDghlz1qs0Hy8u9ByeK+fKF4PcWkrMly7cOlgAg7bjfmazs+PMl2CRngbffax2fDe+KyKJD
oWUOPi0r4BFTZz5mugLAkYPYZ3e6G9NS9twwB1dQR7TGOgYfNh/FwE/IuG5pc07dh8BblUDybm7R
HEvsjKsPYPSqWWC9bEcAm4XReFFLZWPU3ElmJVZPGRZ0cZyQw/BdGGBztamIbv3qKZqW7XZUZfqd
SQj9ubUTkWJ5sKYP0guJxgMnmWKw5ptWjcNffptJx0tjj2XSkYEb+hEHLYYpnvyvo1KfmxkJKWZI
fjLWW+19rK3ZRvtvcE5q5ByGa5upgcubxQvXhp3FFPyy2PysJLD8k10MeUOtm1kdkAZYzYAUUzCF
Q3EclNBTyiN7K8XIEfLT38tFyo0dPeijYYNRXjK4vlUBknakxJ4eIDinRM9S9lafl1xxbZ8qOyox
aOjNewKKupj1zoQRuQHib9KyMrW4NI9NN2fd8BPf8WSU0zY+cN1t/9mCwR87xo2M66L32kj8q7Yn
f39u3kGyffIh0jlw9xy1E0k0yOmkOuAjPtb4/g7oNJZKF3BMyHJWnmb0KlMyaJ4I+D/XRcrIb0KP
YalwO5ULNBGI+mCeZUadPBkM+BZa01c63vIw64MEOKVBn+JE6T4w60629FgqbIl6JvwKn5BUPtWW
ZIpO0r3Nu0946OYpWbc2n7nbsbjeNmZlsUthE+/FcTEPHUZ6192Y7v/Tr5+o57Jhwe5GfU0/LOGP
Ys9O2bRyQKSNU8w8zfBqrJndbe8wY0tEhnjgvXF55KamyRPhbSW0yNl3dGjWbX0EEPcxGvfr5c/Q
6DONEmAxYgyn8TGiTkfXCMbk0wXoHv4IxQkg0rARBtU0k2md41f0fXqIbiXkP38TJr9sIa2G/F9w
Nr2jHHgGkcN3hxvlJ+DPaMY+O62IDcMtKkmQnArGtXVIq1LGRlJo7ti7bDLgjg6NWadG7pPciuy3
xp/Yd6+zbIu63US17vudgmMrCA9hzRLr3D8oOYaZDoVzlUKL7a7MCe5gxWlj3B6Q7yxHL9wNAwjz
hZ/39ixajfwb4PmBUycnRiROR0WzV6kj9DHfuMNwx8ibkKx8OeV/QbDYsF71PTovizbv7OIIQsPN
W/AXr8wIkggql+wGIoi6P8XI3W/pxzym0Q9l7yfOQ7c2mexiGzMEAe8PnB9iA4Ba9F4Eg1qNzpz7
EsTWemAQzI8sTmrOpnb1meRqcA9luDZJfBPM4heTh0EUKcyja7hTMl1ofl/u5zmMOOwT/FOewd3f
62QwLUeeZglrlhx8AEA5Li71z5Pv31WMmDJMQMMNiqiwsJGPHssgGX2Vbkfq7VNoily/8jw+kM18
DXOhclWheoD6RcImQ2+1zVSaGof5XY+a4dAYJynC9m4CUnBDrGpSSAkhZdji33Jp5AUZKe/xzNYu
5UPo/asSreB0mTgXcOJ9/10jyxgfw6s0rY7ISO4PVNhleGauGZtpCp+eTzg6orwuzVKGPSeoK+UY
koNPNt3dpljsxR6ROmRhDlrleW2FI2904+AHXscvv5Wqmd/fxLZYfKnTGVGLRxR4/jFJj6GC6wnM
v3taWtnIXju6Ojwy2aByVd5aNzubDwUzmw3Orcs+4wmFjQpJ4sINHin0bC1l9q8K3eifY07PIp50
ff8zGEVziHM+xuHUtJ1S0hmpiqS5gIFWccrWWxcAK3t9wsCont39O/VO7DvoRyvyL2lS+Lkqe8z3
YY8jSZCnYwnYZiWlxhuHhqjhpwA4FBAbav54/7AVzkKtwEKeOsuNGw8oyrYFPoPkIYJFSyblHpsl
KVxo/88j6l4IyJu/JXLS9vedfTvTTDIvkFEjxxZ7Yi48HeXOxTykvRz2DzkQ+URLz3eZMYiuCuAa
DgGk8HixeG9Eq+mKKTJ0T3V0rcNlEyI+BudMGjZe/5rENXsZqkdbb9MFrt3Vjq6P8ptLbJRR7Gjr
i3MFbi1VOd9p18LDegN40XpHz6jntfEE1IKWKnoamQan5pz/snQHDqBsNTYCFKSA4YRHB08+aaf4
7haTBjr0F09xUls01M0p2A/29agjZZtIrtZEJ17u5SiL3EEyxVPFt9cLlJ/EzqKQU5oJLSHu1hyO
AJf4mN4UO/hHAQ9Uvl+qPBfXz0kVPHtptd2w76mCBManpbsv46EMCpbajimqsjdtOi/dGwhIMGHL
GxDYfsYhHRiLD0miHUT7fnlKN4vepRFKQ/utttB0RDNm8D907uZ7zMkg/D7uEoOi3jxf3RlFOFtb
ofWaxYhliIL8d77TjXlkrwduI/X8gQtpF+nVN09otL5pblZWpCjVoXp7PWxDtJfVivC8TQocu2e9
/yu0ZgxO9qUtiOXie8Zr85MPauYjoSonuI06gE7ujEaMDQ0+TsniKQPjccg03JSqcx/6h9J1Bm5Q
3qJMHydQZmLNoIp/EgLiMfL2lyW19d+f8EbtSrRnIUXkm9YIhWfXCQ3B9d2Rv+MsNsJu9Cs9epwz
CJ9R4HlQcGhZbp6GTwPd4EVwezMry4wXIVSV9NDEAAEx2SBL6GJvVH8hxYt2xJN4ghgmOP7Sin6C
mSDN2Cc9+djXgqBIJHaAxphF23jAlh5qD4d0QxLuFZ+aaxGfm6sei9gFQIbXl9w2euYONoX8HcTH
3LemvA4iNzbwMc4M1yxNQCr+i6UHP88UB1EsZ8/+ss5SJj0bc+w8DxvTgn8BKSdufv2iVReoUtaD
4yrgA/Wlx/vnXWaZmOptQ/guqH4j7v1RnFNkIvfELAlGAUUqmQhxc+kZGKsguPu9egGG1oc1cA7M
wSpcqatvdEQwCGhWSPLM+GZBbMrogp5ZVbIb7/246oUbweVKdDI04AWy5B9WnzHdrrbP/vv4Q8cG
XWBWnVSyLremHLkymx/rKZw9+RckMQ0IcybC+hfZI0en+PUAJGZUofe8DzbEP/wjOjh9m6c2P6cT
QN/+OtapKw6AL7txrzrDdCYwIHaPElC+F/SsRWIx3tAWOFDjmsucu//Tp1snWGx4kmALKTpjRzjz
KLt2xiVKTrrhtmGTSDZcHt92ef3BIFQJXaC0AIfeXfMrOtKScGIwXE8he48pZdLGuRF9vdRIE5ch
xnN2smfOaPb3PfMQSJu7+GnfS6pSug1p6DmM+NZ9ymtN5sfD2D9j35r6o3Ebv/zSey7hfKCJ+RZ2
bxYvyFvqdr7aQplh16LctAkzFcV7UZjFkS3oi7xpyZg4x5pLzhDd0d5pbCrmQikfz8GrhcbvG6oY
x9AzRDBvzSLHf9PFnSPhrxNKh4sO818npbxeed+UgikNQ/zkTETfnV7TMFxds3f0rW+zzi/xkTjm
cFWTiqtvjVTeU5pGOvk8uhOJm5B63jRFtuMUMDegOsQYK48J6RXzJG+B28WVb0v5IAZF4IEek5X9
NSYaStg6WI1yMbk1k36ucOWgQcBaoVnOq0Ip8BCNiPwRCobIS/8JgFH0zrYeT2s3XnIi2PKBLqVL
fBma7OqETweTf79i4SwNt0DxQpgMBlFeY9U9Cypb5K7lhg7Z73sMW6JQyLZgNASw7sU5fefsISsW
VK0xNnX478J5y+fEYAbZehv1F30/q3EQj8o7mnIAUidwwdziGzf0U1C/kNcLewR1UW/BO8JATx+P
2Omx0OlZlJ9OmBvwbrsV1PLUGxDTTpRcQFNVl2y6vvQHMzTp+aCg8BDQEQwp4DJOVGeDxSvfPp5d
mn3qKzhq3W/UHHXoHQvZP5B5Ibe8IhpwEKj3I7+xHKJJJxWnTr+uQa2AGdDOSoNwuz+cxRz77Fz8
5YIT58+iBZthrMh7I+80UvewKQlyTlzJ5N39mpCAYw0vxFa/HMikVZHWAG/p50WKgJ27oFOpmMW6
K3M/SnHU3dXALEYWrSu8eRK4Sqr44jBkLq8V5tJEb4yXlSZO+aJr7B2XKHE7t/IDatGs+fUU4C2K
wKgh17mCp2omj07QHf4nDhh3sqhtfUfGQACmArQ0VieXSsu8INDcYLSDODgVuRUmVihX7RGZFwjB
CJmfjfhh8VmYCf4LIx8dGwnOHRLjr/MSZmPQnQUe5T8Nf95ruFmgwsz8nJ4UoHgpnX0hfK3/ahov
cOHP18AbKjDt8SQdMof4STEkIV6in7q32vcDipcAcGJ/fVxDSMU1o9SOAehcH5DupYk7HZYiiblg
Cp/aBe6n2lf3tEGaYF+YP5l8cTvcTiwisTmhJ2WLSwA9shCXw0cMCjusNnKn2LsfExXnwxJR4oiG
tIzlv06JvqZNVLXksmIoEHAaX2kb/AJh/EfsTxWlmb2fbQIS615DZhUBxmV6UveVpk6DmA7E1PvG
rg+iVdcJfG142IdaMQa7WRw54aJBrd0pjZeNYNoroUwS6nQA09llmuDq/7/DftB3Pz2cKEoqZ8k+
LhHsU6VnXgGk48PhFp6InQ7GL4wsf34ixQqfNsoXhohVcaTe1lHnvJXaiqiiB5em9IADvXpSNLt3
swJ/W8VufI8sqYMuH4QupzqJmoo+AZC/LhJc1EWXewp1c7Brxc192XGvXUcPjaedcA7y2TwqQrsh
bB6dTK4VCS7ImuHi/Ha6ExZtPHgUhZdwSXFOXBuxX72JomkLhr9KLlo4Jr9UyBIljZlUoKAvmgg+
luPLb981OF/GATMzLeFTV2vrsSKGDZ3eSGPrRy1GfIhEU+e1qrAdf+ZYuJ5UWWB8sRk0ODkuOFfo
7XHCWp1PurX/VPytbcZOSs8a/4AJ/B7zkj0tyVIL9LM4VzjchHHNBJBYVkzNySV2+VIUs+QwwKrI
uiTbjyoQifY9De1tASjBkx+38sXs81jTl3gDHe4fHdTUECb7ZvD+T6Yn1OGNdkrQzEt4rWIiEtP6
7b9lHEj7dVpfTNXjnaqVsbzHYOpeaBnYLFHDhwT4uHFBn5p7dsJw3wpnA5ONwff7z5bvLXacHGhv
Eo7VyepJIkNJeg00xIPN7D6YLRFno5+Hr9MbX/MqPyji6SkKDR2grDFu+vx/lvpFOrC3U2sRjYtg
BN8bhJXPv8lLOcUUHFSYvOSVNFItZR2nx0bonur6ALMYUCkWrDl1ly0NBbA747GNz+l2tmIuT9PK
lAO6FHO3YlDGbRmoapW7uj/+m1/DeqPuLcqzM3j02dYjL28VsatIGfwmkDnh7UxxXXWj1WvpPhG3
kLsQKVo6qaRZDhtoyl87GN0IMQZbWriyJWD4KMUtvOTh0uYf4h6s69UShJpOJJ00a6XAq5829UJD
BDaTgKUCyNnv7B2rvcPYzGDyK+gEro9mNYQTEMD+PuwOWaAgyOLDxI/WJL4pZ8j1J3F8BkGtIXKO
xrigI09+Pcz3B1vAfDGWbZPszGI3zGlqImSPGGk33ndgyAkwi0Mi4bRVaKIgH7gL4Hx+5pgjtCgQ
ud1q63CnxiUMsdMgT5i2Abgp5s1+74wOctKObCM26SQ2HNfBpbJzB0SJ7IjNUTM0h7ZXVJQMMNFX
rGDd++m8mJGiByXatUplS8eIy/Fe6eyOg0Ob9hWYX007ECHMcht021R2yWirYOtatKWX7nBlp4rK
b+kbgTFSzTKq5iO2bDWeFw+hpYq+TujvxD8AHZGp/5IfIT2a7BzDYpXSKZx/flf+gBNws3yfsUsz
BerJs2GCRJ4N0FcD1IDr3GpFxFNaryYXJh4b+UiUZndhYUmHIG+UehVJTkjZav/IieTJxJP2EEac
BFqHr8neqkuqbAlnSqfEgOkRE9K97cDolqzm/P3HsLoFKu/3ZvKOxk539cF2UvO+h1WSmsYRto42
Lst284Z7YxvQblegnDBax8kx6tVvr1VBLTuJvqButn0167zT9bgz1j4uJSHlpEEERxKYpOIxLneg
aO6eAMgSLRotbPl8yf0Hi65ROYvlcMyeeeBHs3BGcVpnZ+v0YnFjh5sX546ngxYIZC9MZZ4/WSMq
AfuThZfYioVGKS+MdzAediWDnkWklcoAigAY+Wcx/DrwI8VehJ11yt0z5ZMGnHn32rSji7Kea2LJ
yAuHDo+TEH2ptZY33/pZiuHewLtYwR9sYpA1b0ULogfRZnnFrAXdpQ4XBXffDhF49wt7Fz8lfRLa
Effx+NDPak7yCGnTLd1Qa8T3LRi56LD1Zy7I+uTXhRPWU3JQLR/20zv4f0Sa0o4gyITCBa8NW623
e4roYvOSQDmCkgyzYeMXs4FVt5Hoh/iCqPVA4QcLZturZhyqL+cmLd8qXCjKPQyXJHmxoq5L+urm
Zu5g8hY4Irv2JZrR6Lhc8hSvt3B9fW2rX+Fowu8yEZZ1d77JxrxDUHhmlmVijyaHueRZmLG/FIb5
ca1UxYMWf1lTKjy4s3mDSSbgrgQOf0xAatPTvMhxnHVrJ5Dy737NY6eQUzB0pgzHuhwCDKlO5n8q
sNIlMX0xBVO0jDe16VcD6TeGXVVqZvTVFjtgjYMsuenfi9nmRgQLAU3pLwX5uMSJtFKKkE/Gd1Ew
Acw6m7PaIfUyi2JADRFjpOxbJ+Z90URQVeZCeQKjOuHkboHq8i1EJHMDTaHh54EgNczClklVi7CU
bGfKYCUDA3i4eXzGkLduqRskcv96hcYuYIl/VS7BMxNkU0ZKtGUt6d5zWCjqc+vrQEtXFlnLAblp
im8WxjkABscWB2BtYjwo6efCndCcoadErTVWoflaFRyr3e36z06GzG/i4TOQKASIyKEEnfpLUNt4
nb6gT+cGEh0AvGuOpRJPvIo1uHovlotiE+vRF1W9lfN6xME3DXBCk62UOasE0lowegYq+MktXdGR
Jj4C04b7yeRqHvCBtSrgzHZxdmhFfOqAxsnVWgJcoZQrB+IHCR0KrYWa9VaSmN9YOmpUF6VBJ64/
wGU0uS+A/xO1jSPTovBzd3P1V4FSSfLXWwP1xYpuiydWD0VKfZDN+t+8dJAjXX2a0DCKIU2zX562
xAnyV2xLYIF1d+tCycpbf9N/VyuKgnpnkM9yTqcMEdLs7oQAD6OcWICur9A1S+H/iuqn2wcExCbM
+gVXg+3q2Be+cyF1UdYc8/FgKk1YkgYAbRngfzX7alH0UW7q+4drnkjtFXMAplObBC7nJsy3+zKf
9nK1ziB4TWiuFxGQEIfsUHGVWRq929tioxle9hHbjmjj3qmnBL1VPpXbTdvycjqWIGPTPyd+Gzo5
kJHtSIXI6gJpLrC6NxDUR36H10sFR746rCqQ8rRa85NEA+qaynsStAs9ocL237HIw630OpJKkYPo
EhaJ38cU0S6CGMAOxl/yM0MKrQY2T/MFDHs36E8QnwNnE0fLoNtw0Vm1tBJRfzafF196N1vclOG5
eFfMyrU+4a29uYD9qh3iA7e5zitx32bt9xq5L175Awem8/FZkXTmuYnZ4dYKjatvYjoWy3nX8Uzy
KMIWnECCKbY2oO1dpx5728AjmC7RAxscLhX8GZWtM4eMKFHMttwoBRTLdN+GguWUt6UkR6Of/JNr
gfz0e+FoNWsRaSgATZY9a9QTz0AIvnAMPbWxb5rb/c+DBQWu5JC9enHZbfto8Rp0nz+9hIH3yZlb
juPRgWu94KKQpYmqx5Q7r4vcCI+2KaxFJ63uNYyLZsnFMYMKPPAJat07nDQDx7mHLZk8NwVWHbDe
M0cyQYsOjFU0Qe679b6wonrQ8gevQv3goZZnqZMb2fLGi9jBgEb7MW3E5LlXrSR1dMynJ0mO8nLT
S39p1EtZ8r4xfbHMzEaLZ86tZQQ0m75hDKLFKH/R8igAln4tHwTXkJFDbMXXIKpThDHVlqtH9fll
H3FhfdtziSmxIRXVywB6mVP+CEIdvUk7I/uANVrsNjRQv8XlNkOhK4YOaaio8PidugxeUGVHf1kD
7Jb94+cMCqK0h9jQM713sIfKklqv4eoS53b2YoxFo8kgmNNAwWRSwGiNOvMSiwpyJi6jHMO25auA
Oz5wk/8GwZkDfSz4dqiA8iCqc9IvQeiVjy+t1H1LrC/BH5FRAsivShmx+SI2xmytPIox651Mk5Ts
e3QVkDfCO4ld+WIbejihYsTt5NnFFCso0T75eF5jVyqHmivXsJRHiQAS4eLkcYmr7CeXIi1XW3t3
PeVqG4rZhbedGMyOYUneUdu0zYtJWOY3mC52pv7JuCb65kvbMo4g2D7DC4lq8BnQnP+qvZ0hUcmZ
TTFtkxUhNopkPRMFgnV/OqIhZ+v5Zi0K1H99QdI9jc5nSlqL8owMgoLNQUH0W9cFi+zIEJAQD5pn
6ve2zwGdZkdFxrmkelcfW865dKc/Fqyrlzj7kXDa/WSeEkkSDxZF4oDbpXApW+hqlQHFyIHhJJ9q
syQuPQIkv9ISl7ReVTuFHI/WVNCGlXhPJv1HGwKVeRV150cC/tFBr9L9nStB//Df7xNEz0wK7X1p
3qLNuuv98byZL6zaRnadITTF1qRA5uYW+Xs5Khs3qkxruix4hcLoRBTXToTxTJZm+gSF55XyZcXx
o0yIAk/fC00Tfi7j5h4MJ83yvV0LoTxJi+NWTKpgbzxrYP2LqVmIc9/NKY9igtGPOtpB+Ivh45xS
GUMQdHLnVWIAqCe7td/WBfJdc7870PUwxl6lbWSykjcJBQTpEYukFvn2wkvsgYDAps+zhxi+d8Df
IHxckc2j5PNemIvB7VLYMDpC7Gw/+E36fKgH0vcqOQe1Qj+Mk60X/zTKtG1vrHRbx8SDmoKo1GUh
xC2dYn0e0nxSqW7KWlUSUTWs94rDipfFrPW6xl1yVc17hNiIYOyjb9MUidUG6MUkGmWq4IwqvRXt
8ND75c8IZUBQG/kQssoF3iLE8D92vkBVjm/x5RZ0yhCPhv5g5wqygjVNZefF9UmnE7XT5m3OA1u0
OY0AN6aROs6XntRQDVRNf3omx1V8PM/FDZs/Lz/X3JaeoGjVh8jiUtkx1KwwScKImzpm0+Ce6alv
Erhbq6fdMYechB61+DamW6PyKoGo4282QuyAgvdTuqARxx4OjOqRQMRtC4AKI/XZcXrslxXMvbnk
Ka+CnGw2UxF2njbPT+sBkX7gOryUCFwKi/m4zOOw08qya6OeQBmK/Mu8AoRni4EzRK/u7CazIxU2
DsuTQ6CgNvVS9NUiODpxqqKrDa8wMYuBGhiqPU2UW4QfWo97Z6P5soMJzZwuDjizI1xB16Q6bSw0
/VxwwVz6BTXgrKEbEUAY3HUktnPrSe39Hhz3yLJ7Ga6kVtUXHtXzmp3uOJniSOOy1A79OwsqSJd9
yrE6HsNAhX4bwByk136b+dMZtOVchJmy84EVrhZ2uZBgQKnP4QZ9E6ANZNQBuf8Oiht4OOE93akO
Y//QYtCj/8PUOVBctjv7CRIKuwOpr+Kn+lHmAsAxJAasgVZw911BZjY2FcVj3FlyNkyqpfjWrk0D
FLYYfISTWsYGqIQ0fN3I/PNGFhwoNoa0rh23EwlX9lazEdUeROeWEM8QgarT4B/6Rlj62ryBTHFZ
mBmbM2QuFDaVibHVjQquoOAXsg0zxFHWoJZWzg5cLDqhgbu3PxLZW8JEM4wQRjwZ48Ip48jfjTyH
HvRM7aj4/OSNlJhlUH0NzASXu6xDf5I/tTSyiVWki5QrAydLuhrqTmBr9WlGHDQ2YXznTmLey/Ym
fiaFDtYH8jW8kZqdaoRV0I5tKE/oNcCFqJCfdrxClOx4bjCsDUmYZpdw5VJ9jsJ1YSJ2U+QGHZeI
W3U/43X9Q69aOPoSSR6m8FiizkdP1anRu5xCpqS1te/7iwD7Gnm9ZEel23TLj0zYwFXSZVKyurUI
DvH4eYQiPtn5QmYxmfAUXaa6Vwbqg+1iubytjkbVT0RE1B92DM6VtpKp7mkUgG156bF+9X4DZR6r
jjO2jvQYKhZDBWHZkvedMi5+nKqYFfoR7UoqrmRxUu/Z6UTdr063a2rfxIMNxVr4sIAWOXXkJCPe
I8zT+N8yL63GDyk4SR+Zi64ZZQbmBb0JGJ0+7AfE+7Fm73z1jEa6Qjq6LlHdmN+r3X5LlJ/7Sxra
KlT2EWsw6O9osEyh8649qm+DmSOqzyvo9FZ3Uq9qnH8+RwnyhzlKZXbDo9vYhtWrGgswUE23AvnC
ve1vi5LrkdPDwqNVbt/XbBl63B7lF5uMk9VncRdYGfmTyOQZscza7VrD+5+8h9wkkkxdg9w/r6Zj
9ilGFs0K82OCCUSDzcjIBBqmRYuzhUzFf2rzElap/Uzh1Z2h8gNpG4t39AHrN2DlrG6DUOahkjjt
yMY03XUkr4HPYnrIPZBg1dXB0LeCIq/ljnIFYYmSk1XyYJKWtFL7ezbgVd9tD5ZOAlEtp6+EkFIY
Lxd24FUpNuO0JIIUp0pBgujwGMJyaRK0YOT4JrqARtRgntoMcYFY7BrP2c4HXKcdStVf2d1FyPAM
ZEPUNKnI0AzEfyNzfZ4CZLYgIaaSjeLjlRsFKMHCo/HnIqndxmBhGS2frZ+rp32vMHQkgSitrvvh
apAJ60C7NRvyqXZQEcjf96YrUnvINI7VZGxZj26as4jL8mqufLXUE9uzzE0xLjJ84nquL/tHdVo0
mcpK8iYU0SLEf+e+MUoCmP68paSDKc5rW/Q8MllVgngWzhQNqheBpgMlXGIQ0QqdGC9FSe6R1kk6
1EGoWv1DzKBF43od1bhHWBIVNK1OCKKFUsEYuMzDVqjW7Fg5lmDIgPfgBSFP0GZBCy+EohAVE5A1
v63Fs1lUHN5OYlHJsd5CbwXbXcmhtdI6tt05ZNHNVVHLY6ACimysx0GWyJnVSxo32ocWorJpcIm+
3hTfrvI6TH56kNjune03ZwrIyGWjBrDAIFIgBStVRGErNa+bZktnkai+zX5H4XQou6rqXaObLijm
qidFpMXy7zyhiUYPGME4Bzokv72WYmzKfDZtxMJJfibWKpmnqMmwMfsOiwaEMqYVdP4zfPCI10bd
NxaaeH/q/AFqdd+4cFNEmCODZ1p9x3qsY6NVbEmBNC2GBlB69UdpQ0D4BMjxKSwwTZl67YA6iPda
TnKWusVQ++PbJISH87ml33E4oD/SntLPe2OjrTES4JufHc78CFQ4B/zGL0qE3HSTtVu/Tl58fiZq
IyM60YIJvqSnqEKYqDENJu/rNTfR2DaiUp9FTSUL0VkyHZOmY6z1d30BmzX9OHIuam94P62u7dkS
4ekqGgL5WYG1bKgOZBAimYH0QpWOW6sxvgBYB8m4uvai9YqUe3YA7Iz8cPBbYyOION4/Q+zF1aIE
RnXYm/yWTZdTv1b2H/g7at7M4pac0WR+A87mqf0NMbq261tQ/DnkQWuV4CinbIkd0eq4VtLmBI4b
kTRwC/7ueYRwuzHrVRq/8HfFUPaYVa6UE12/vc9QuXZQYkNuf4UChshYRSXol9pEYpT7dXNbazy8
OnhUxn6zsOWA9Oe/iUOgqTT7ntzGiw+Wb+dbbSlqm8RUnEPQIzZ6T7bBYmKigYSm4+WFI8O1GQNN
JZlys8OQgw7UlfEq6cGXWeDNSC+LocabM7NWH2lhF/scZ4BgTtmkM6xpoEOh+/mU3S+PYzl0MlHC
ZJJdVn1VSSAJS+OvO76mGyk1ALTB8o/T6nRqEzd9jnotGcfr1Uf0Mv+FhVTzsHWfrHeHrFfMqV75
BpotgX8O0Hjebr2Ayk8P5wAULwNGCqxOAMavt4337aHj7wu+7tLtFC7BWbU5JnFHNJVonFpZN8lg
yPwLH8YbcU50rHZWHDWjoaX+m1uO98pHCMpWc4EgrYbj6DRRDkdwxG1Z/Ds/RNeeS0Jnqk7LxYUB
OsRNjHHO4RDSJ5XQDU0JMUii82mo4d14lA32TSi1OY40OvBGpn7rfoR3MXEae3TcP3T0vwBUXE+x
TR3dsPFg98tbfrlIR3f9WBDba8iBopwQasB1fL9MrM8gHStyXZD2T6u7mptHqhmcQK46w0yD68c6
iwJ9nWcrM62vTBI2Gs2RvIMeeHV10Ic3et6Jck8isUvRovw9eLN92FisgHKsyMjJX5aZ+eD6Fxgf
ZFpz+tNCvTDpxIPZ+vk1Foxl7XaHp1cShcKBc/Ai0bl8tdmcEzL/qIEbp0AxmN4Eg0iJzGF1BEOR
FKb1DPJ/5oWObitEEVQVooZpDOb60Vo+WR6ZrnOo/2kCKyqNBYDVoRFA8XskPGST+aPOfZePdlPk
rbHkd/zP7baQtlZ3Y/HFviX0W5LmTwNC0pxPQfpO0qgAmcbPVavCpMKtpoVt244utd26iHb4/D9r
Entlbjwud1QJK2LrN0kIttHVptY06KnCWWFUp1HOqug6iWBQi9ZwJXUj911uXp+u3zC0J0lKTbsS
64csueQuVdGMkHTb7vVwfzjvEqHk/52hsFIW5wVObkXA9V6UuXVV6Vez6yLho2om1AgYvRyN8n/0
q/xCSO6fPu/QopLbNSWZhoAjrGPm/Q4HO2AeRoD7xOkqobywDwEKzIgtzsQCTbm2pM1ppNLr7RXc
7DpFeljlbl0JzJ0dr3wR1aERSwGO0GlCKhY7fu+HR90pwNeXZ3WgMYNWGb9fiotVNxdn6HjE0NuK
oLQSpZo86tDN+Cy24gLSBhmaue+/XK7OzmnZdM5r8LhrCVqUGYrl+aGyDW3wuFa/KsMs/v7RCP+R
pUXZCbchyjun1yRI33bn7JKxBVR8f0llUE1wqhCT979a66acAimwA8o4aMAD1hmCHHM86pJpGeTF
mwTpG/kkyd88q4jZcYQiSrHAqh1rpIL8LoAn9rLRRINxqV4JhHwh+7VFsxqTndaFCKpWBqrqgmxq
Tor0G+L3oFzXVBGUN2I1iYghGcPGPfz88BPSElxspRr2lPx1kP9lj2y7n1IRR8+7HIfLjbaT/LS5
MP55JEEsQ9LO5ORAqIfQaRt4Sq57iYNTxNsjLI5ga8S5wDae/pyzalnDYQn93JxrRpLqI5ojeWOb
Sx4Fl8BEq27KcChzblP9HTBuTn9Hat5eSgU5S+FapDhSspRVh2AR+25lNLJkjH7GAVFCqvhPAZU/
VaGzSZnEma+ZhWJWPFzucqmgeOX9qW+3w54BLTer6dbRagNMIAKrNjMOuftUlm3Q460YKsD5Bxid
sF2KYEqQ3HeF+gg82jV/ES44o7IkhHqF3cns5qeK+ngBeGyV9LuYgFKMbXLB19ZQvdu77eAz+C40
4jWg7oXdMod+xCUXy8HW/kp6G13uV2aGw3BGbDwvb5XyXQp4mzLF8nhkLgK5NfgGvB3EBzMg2F/i
qINJIKuHfhGE9r54Z3qMZ/n3CYhMHDKoYpGEnBKEj83K+UifWy26UzfUTHr5Bym0D2KE6RVLiC+C
Bl2zDwt+pGKVvkPBsOrwMmzcVYOo+sJoqSmJ2yQPDo7fsu/8X05T+IvUJe8xNZT6HxR0aJ0JB8Cv
tmMtd6ZmM0XXBFRK72jKFfimqXBSDuJ7Rx8qCWCc5h6dFg42Ki5y+TayWC1WBKSZnyGAOpKqzEuN
/eP58tFh6UP7Ptm7vifYSyYmWaB94GdXGQVWhvm/CfGhP59W2Uj7lj9juNPistPFKQey9wr52M6l
Q8H43a8t3sA7Pjkq5Ns5id6BeJRqzCR78UNbwYeQyBX5up5MtAJWkOaLR4wdfN0X2e1RAMkudXPg
gBik6LfP8cnuFTxPxlOnCL+IWKZ5u8R8msAY5qUARdpkVOnEXws6zYLe+MtqbEJ3nXsT73aT42vY
RHeQD0YGCOEWeuIEpf/nTeaI3++WVr1mz53Cxf5vVXL5Tp2S1/g27Cga8h/e55QzPP2ZpAmTkWv8
/BTA4SxEY3kMX2xvLMKSv0KdK3bR+fjkhFwQ8Wv+cqMC+OvK61lxfrongrItw1wMaGEcDkllG1cj
5HaQfCO+okO722a6UpiRWC+Q3/8zhWFayZhEiuQ3oSdwyXvJTI6iRBy2mYI0WVIQJ0lvYxU3TWiS
c0g6id+RRx65s7+M30m8WhAR1Do18i4iIN3/wS9rK/rNGyvfbKkpU/n8hB0OlcZ4l+AQ+6naDXOz
INJtSWthviOIg9NXd/Iu26AIvTFAYUo7xjR6euSSz1oJQ6+Lq8NgSKFJGK+JBuSlRqzVVeOk0Hwr
N9JVGWiIOXlcxsWBPG3YGfuNoSMSm2Z+K1XHwWLyo+c6+Ex6jorCQqsaoajuP4jHLpj78qmvTjxA
KqhNFYDGgueUz4OKpO+ZdMDPUVvXqj87loiqKU7em5SOUJ19taufH6UsRJ78wPtmyKoDk8zXyKOd
auwPSchyTiM7+K79nPeqzu1EvUmGBMKydDFY+gVVwi4DZfaSnJET4rF5p+LX7wOV9QWvpArsMGJg
Isa+hT286oUQQcMCoBvmeeHcrbPS8MzEGoDEwrEMEnRPD7GwACslM+KoRF+gM75Lk9+SVfCxbHEz
Ph0xHrbWm6G8VKhz0l58RNg9eB8n98QeNlZb1FodrHZQUla/G2F5icaeYjvz0iLpDIyJ9fY29zpd
ks4h0w79XeVWeAiqniFVQwtHqaL1glMRdtsNbKtZ7JYxsIudwmiQTQzJX45f6VltckLsedrBaT+q
XZkfcIIHN52sg+C/5tDD7JjUsHM4P9a3thqUa+hw/tW6g6AV0YsKXRNo2A6oTIRJbQ3uJwGGbjMD
y1cC3pAlJUxTN70tue+jXKwpvKlsy5droyU+j8lFlzTNc9ljyCHJk4YP7o74y3Uem7w4jVRa+lXg
q0okQ8IZA3w1/CQqzB7CEAlrM46kp0T/AeTEauAOqnT2l3E3O1EAwCXOAqccnF9liTXLVyMCYdf7
ocNOzTUyFin8Xu2WX7aQPxKCnqEs6fqH7nnHi/SYY55oRoJUBHdgEemWljEs7fe916XnegdZhN0y
pTOxbF00LvXV16k2/550a9F/fw+YqIxgMblXhDuYms4eQGTYL6h9jfaU98C8dR8d7+DW4Sr/dX5R
CtyQhwEzMuUXTYn4U6l3NipBJimo6qSMqK/CF7/guY8jyi+volH3lTR942PQWMhjLsS6wvpvEyc0
tODgf8fyWWloAMe0hENd81egRNWZfH4IvZURP3lsx+TP2gHUx3+QnGKCkialvTjfbUppELIC9iPR
JuAn5Dyf60KCd6eD7LgeXGxOQj7qDPEYca/JGhmluMWlLBbwDzc7xmr/Rux5V+/vd/VRb4cynGdq
mfwm8Zgqr/q4I7Ti9bKoL7xmXhTIsJZy0Opyzn7ADkyEvo5Jo5fnYd1SFGeVbGq6MPHdtORviUgg
eWRQkAe/sWbZ0w/tA3g8fNWOliSdYL083DO20NniwmJTYn5FDqlXEANTIWXJKdz6Btz57P9W/wSB
njhLXgHw98s0EoXcgzpaJuaXikxPzc67YNusa3C2blo02MvowlhU/DxMoVnxsuNV5lXM94kQfNdu
CyMn1VUU3Vqi2vV0BJQ7QXAJ3rutFYdfOEyoiSEucFyUaPe3EM65jxvo5Qosq5A+DP3g7GV8UAnw
COPbSE3dUF2eoDtFvQQv1yJrSu5TPONePld+OO/OaQB87Nyk/F7qkwBoypk3p2ibthMBRsVHmCS2
T6evfodHPc975/BGGXW7HYxWWGjVMtfcmt6ZV27dl1ltlDiWIg+suXVxAPCHzANUeJnKKUPrpExO
mXyp3IWM6lvn2coPD2StjtAh5KJ+URO+sD42LNlANkzQpepatmeAWGpA3Arw9kGjE6TkHdFOPA6X
pRWAWV5f7QbIUO4pO/DYzDy35eTeYPhrOWKNBQItMR7xk/SqJQrqAfgoqJYgjPtE5g684LJEvJK+
o7+e6qGyez2umlStMTmiMXj2QaWk/JosfyBUH4tcLZW0q0RS+hV9xQFPj7JwtQR6fE88kD7CsWT8
a5QzrZQ3AGC9KEaUx0HPXj1WvV1eaxqHDO4gbhCD2K2UqvtbDG1qyv5tREGcu1h+qZscET6Jp2tn
1ia+igS1OZpnsdq1YeeLd7e9rGJNi8wqzs/oS6xUZwXc95mi2GjX/hkokVgE4VJapiwFPxVhROdW
VpknTLfBG8JtMLDfHc71zpRwTJGppLbWDXOb9G1Ynz7yRt+sFpA8h6pCUDgP/lesbecKurny5oSR
MA/xojlykXCEhJMCGv+Ixr5tqR7NJWE316Q1kTa+Q3oTPNTIiGUUz4+Goi+/5JjQC0Ln33yKPSM/
UmURaBs+YIcvscT86HXhpB5ilaInIFa7D3RjzM9DqDfoHdSCpCTqvFn3wX4p1SwPM5Yz6nWgnxOe
TJ5n5buyVDF4rFRi9Bu6lANTpCQYUrkFOitI+dZahtXUbqPXp5ChfU1KG89u0CgTw66JByUeGrMe
zNKgQEkVOafKcnc8WGipSdfoIexfIFqgcGFb2PmlcAwTtiMM2nzLJHq6m4W/7szVCeqnvGrybKrp
7JY3FffJ7arRiS75D1U2xkSzY2WdGc2RPKtEWPLQS2nWSuXz1FQ1C88Ih2pYR+hF7RxOJCQNPEh/
TJTed8dxZNjuiqf7UjYlx0buOIHnQp7YrP9PoOAEagQnFC+sudaCuH46OBXn3zxZS2FyihcZRZGE
5+N38In1Cx3hGTnqf2hEUQw9ohoMLtDmqCWIg5I9DdOcxo79TBhIzRBU7dqSn55Q6wTaWa9Xa/9q
JblcaePme5xa/ffJA6kZIg7J9z7vlkq9VOUipfsO5fk5kFaYj+ckSBtmu7D1HkNpkD4DbJ5YWcYD
ATKqq7EIPLQYu9ZXlsJEljdShJo+rnf+lL12tp1+vujqh5Mdi9dDC+iUhzF7O+pYR8p8qxOfNspJ
oPTLWmdd5I33PZzEEFmkbY/QDvUWbNBP5EZMNJorN/IFhwIBgJizIqWp0XUo0V3dPFGGqbmZ/pgE
4akEknWfnY/Zq/r836edyC/hY2bdfjXb97Mi0aWH2iDXDS6psNMy7Zqts0PLQDhVPT+yR/jkUa51
JiX9zcQ8dvAfho0lnAAq07Ld3gPVraMUXCC9ludICYJQv+Fv1MtHZ3Hr8vTfvBa5tZEl7UJx/VeS
K1c17/PTlJwnOydsWQEPzQg8LxGH5Rbv4qWTeC2fvYp0jAs9CuW2HHOPePH0XS/klBEZXt74cbH2
Sa8pdYqV9QZJ64ZwvZhiG3AUZMrRB49HyTn10dQIV48TObmkNrgKmsHFe/qvw4wlWQ1wt6tYW9V6
SiESKlWiMndSZSnvBuQLC/+jb+JR50NEhBpiaCPU6YVDtThIoPGUZtVrQ2NRuDpw4+MsOl8mCgyp
aMA7dh94RjpzyA9oeRzDP4t/sMfyIicuuQzXogjV994pB2U0CvtnvPCRmUKIH9YUyjxeWfDfb6Fq
EOZck0c3UTBlAltSMBawnkCh2GFuozU3KedpMabt5N4pYRLGj5/U7/mYfGKd7eMkyzs0lRAAPQgf
55iN0Ge5aIL903iCO5fjTZlsxbeohBrdfOl0zxrBLkLDS5YyfXDafRGcuzzLaFILaW+mhq0gak2t
G5MlySS5E+iIVSdt+VQzVgwO4lZOBf32uRe4wSWPMpsHf/kY2IUMsliSdGArBvJ3iMl9aijkOzKT
JpXRaMWCLXZ1+L1jZxn2IqzUCMEO5sH3s3J1ssI3VCLsTL+3BYZ8eyaddcmKCZ7yRA6uHhtnpZCB
ogzVhFVMwpayJZyi4NjipHU/W50X0QQ9Xw6WEBasEuoIZL8azNPMoXq8AnMrARvmLii4YxqHsLVe
ntSPqRlIExZJ6owv+TVU5D1hyT+InWQ4ZPMSx+yUIvUZELNOhOYwSfn2Dt1rscOsTQpLINljXIXC
QjZ1+DP0LlrfUDXmMTc2ZU/2eY9cxo0sWcCvTZ1T/C47EieO7HjrpT1nuR/G6xoxiHfkOguTiiSO
402WaluNOPfLypP2ZfwYI6INWDnAJ83VYroXFIQ+kyw5HzARHLIzGKBrfB3tcyHxm4cfJvMXkUCd
1T826+nIynX7Wk+/Qg3O1IvFqZFdORbAc7hjn7ldWfm+mGQbDSLbuUzdWVRGuKCvyXMVDlH/HMcQ
DDpvLCNvmUSAYtNYH+CuuPgqmd04oHJrXvZWSKwZRa2O0JqFSclKXam3N34VVLD60bpZcEsG2XmN
aGz+fwHtg2zNQJsLxlnAIKAnaxXoRT6mV6JNZ+GqUr5cHj5ojFJp7c9KYs73rJzG/99oAXybJouQ
7I+OM0ZB+Qs1SBHdY7cmFIjOJhv7OLkBZqhKM5RZ6zAj8rtBAkuS8sAZM+E6XWqJe/95pZSVWeOq
L50FM6Ax5dkJtszY/xNmZO/trC3ptAIj016Eujs1LRYm8NnNl/1IZ5nBywN7EUQKgxXLcQt/mmG8
nGrx/UjmtwGub+b9c9Y+qqGLqHnhFnBRYWsdemDaTcvWX3w40xq68Eh6Iv/BDtfo9vMxd07xnftN
7m+SV1o4Hh03BcF+nlRT2E/BAk+RcSt+UUx08zWfFal8y+6cXSq92RnBtcrEaX1OlXR+1zok0eCb
ww20L2J+bQ3T1YO4lP1dhkRj5cFtkozoAkWGThMtXVnOnJ8KmduQVc4bRaOMVoIG62K8wiN51v8b
Y87ho0HtN5QweSuwWHHHb3to+qTWTxi0nTDLJQ72UHcLJ0lUXnYwuOcjfn/HgALCPikToiemkxwe
ufPP9SFhwFZrVXebvVL2pIGoLqYzRrPIl104MUfE3vgQPrAffAKt83JVtRYTMyHM+CVfciygZB8S
ZFLCS8NYT25AE5kFBntM334/X6jYGeTN9a8Srcgqrs93hHJcb7XGEMxW4Kuts8mjeAXz8b5qUORo
u5ZlXmm5MGFxHULrv12mpAIDLPCCdCKm0t1nvichGGQ+9lcxghgMSyhEIEEuz4Xzf9UJ1L1WcCSl
FvsF7uH1RrblbaRUmHE6c3/7cknjhhelw7sQKXydAJbJgyRT/XgyRNKv0p+x4K5FZKmy+fOnBEoJ
PMLazKqhyGCcz8jDpmw7V/zGkrmoTzBUtyz+RiwbuTBf2I4bbauKs67OV0FLBwj1aOshQjbFrE9v
TpdXsj/JOyel9UxmkiVzCbwXrO8mrL0lCkqk4FWxNZTd7QYJXaPoqWlfZrx0hVFgqv4OlCFsAs+Z
5jpWTzCbswuzCWM2jjATJfFHJbaQtCN/yAE+VCqrEiLuyu6vcdMqSnqmZuKxJVmTQVG7v3TqGRsy
EkeYRutov8Rczm/Zkuqwh5D46C9XtuL10UVk2iYzcdm7t7nxskYvIWXEewgokat+9TkNACCGpJ2w
Zmr1XoWFS95cHfS1zxpQLI4LH1zltN7W2kGj7PZMC9pUGMr2YjUNed5YG2J9CrYkHUY42bVYFMj2
ukmHvrrtMSAi28qKwrF8+7sUaHLd3n9gTU/2E6wxY27WC1f2Dblk26NddsKEOdU4brkfrT+3icWZ
T3WvqHVRyxNyzKSmSEetUF3bX+ZnLQGs5EJ0kk6CaGBg2aIgXuKMaKPyqn4pNNNmE/yRcauxlIzb
XZyoK2bm9YjrJ0SCSeUuSNHtLqnxEaeWSni0w9Bae11siTCOaboCiLbdB5y6kFbL7JBB/fcDk6rW
O/M/e8U7b2mMnNJgkotb4QQwnz3dDEDnAW6g9dkkEJXIcJA/oBs8jDfwFqHbZnUn3pmaT5GGGdHJ
QZ98N/spWtYbjmXoeYVOyBUN3omKJJsnOK06nvgR6GbmpPYCMDtGxjGa4b/PJ5AaKePNhvIoiRAh
rZZPCR5fDmNlZ/dJaZLRvif0b18o8sqK7Ou/uMS/oxvUwi9PR64+27RVSwUB+8tCFfD/PzCfE93r
58IbOtN1N13YjB07C5etP9kyZ5GhoeD6DQMrPWXAFqOxLFcP29dqyFVi/v0bSkXz9fqPogrdA3zp
pMMSDV5s2x1wvxqU90vGYbRfzEeZZi+yLhVNhNuX5VJwBHFy3QQZkwdD52VMBKdk+R8t137OOVuE
LFxYSEVejWaAxDjk5FYJyY287exTdq76ZIm89wX3lbDv9fzDWGIHpkAym4XLiJEqHvW+frBBzW3C
gEw4SAihfUfMkZgdgchHRFs0ivsmPAAENRv0fHsV1P4KawFcgI6l430x14LwoT18zqiPUMI4Bd9S
hgrA6NB8SOtZjKUkNkAOzcbcTh/ms57y7UV3J9UqLe0HYF1JFgaOr+ms0VtbuILtnyqcOSmafUwI
f/tCdKEm63da5S7Bp/9ySv8EQpZsOq1YJZQOUzHidejisNX6CZohFS3AqTrAkaDvFXZvKZudnTQc
SGkTcVmwCXmuEGqHSdV3yWtWaDNzkrxKtYXIcHgZsJU9AzPqwHcQPcPZHkC8HyArEA1CnGrkbSMT
lqeYZXLCqQMTiVAptnOCPwNKvrNEXqMf4bMhJpOT1ekYHUfiFS+BRtGHsywLierKof7la/uXiO/G
mpIdMGWWPwPKVClKE+sX4ZRfPis2rRCMvOb9L9au2N7ZJcOBePYcEI0H4rqN9oiGz1fcgWBlWS3d
WuoSlIv1RjQVr/Y/HfjjS+HtPSUH0lgCa4Xa8j6NbwyYpn02iMsl4VL6tXdW/oKUGoeCW0kOlHn8
VVwqZID6uXQAwvnKZ/EVIZZNW6HI9wXSQzsAm2WKw8ZvNxzQDR3zJnfoOfEeQVIoWfi453MyeQ/G
IBCuzjwsUIQbBENug5YtrUs9UeuQY1ZG5rd5SbDuOxoH2yt6eq9zvl1BKwLt8iZUTR3s232EwGu2
tl7ylakTfMyz8mBghrxMkXb1XCmS53gb3rQWl1Og2EzKunEGKg2xQwxSkBaY9PmcvxwuhqIUfuvQ
RgQQgkQ4JCs/QPXxAKwDyaAG8fSbTK642kT9v0hJa2nTrvDQ+Q3mWOQxXsp1aNXb42puxM55AcDI
yLQ4coVcIMduJm8qFxvbVmkUfl0IwCBa6eQGvj6BApy56m5fO+HSRmWZtLT1S1MI99h37QfmhDfB
8UxzMKmArK6QqYqCweTs+aLbVGjBlU6FRKOlgVhvpjTh+sH2ShG3XazGeaoZxpVEnRiTi/KXFYjC
pIvDi9bzRYH9YjwYppJQ6M1l8RCq7uZC/4gHgaKQy+j9rjjsFsNXAZm3sTX4cGPuYC7Fza/3QhDj
ZdQMh8jMqf2U5IJ0z8nNNpYOmGdvBTsutd/tSAUUBffHctQVg1/afsDR6Y+m0BIMZtTV8systPgb
KpY1iLCVr2VhqZYbt5mQrOepFvKRc3QaER21HDqM64Cc4Hnvux0fWRlyPJPeAQwMz33B7c8WVDhp
jMpszW7c2tAdQItifYGYJtEkRdp0sD0EgWfd7GhRbdaxM+Q4i7JULbNINQtdKtbbALFF3CD1k7tV
SjytAtNOwAzT0VaA8+Ams6MP0Pgt7yf5FtcHcvQQTwgGjVnMzfKd9MHe1Tht9OtF4kWFUd98hoCc
bEy8SgmhSindQz6KH7IBhkFlgKapt9qCSwb5JIG9x5S6ivVJ5BxSW5+LQ0xqfOLU4LcsQ9b0QcSw
DJVscGXpGM0uesVLbQMWf1xp7mFurCUv1lagkyYHFebRvVHZdzzkiUnE6Uca9iKG+yUek/1mURsr
bdLTrN4UhQX8i4FYHq5XfoMeoU8teYofjoGCwnPJK3BEaiXyxRaIkcSCwzJJPnpvfL4t3YQBDmIP
/6CkUcmll+X6c1LNjPZrjQ7zcok73iKScZ68OCgCTj2eeLET/fY2kdsN0glExK+00eC3ld4sL0c5
izSOGiRMvN67ZcpXnoHdzh8G/Qk+YsTOFnHzix7JrBtIs3W5M2/n5G1QVcNl4YivW5qr8Cyhuedo
jb80uD4btzj8nlydXrXSPrHBg+W9CFDwbi0uXFahq/bMq1XZ6rRgPhbtSyDK2lSK711v3TrFPvmD
ZFvx8liTwEdcwkbxWn/KDIZ79cE7YJIsRoiPFy3f+1c7yqAN6IruoIIhwNj5hp8D3i12/QGUaSEP
5n32Cz3xwVfkrE/MFzOJ1OOuPiu1k8zPX0Vt1WKNz29RMCydhu2eylXJJXhvmWfz2l1+5SYZlD2o
8MdVYTGJ5iGy+hFuqa7k6jLs4PQf2NJ9QxbUE8zGJru49uTnABV2KyYwIPditKz7qddmRvTQrVJW
NggxXJzfhTL0QNDqqb0D8XsHoFsjsTZhOjZUyB/aHPxIkRRJrMA1ycjj1XXUP+4Y6nMbcRWbNk04
9sy3inBmhFr4rRwu+RKx+SfEr7fNnjna/JLLR9scw0IBkHXE81SNoVk6xcnXu5eJxEfy5YLsbXX6
O7Rs9tVc+N+sdFmdnOPYPH0XNmJtZCETXn8wTn4/CxxjmiXIVUgN01A9TRDKowsF4F5HYfhPkXO5
0J8t492ETrzC7BmrBsmo9SNKAizLVVLv9cqPl9DFW6e8lggzuZJN68CnVd1odoiBSieTMx56UIEg
25k+Hw0eWY+8ALCD6b2P8xnmZd3TdtE82j681Rnq4tCrkNGyd8IyWgwz34G6f7LTzAnSJgaPh3wu
oXuzEvpsTX6RbDg9fxF3rITeweeqPDjOycSAbMuJ3dH2VYrUpEFf8zAjqEB9tXjXy5VngW4eneV5
F09Ilt6ttoQj9jGPeSCfjdRB4wqtzDkELIgx824RBOj9AkvqwDSDwhTlvGq0uhxhtnVgyE3Febt3
4cWVnu2f+0vtrtOaSayKXXtbqoAUx4Dvnof2JrZOh/8/2FwV1zL+ZyzcW9WALQKljcCRKmF7Smj7
k3OkuQv6/nlJw5RM8A0zAuoUlu444Y/j9Qtpbi3MJ3oFI2FVbb0ViyF6hvwNbh0sUozL2lvPG5sP
x9Pc1cdf5R98rWFVhKYcmWXQ5Be2fFCjRLOmUjS9qf/IaNI5Rz/kWBW/9QpNWGbaCpc7SGf9S96i
yPO8zNE40YNb8oajsdFA7NancoWGaWqIhbqaWgXmpX1lNDCA8/BFuVgOGKAHrcEmSNnsrVM1d6LY
P32MtHpNnHqDMnJJSAgUO47SbNtyo7Kgr+dkzUJKVo9E4vzgLUravpa9/ugE5Gy32r43wNtxs6IP
0iNfDhtzQ8hSVr7rwvH04JYNJ+7AiUV8YIvejx3k3OWziEph+GspqpFlRfTzbjKURkSLOOPIVRSI
5axLteYXa0uW2eXuRbW2547m/z+dPAO+CalFWmfN3O71KhycMMTaHOr88bwkcsGuOZ1qrN3RtgsC
jRGxVHreHdUimlu1ygMrZ9kc4JSmEMYaaNyMiDzxrACMF32/x+YmBpjCgZG4HqBGan71UkK5rCbU
d1cLtgbT6LAhLjv6xxwK6ns2naIg9HsEYIHGSJ4DVkXgL6J2s+BSEFkDceaiHD2ufr7jdfPbOTN6
VqlxADbSl30jsJY4QBM5owF2ZUSAdMC7n1SWgJeP7AsgO59JqkjjUYvZH/7WCFosMYiBV0cLP/8d
/LwzSJa8qMDHTauSCXaefyCnYchO218axUCsijaBlM3wrDonc1/30YCzxG5dOOG17ZNTfRjE4EIG
N0gPEXAsGeUWhOg8r1h6vt1Ai1kQ60yJkE+qMJFMRrWuBYIxlFHFmwddhKRef4vwWHJXQ5avpfoi
1PhXYBmIzRoHXK8lKZ2LAdtqldlA6fA7aVzpwhdkfhG/JpGCw0lBpuJmf6Ud0nJ8kxyOJ4xwdQxT
BJctVK3KCr20g4QZ1GtfTZfufSCiY1srjiQhCYV5VrrA+UCAv9QjyP8NvCAv0AnwwrsCCbAmOv8K
zeTtJ/ukjdwuK22dpWUgDs1AJauBit9yipE84ugp3hxSlfGBpraZ0i2DsBsza5CYMIpyE37kpviC
Jik6NB+OGTU2YRvr7wcWz4B6lvuv66etXk6v6UUhrxCCKzI63LBCVSaW6wHouqQrdrruw+4SX+9/
sPzCYnNHovNLR58u7MwZy0NJbglkXQidvD3Zk9LqxlWMX7QwUCk3zpEZZshrybW5C02KP5bRMIIs
eYGkpTSbgP/qTK3nteSPhgxcKA+/hKknSkFyBrMqzF/wUQhKb04/TpaGOsAl22J7h9hF5xsGulwP
wvHkjdTXVdB5QCD5lHc7SUtnLawPrCAJkpEsx7CtbNc58OgMfIYBloay13oXOMPOkENW44tsYc9G
K9u3LG1ChejxQtXR4yg9MNEGRg7QuEEnYvPOIJpgj1Clat7g0M9WIZ+3lw425ctnZ1pmkAgJwSMf
hOYqqT05Lu1elYxRUWTkP9D7vmv6IO7jqf/7Dvd52D1zs+7JU4HFdoRDujcxULWwLsw+CxXGonUh
+qSo8M6YbdEE4mrTC3OW54TPX3JwPD4oS+bUv02/83HZ+VgfAI+OLmXdA+beCwJhSFNv8gKI2EaY
8ywCmp1yFGSzZ5/fPrhdwE93STiqqLlWjcFRY8nvSNt1aCCKWROM6wsLUigKtS/pENKqlJlF95cI
NNICquinwqimBF8HfbXxDTA63Hm5YkJDFZ5zkoIDGc+JRSYCqEZFl1rcndsgYQ9qYEZHy5kA2lYj
4HflW0/NooEhC57/HYun07aB1klzaYmjTjvWAtpd4N1JUk2RsjVh1vNVeu5xDkdbpRD4ZRMTVWQI
bn1o0VzYZlrznn5edck7+PKIncv4AnGg53xTja9K3ixy1GoBsHNAfoVK94XLq6vo8oSjnjxkEMzA
4CCK5S9RY2BOli479KS9nphJFGu/ditmWrLzGGe6no6e9VqfXYAnaEpOWVVWCWF/S2GlVxQgyUal
AEkgIkUiOL6wh6gIw/c9gXgqmNfgbtJCKDjAibaDyzIrDPzM7zhb7UsA1iPm6LOzHftZzlnuS0Mf
JMo9JI+QHImaIwOs1xglwDfSAIVnaZqF6I4ypFSclA1+V/5S5CarBOVWqbvHSoi2C1god5pKj0AD
H6AnG4DMAE7H5ehNY9YZnFtPzV8ToTHsJycD4rIV8yV7bgYZL7YbNkDcuqAqlk1of/jBezSpir31
DT//hSzfoTWc0hqyKNhFQqp2lt0zTYSlsjcwW1LEcODNZD+vLwiwVH1d+vW9C3EJyEk1NiYt+lh4
Wr1dITECidvlZiRYUwOqwcqmWF1E20OkMnAFb/UejA/Ei8NsWcTzw0PWowuDtu0DImaqKpb47sOG
Fl2Skv+gaVlR488c0kiHN71Upwz7Urw7E5TiK3OhVvcaitGlThBcj0rvtntZSUY+9IbsMyoW3JxW
cZC/I8DotOuPjX20Cy+KvM7AuU2QhqKOc7cM9/jOtl6T1lfGORIYxCGklJEqsSphzltaxFv0UFxw
eOS/IGmtPa/W7dNwfEPQ0ziEAU59fjOpotjFIWi6n0yWwozaLfNuQt3oBivCPZm+OHug6ZywMfkC
Zu9UxSv5E4sdJbzCPL3DX8kUPaF3vTzBqepxgfVI/pMvd0EXPhP2Cg0FgQTGTmbKUaxnn47DlkfP
t/ff7ebMBIp3MaZj3vQrdIofJbau8C+c8yfSEhD/+giK99epaKs6OfWGqM3K4koyF9aQK782taBU
HWSFil+0K2LpBMmJUQ54qdLbnMDKPBw8zHitT5xRgbJQ1Yg/FuQdKaxy7Kh6Ozjg9ikudrNCCdyZ
vCsr4PdbGNWjfgQPaf0ZXayXlUZ0zmPv0Wla3PPclKtsa+3wkuk02z57AMuCk1/dMgz4zJW+JQEO
jcYBh+YPcnDvBRnQYybVrTu26k4lJ9q9Q5SWtZ+oWCm1VeldSuWovIiM53yjk9ASIa0/xJCc3q5h
1mf0RskEEZn/hxhT6dkRBXUJs5KbXMn17TeJ/CuE45D2x/PL19DDjaakFdQNQVXLoOBUqLwWuAl2
56aREdwpTYaKCqFCcXDQrl9epF6Vm3iBuInVMUctZD5xxojY0jnVwNpeM2W9F8D4QsA9nuyYnzuS
kXOgIfGHel+Wr2ncMeDcdBcisE7IZ4LuGzeit6l+nr6Qml1qQDrpLu7YwY3kNXN6zGWp6l/hxStX
xf1JfnvssgmLgys2ae1V28mkYkk2WMS5VTjCqqyp3tmNw5KUArIGZjBUmJgrCG4IQDvddaIWgbdc
MuXu/jH5kzG/+0Q361oKUYfSywET8AC5+ky88tie8nqqPXU0bf5VKWTn8SVsJrZSb2KuVQA5XG/3
N9CnyyzD+tejyOxGfjouZPosyrLK6NlSE7Rrxf+msV0Gi31KRWnXET2whwx0kVCKGGbUKXVPe0nS
kEHkragNxOHHy1fIojjwcexlkEyTimROgLDydNi3o/XYl5oscAV3OYIgBAQEZBW2NebsphIkUetJ
9VKHM1Znz11rqRMUZ5U1oomGBNQhw57vKPmp6XdBw5FIrafD887jakOP6wjf51MyHu8CDWSqBed9
cl0KhbZB3nnGJwBcykqYzepfEY6RcLUqLFxLVwZRAr5RpCSsi7OyRlbNCW9Xvj4+VHsX9wjnXBn8
NTdTarJ29c39NHYCmoFnFWr0MIKGy+0AgZiEsWO9f+x3vTLZkcbQwzBPnYrXFIv3clNghjZgl8ap
Ha/3CQx+HB/5KwBpxu2I4CN4YotTbw/PMbsQ2EklFOEmyrvqViBy4i7wKkGROFpoONTa6s6lQXoO
T/7S83VVEECMq816bD0rpP7pCRkWlBFUf0xMDSA5BYQV+lLiuXEqD5JU4EfNB0UNIWA5rXIsrIaj
27lb1I21011cS2mWtsC42NIynS+lhUhcz0N//7BuyK8sSvQdyboGohbv+fYKm6+0WpUGtTBS/fi0
Z/duHpzWeYlD/YgIUVnNdq9bi9KQ3h81RnHNPpUlcGzMo0j1P+vu/WtwzxJoDXOce9qAL8AW2Rr3
QV9XxUebPb4C0eEEWUYHXExfA4xXjVUSQ5c8qh2OCnnmY72Mhl/Der5dw/JlRUFia5envV1hSP3K
m60k4VdSqKdTiTkYVRSWQEbPvBBIZpT00KLPt5R872Kdj6Z6sHqzvDcm30NqH/SVrQTNexvEof3E
wQ218uBRG6wcwVfDzlgSUIK9pXYKeZPBSdeFABGNLPA1TUd9OKvJ/IazoVUb5PtY6MYFoT6Hyb7f
fVLhmWl4QYiNUztaSlesgRFyeYXuzxmcB6gMvZiD5yjvZ/6NbikXOJpK8NsOtob01y5RW4auCsty
h2TgRpqLWwVVfutoqU3E79vMvtIhoBDyDEhQnmE8q8L71J+dbRjbxptKhxoSKaklC564Iw9I2TtR
eRqN2kM3hj620Fby5ZHfawgHL/+8jb2VR9xd34ga4XsxSBCk0FtuWg/27hq7pusA+ZDvmRqWM8NS
lAf3rzZClcJkWfQ/RlspJ1NzTw4+RrOGf2sAAquifnA3IELJfseCKw6J27ERR5PpO2PKdGSfq8dw
WF+b6MKmB159k/2fxMXkbh5MVxJuAUU7hiQ7MWFf0Wi3HRWSE8ck9u6W+JO7dGInApArRtGW17cm
7YQIy8XBQlDSycZDy3NNYEwKfS8nsDHpfjAvuKWDOanfXWrg0oGCG0P4ze7HemOwkfXYYOT7aY0M
teYsdDAb3SA62UZ5tXX3QUc9sxpRIDWckjmA4B/1KYunIG8MVDGuvbeXSjYl2yCNloqrOaGqfue4
hYBI6vqea8m6rppYaitQq33uFpohHNtFLIsIXQZv6gpokPnAH01Bw81YdhqTU74N7w64r82bZaPG
EOkQutk0yGsKKoNz3WnKaTT71wegcgpsjg9isB9suZPTR9wfTXqGNh4Ai7vj+UrP9vTCLiUZuW42
Wg+aMYIICvr0Y35bN7z9T4uwHNj5nMFjb0oJrYQO+k1yX5b84F7QFl0rJRiOeA0eesOZcZzNRdOE
aIRUwrdqJMgJK2LaugiskodhKkUtcSShFjhwhKV5TvAp9mxAOC84Burlz6TpjOJ1fHy4R+g5nvUS
8uXK+KzXhSNcsAiO8R16VJRDo0bBpwJVsprVpFRfG540X06BStBWcjuqlM+yALUgUnBRNiHHtlOc
GrSA3FYjg3miCnq3nBMN546c/ZJuVwryLaLOpSmmrRmaOIdmQVTseHTq3c8n0YLPgr4ZzZJ/sGL0
j7ui4yzJwpDcqyWOoz5Aj/ZESw8dkAfEKmdgbx6zSwCT8PLyagjHXuITku7KFprI+FOXVLhJPXP6
t1MFb2poDYK82PwOdJGWsxIdRfkar2bFv0bwCsTRK1NVrhx6cXW/5grhKzGkvVHefG3QGQd2v5Im
mvDZ35MGelKyNUVYSPteJ8egoHNMyZJoy9GBzIvz/rZEFygKFFozcLdiTKYnRSWcMqYpKGYeHnyx
cQoJkSgfmCLggJ9Sjl/pP9LKvJBjhQcIf2xXx6L0qN/xB/R3roqM9ha+L5tZWxwMOf4Jw/FXnII6
lBwaApBUwZcJ6A85BPCXAZROgBytS5u97QfyZKKsjhtQFGlCmWCereAYFi25N0YmPL+6YSzSLf0x
F1bicyWAlj7LYAvkOR5FG+0NiB10GaUb8M8z4BuRa9pJ4rL6ocs3e0+q7RXgKAwNlpaCvnf/mrt1
3jj24s/TJ8BipPPZSqJmOxI3mGcIlOm/cVyPRkbGICUlBeLh34swa8A0AHgkhLNA+ufx0/+4j0vQ
wlGdBo48nKri9dQSzXSKpR3qxT3T1ndUbDQ+JVl6VU/PM56StrCQWgYvh39jLJxg0f6Yqvh2sZYg
v+lFhCRbC2U68p0h2npJvKVxz3Yxxv7QGGcWEcJYP1wLEzgSAyISHSn8qUT1kL0tY8vghWL7u6hA
CkqrvvTrc0dqjNYK3rtb73LAm8+7ubmifBi3Cl5dYs7bYc5+jcR5GOKQjdZ84d+qAGnLNBJmQqdR
/0yOALvTFULRfWHvUg5qXUlAEHxByZmG79vBCsWeoatSYK2+Jigv/vXkW+DWjcjlpDAE/sh7qbtO
2vIq2tBnQ+TebeHVfdwamPJNjIjyx3OWtCHsJ966jQ26vOBl7WI04ShQlr+tA61ml98Joqk5nWWU
/DZrTyQ2JMixG8AK+qrUt4+SfuWjJTmF17Zs2B5nkzu5jzYFotNwBdBj2qc9AxI1LiEBbWMLBe42
zxKAvu6JRhUbvthQKQxyuE4SCbuUInKSKLJOIp7Kq5m7i5t+DOr6g4YfnTG+QJCDNL6IuxnrcJ4P
2FXBT963Rbh/8+hb3+qtDnACgotxXQbjpc0ZbXvHhserfUGQbU1DNbLEwS6SngM7ou/+pyQ9xvor
ncoX1BcRi1cyfTUiClX97T29pSFETesiY+jTlz3TATYrtQvigFgne4SGN+k1SCkz1nlJAVCFGjIZ
tp0B0UoKCeae/MGBU8NAbRJmFl14tNxfsFOKA9Hnb5/V3RVtQeCnSGAZCrNmtpQNbhQycaHRailA
5VoWDYNsXuQpYS1mpEqWWSdQynn15xe8titIHOJ4JV9QO18JjAoB9hnmkWj2iwEpLA03JbwVuZZY
Fv9a0GgNDB4PsI1YIXk3zyuIXftGc9hX6OJlwJW+DgAH9EYjWuLTkRiePsygbikavzwu4GnLUgjL
JjY4996XR7GuRq+EhUL69vt+y4n5RHMJWjsJpxvAXxuulIh+2+991CYeTesV7QjZ4CykSUTpIB0Y
DeiF44tKvd2/l2vGg9uK8eg+fJ+8Uix5WXrBywism4lN+KNJ5C9CnpnMjr0Fb/MYXG/jFTCZCJFm
ahUST5agc3KHHEBUuaT8genp52EmEwBsglp/nhunnl/+3dD//78Ul42pf93SgidRZRAr9Nao0b74
men+BZ5fkXgp1aHwS2DJcflR5yNhW2MrAaBtHjerCKUYCJFHp2pM0qc7zw7VtGKot5HR1IDKfNHE
vGe4Y6rHdgxk/gq/wjyBFGJNt3JKgSTXbWkcjqO7glR3JXCcg4jwZdomIJlU+4yo74C2wj0O3LjH
DuBlAQZkd+In2U1g1SqxKoXStC8K4KovO7SqWCXd34UkUaVZ7e5qoTkCXxsN9+cs6SvZ3SlL2v8z
oK+DACIq9kE4yL2YX+MAfx6WlmzVfuzHqmPshqy17TT81J5O+uj2mAW/CnsfPY62gZ1CZ7QtIng3
sIQBjqA5cHNIDczbOoOpcr1Fx4pBRdlz9qse+bR3xU4Fv+N5qWeQqIX+FjPb2/7TEhWQndnSsdPy
oaQndkEMwno1macoevoh8oiA5VC6mI7k3tYF/ImWteTe7Ue+proMZ8fH36wVSZBVe0uR0tYmeuNb
jVGbkESEGxcEnNUySY22ouY+KUDD9K3ehFBrmuwAvS5H/Brx/V/YbZ2iH38/zGXSW7DJX2RSGq16
GIcuRySQBKdA+g0qTvBvXl33VaAbD2KRm8wNi9GmqB2YmzLlkA4DwtzG6Ccto+gxvJ0tvQSKvMHO
2MqhS8YvwUUqaBEwnhtBkN8FxCD7hezjLi1E3jstKFwN0FyYtrMiKwMflUS1wMuiw6klfHFTE4Jz
XhcTH/yANL+Dxqv+mAxL0mKE5hUPeCYS7hAyp7xKYUizAvOZljsBC4wWK4E3FiVOzHMssUNMAE+b
JotqseTD8drtoLEpDyQ7Ojg+GA1BqMoHb6GMZe8SNyHNMMMgOXSpLCLjqSRdvFO6RHZ/Ft3/EoBY
4zT1jocyMJU1N2JPwHP9qOMoV+JFAe7PtQDul/jq86QcnjU3kISaLI078nddkP/Nw4Zz8eqNWN4/
goXeWJQEk89I4KHxExr7p3ZXImv14X1aRZYNkkmkPVn600yhvh6Bv4QXrYTxWusmS2lJ+C/Q2vRt
2Ntg2EQsxwttfRKH8GUhO3VVgCXDt2/h/cB3BgkTdMxaA0YasMqHBfWXaaRGT48K232uC1/HSF61
sJSbuLG2MRXlKXJ5MPHgqE+KDB3yKFwwS5l5Gqa+aJBHm1oSDfmu4JQdDHGThV3cjO2/UbEXpVWc
lZwF9fuHR9TdvTT/kdVm2tRyrWPcBYmtTz3O50GeN8+F3vk6AvGkejg/iliOAsfwG+Hudvu/eyhW
SOIvmdjKO8mGNDheqgYeZvjCgM2ZmUWhHHOCBaS4uOF6hD3k+QQWzyBrkyzsB9NfLjRPp0bcQQq0
Ua3a9dAESoS4CvhPIml65cLGTgA4bvp/JJ3R8YjGqbdd5Jz7L3k5kROT7TA0GB7B8zS/JgThhyMB
RTevfu5mevas4gkBkRyx5qeY72WwSx8OlIZFMWvft17GnCyfMUAhYYehVi+KmyZiTamz8KTNXVWa
LoKjtt9JDQkXu/CKT6HW0Q9OiGRc4zmJN7O1RElDmBI/84WoSgIp5mOSac5TEyw7jYKvCTMi6EDA
NpLIG3BPn0c1bG593PR5fqZl65AEVia8gekaCcaYnuQP8OBoQMuXnkiKQbT3fnus2ZDMYkLi075t
CYrIgZ2AeK0rMKQIOjwrA0/Nj7hL+dAn85L17Zev2VWCk6wm4E0YLfy5gqafA118y1pgIRHHlRb9
/KJyWknFbs1D7Ls7RhobXcUl0SAxh7qkUEN/Fol/sdSATJMSN9mkGilKp87yn7L+OmvKnkkvJKWZ
BkNEl8emZVRjs1EV8ub2u1bFs3Na0uqT0J87ITlTxJGhTXmQEvZI34UKj3N4kjR87R64G+c8DpaM
okw1sIXvDhBkvUFhBPs/sV/6Dq+XuSezSHEVC+xdYh+d+QcS++RgHjFH+3QWGgJmi9wbzQx5wy/H
FwUkNgQajx2SiRbgLbIrpYSVEh0n+OUpkwaXNNZ0q/UwUVMoj6OLnWlelQoEtO+Ru8DBnBYcJdtR
dpVSSixoSoOq7h2g0AJdClyqjvQE0w4+CZidQFcIvGFqfIsSvgLeDXpou5Pug48zlcLitavh7r5q
o3i5jpUMx+4VFDJKlhnHPTNeimgloxbKYv59xtGnTpaReX/7ZexwL9hCVP5jIVS4xCr2/Opk+jL1
KOEloh+R8Aw/n3QjUY0wTLCV0vueMKubS1GXgBvvUZBsSLh7NZAEN5ANBM8FOR+gOtDPv6znueLm
QbCZvfcQlvwtLGE9gdID7X7EW+Q7LVmdrYn7jMDN8WrQua5398ZrkGcmH+4EHMBV87b8jXzA9H5x
577pcfXX8ri64jS0GNkt5T28c2Rj1tAnYbsvrLClDVzSi42shhuH+vsyeAtFIBW6O1Hz/z8aaUI1
rUcwKrCNnbNH6RRAiBFmgIoX2SOKk2gZlLIZCPuLt04J1FD7hr/sZ0JWJeoAd+8aP3dcJF5jiqnS
Y8Hf+vv9KW7h36gx3YbIpZc93AOZCQzkg/772IwcPQTvVio2xa3NBb6joPHjRrzv7iel8XV4JPUD
jPHonmXZ2OsCpXBwJ2rLIbFDd4qQj96chW31+Lr8BZVi80lgiv0JQ+DjHM5rfF9mHE5dHkalYr4w
7HOBC2xsbsyDiBW4rfCi0uqa2gf4dUYw/aPgFIKWrQlPTtLmoZdF6i4O5KVg24ARCxwCNqNmuUyr
9jk0oLX2atuASvL7s38UNv79VMU5CmSgOFLbcPP7rPJA4UUuTSMc/B/mU8IFpHaqx93y65ZWOoHP
LRb4Fk1v6Si+IeoEVgbT4lRLXbAgVepQg/QrD3wp/lQwkyDAc9s3xSIjwgTff4y5YVkVyPEq6laM
xEMRJCo4ROlCqdD/iP2zhTFjDoajNpQHiqTLaSOp/IfdQmJgqHUILX4OddVaYvHZJ0Q6JX/H3FQ7
D2S18BEbvwmfMciW6haC6utVNxzhmGZKmV43eY+ykUe3pHTcY657F6v3BFzoWJktG+rAsz5eNEnL
C1e2bn13lIha8qY+dxXMBbVkCQg8yOSCZ9M1tl9vNbt6zRXEkIz1bazNhHfl7UCZD/JKWR0LWB2j
b7slm0zAvIQnWCA0sMSRWdR/NFliyBWqnC4UAnF1smhfXtWXgi89U65OCnq8vCVSmfdOE1MpX9sb
oolH+V9hJeJzoPtfI4SfzzxuimcKBwyrK2vprTRDUP8rVGVOwiK0tc54cnG2ztiy9aER1s3DtTDE
/l1BHRdW5zyNGtNjIjYjFHPA4jTyuCunIbV4K8Rr03Pndq5AnROPPqYtSv93POglYjGVbaCgExAp
PP46TlnsrDjbFoSg2UsXiO9Er0KG6ClNcUkuLdUQIThPfNyTsiXskkTFFbF/H64KLcR4AsvadkqY
1Ez4wjikkx60dZ4WZaLFeVI1VzEj+/nm0EWOOPTWfsmUqhi1moIrDq0Ys/4TnoflS3XuZEfjnsGq
z5x2qx8iIzV27ncwWvG7bftc2Ma3bwXyXQHNNEvR5a+zO3+olzi+LvGEujb0fYC/4IYwLVNnBx3z
/VOS6d4UoUj6179OSwXCZKR4qG+9mBEzGpCq3aksAqIZZfimvwzjc6VlQ+4JITozaIpWEkUG0f95
DF5mrSWgzWNd4dQFBCZtTdGYBYF1gAXY+h4g4JzBKT2m7P6b5HJzdHrPqmr/u6QtM7QHyw/z6x5n
Y1Ci5URlr93tcZ0hJ2B58XOAseziDC/tgfPhvbQktCeGvyCAYAPIaGFYcD+ta26L765XzPpay+D7
CXll0XDFFOnKqOIDHXk4/wH2+ygHWJ+UFe2Po4M3o2cJAzE28Bp52XOhy4Usq3Wu5rJFY2t0QM90
IfIT2jWH3aFDUUlBCrUY0LjrXwwJ9iOlXzewxTXgPeZJpZnffuclSyR5YhhEYFbuTMsEfO0Fu8kg
JqoUvUOvlrKR6vnPH6j1aD8SJHWUqe3VT+sYR7auLxKE4mNYaCEsJuVOZgBBtFjxUnXBREmMO8XO
dS5ZXH28RmN+KlUO0E055iD/VM8dAbUWOh3ntO6J807KndQu4VlCApuoE+hlo4TSmWah5SN6udmM
U5Rc0KWoc1x2k8KxUaPn93HMoKI+PCZbMRb822l3wN455VOGTRQpZkmpbLxD4gh8fBIny4wX2Alg
aNjmNhhT46ReFPmzH96LvJ32kKhsDlFWn8Q+yY3YDNM95a3ioLZ+jxaDdgaukCgPtm17qI1s3gv3
sPfoRM4BxTmrmM3WH89zfxJ8ekHTR+hjU9klY8qtXbHXxEIGsU+9Gr+YgBszpP3AE0aEtTS9m6w9
N6iIefDzetqvXWG+SulRJCNvLVhJS2DPiF9zy0A0Bm75LKbhQd8QlJE0sgienbIhrJ9qZLokuW3L
bf/itGaYnzyuQ2hFhHb9D0eVYBhhTP2YqsK33aUqCEuRqLiBWdv0TYomBwiJR7W1I+3qlKhGm0fk
M/H50jMj4XAcpAskuOatT58KN3IHAen0fTbj36dhDkTnrOXbKRYDw53vizo1AfSWjzaRLRieGPxT
NjGrls3tHDBSW6kR3LXDuw1KhJviU3is5Wfdk765oPeI8wvK65kNcRoyMQr0bJxoZA/T2FmZ1Y1M
TjKGQpybXagQkZ5fIZ58pgG5RxS9bC09wQfAjxVGilFOplV7FexjlV6wB8ofA5Bs1vCxecjwjdnJ
3TJ4Y/CCUCRAs4DgvG9JsvinjRFjpFagMP9JDjwX4ohS8lNM2gTJCaJXx0Wq85ttPzGcrElKAWop
xKiacETwt8QQRrtL0YYwCvan69pc0To3KnXW0rNHCg9uE43rvwq6v1g8N+E58EcPR2ELLSd+hKY7
DrBn6ES5dxpNQ/8khD65AbYKFdKfjYtXOH9+wnS6vPMr5kiSoq6S7gfv/hmtf0wGC/s3jfJ2Rni8
uL0Kz+tTNibIF22G2A2Q3K/SpeLPtzLeGZxISR8xMRbF8mBPKz53aLIhWpj5q1Oi/Xa3OH8289VB
b18hk0eMT/XO1VIEcjH4XMNkaw12WxM7NC9OnKDb90y7DE+x/Af8LgNkl/v0h0E5Ct0zM/uXhjhM
WOZzelDUdMtVuNu8xnxiSKH+IN7zs00ZXsoc4U9GGCStZPCplelDi70uJh+Wot7xX4fHyBs7YFyS
Y7IZNj5BTM8w6FBoK9D1K6jaWtTFB2aATAfHh7p0p9J044YM64wpXSaj6GgY55UufAPPC5sostjh
oZcQdrwWQZ1+lVmjFEqtJB0ixkj/NPCnU62kbTrlRu0SyRJCqlDShgp4g9rAEOPpPJlkw3rBKgxG
URuc962EZggXPGAGAntyzHChdoqb6W4pY2TImhaDOb1xfrdupZUaFoQx/VBa/RQFPJOfEdePNebH
FeS706qT2fa3r2BCVTwluq5hlMxLl8rDgJCiNtq5tDd1VtXVW/xJElEjVZZiIi0PSGQDX4SCTDuP
pZWXP5+39/zVroWhyV/xGSWcqPbQspmLA3jBhHOJI9BGYuUEH23OLXJgihClNZKv5HHTp3CqxAXB
iqptm3Km5ZjelWIM1ajx0Suga/vjIwVx88qSg0m9EhpPRLlVNX7Pe0XGHKcA7u1oEN125/tTwGQq
XhDVXqWNNgpzZliD0w6O8xcA+P8GfA+DuL9zFZAoc8E4MgExI3qNoyQF3e2i2Q41NenbyF4a/zcH
EoHLKzi+B9qh7tQtVHXlXyX75Zbqc9SmPt2pbPctJiiQIF2X2zpqNMizHB7oYQ2t720NrLxMGGcu
o3A3h0ywetfB9FbrnCuUZUA9yS8rAsQmZm/41sBB6Gh3FtNp1eVjUd+yPKsTrzvKynu80Bgsakjl
mBM/XIT38FvTCaBapzo4ipYNYGTYRSf3Qal8UAePF5IfIripYVgbpqsH4QCK4WXXhHpDfUTBsU6p
gE6Y0cU7xya1qyOVe6meSFGWNY4xPt7gnu81bXWYPUd/y+qYueOvUzEMWUebr6HSP+eMXmYUx3OW
it1lyUn4O0JZqToykbE86zeyc7l+/5WadRKO0rGN8Ivtu3P/a0IJxmKA4gXJq+l8G72UiRvarwza
iQoVp0kW/TpXJPu7MRzOcBno/4NnF2eQImYfPczZCVtBEv5y+XshrC+VeCYowm34q8bVIYnfl71u
8SOYJdc8uKJeu660FgcAi2B6HapO1C7lXSg1NmVxR4xwCzAfrn6QaQBIML9/TZ8SEMpRK2PjJZoC
HNJj7qXvlC2gIXzaKvPAdOYMO5zWb2V4kjndUh2/c47raUiQodbbSsbPAeaIMk29jEnYzLObRsZv
HWFqYvYHpeZeDEIQKGQ9T7+EPrFIAgvl86YR4Z5Dulqj2qzibQGQGvNQchGUxVeRIE5EqLLOWbpB
IxjoyNOnU3NPk/NuzbUnzKSE61hnMu8bdyg13sJ9LwZ2XcZekIobwuLRMFSCXp7M4c5VDls94qf0
Gg7xdViX4ESLbIoTb0tjd0B0G+8hsqszEEjKJd7jq0FG41G6xUUB4tWZcZqQ6KfFI7cIS6IAOj8A
kCAsVN9qhDHJXX/q1mX9k+oZ2b4yQXtyil2LvU+nre/3zwa/x5AKuxubDJkPWpJAivl04gcKVtB2
TXE3yoAEij+VWumoG42UfNnnxqwSmmiWxPf8pfx1+qAgUTipHisrbOUs1CnOTEU33Kc+Es7W0hwn
k9Vg0nVlMeh6NOT9rTZqY34y7lPDMA4PakbeTZOjcYfuNGAd+DWURFK28jtmSFgQuhx9T7GU7AWl
OenWtpjkOLwh+gh3mweteclXZXu9Mk9PtB+dK4ERMtAp6YO4r53Bb6WB6JP87Q+NPGuEzcHe4vl5
c7zmlbEJfDsio8eFJpEa4so5f/HCKeDbY3WUmDLoR81WeIx47Pds+A60B8UvSc+oOSqv9kot+LDY
tJ/Y7aBG9KcO7od5GfQnZ5/P4RNp1eiNRLmW6Uah7MqRghgeNY/vhA0d5W4Hww8tD7LcFQ0KOdHs
KdEutPQR0ovinBDxRkLawdI27Y892XagW+c9au9AGJlM6s+Fh0cVNnX9OMFXqPuLqkH0TQGmpY3z
+yoqHXnE/N4BzFyiVBMi3BQ51wYyu1ZAYC6q9PHEOWu1bYRJu5/2O6eY9+CxUZhtTRSF31jhaDr1
4mY3cKX5oPfzP+JEfDbekDrWx5wzEftYCvGm397xOKyhanCsIQAxptchmxVd8qGQB7+jKTzlkvdJ
J7GitWWJ+TA7QqdxjQR267DvXYWF5pmE7qVwPQzw4Q5zJwIr1E4SdgvHa9ALZQlzW1eqQ8+NmEXC
F3ZkmaD7G26B3yt/WwwsqfZm8qQPdPvyp4Ge2VailbeqoQJbXhvYZBKwmR0y/T9qgTWBrLl2WKPm
Gy3y1H3WEC1NPVc3KX1iKEA6BQZigyjUCej5LS5vVPh0dqRg7EOlk6rtGXL2sbY8PRhn+QKcm7N/
sEo5yVLvDHdRYl1/f70H8084dMYBhkUIqnjSEjkL1l1DI0m7y+YrkdGYmw0Czp2d1SzvkngzJE3N
FWSZF3l6iZkvZ7dUi/35TkHENmV3d9ckAdzTCqyl0M6GiFuaPxJKkMl0VuoTHxcvRp+tjbnHYXTJ
ByE4pH1DYB8cHLOkfsVup+rYhRPYQCRBD16c0LFcwXKX5286UhbtNTHG2+4yznuVNOAllHvfRdJY
3Q8dBbsQlmN2gOh3yv9G0Bdy4kc1lsEPohFZf6sIEz3K2YzKi+3kYsrRkyegmNadfpBmfsUbM5wI
70RWzImEVT28CSn4Ri720iLV0G6+N2wAv3fdsuQShvzf7r9CrANL/0bSuVDQx59nef/QKsGL03KR
FJvE52xzmwfxBbTbGu05DcR8flFlxZ4vfHPMlmWgqiK6jGEXeL6NbbjsxMUdl3CyoMxLSad/Tn+1
BUDwcOqKC1R0eMnw0x11D7bqrFji62gOppttppOiw8+sHot+xRh6AT3ycm4WcpTNIMcY4V5CCBtl
Vl/gNdBv3WwpCgouaIRnN61OpdpVdqrnnJjuPVPRgsv0GJ/9nG8KCLx/oYIBy99mEkUiZiemW1Ay
nWNlX8MLL83mN4007q/rYNodbdeaYJfKcgDIy4wu0THMN14L/mAi0mcP9WAQmMiOOHt0nzyXARKz
S+0vIqOWMkwrAxDYX+soOVtsRNlUIdVrSgeGIp4iaoBVSQ09iGC2fvBpY3bqHWxzMOb/6n+wm2Sf
SUQNPgMflJv4Q3Am91dwappxWf4Q8nH9NWAhEwhjufQwxy7E6+MRYlaRnO/m2fMtoZqxgdXNb59a
qhv4pQnCS95IqnWyADM2nG3KcsbFhU8eB/3G5GjGd+WvT3ZUdaWmckrf5Hdy1qiAExPUWax7kFLY
XbmJ4IyVleqcD/5Z/dgwwscy99VCwyWj5zNyiSv/UPjDxB4b+qVDHBTxbcxy4BoAaPRPOQdCoaM8
jWuxUQvMn8/jAZDeqKm1aSjcKMS8M54+cSg0OZSQXoqWC767rbwATvm/GSKj9uIBHwhONr7D9ypV
g2JTYM/Alkl8RWAOcDeCzHKY4K+tng8VYceZTM5QuvJ0W6xAGuE3lvunh5t1nJx6pqmiQ5fQYBzL
Kpu1hcEv7cUyj6rOtx43WzYwGlNKXyW7DZCJTl0XWQaf1lQ/L2BqTKZH0DHP1Ao1AkjceRkiQdRW
yg4hHa1CtWsM2PuuWBEEBOLGHhi3p7AFc6APZS/ow/ODKf6BZP/e5pSRIzTkAsKFWwX4ptSGNQ9K
rZgMIcD/2wUQBqYA4P65vtI3qTx+mTf+4sK11zyjXR473i/UsMWShPwN/xVIbSYvI+yLEpQ3n/nS
EBfYvcq04k6GusinXCQTWkpBGigKavhH31UB0oWcjs7tOA6DnaDShWQ4dpCYmaL6hBBgZel3JtEh
LDknSkabBdGkElcpeDx0S15H4eaOgmWPn5/XQeepXemXiOIRd4I4AmX7sGMm3hAIt4AbczgtYaIq
iYPMCJIRBqW8aNZNOpdrRXAjCMDa3CIvNe57st5Dr5fz9wDdQdUVjOm4jC5SLWDm8G5eWcwJmx+H
Xdlkqq9yBer3JG53+3M4y10Vb3ayi+2hZ60CAAEYadMNXrMITD4eJ1KwoDEMslbNOf3Ek6nM125j
+WdnOVZfUM+yLsezZnPadD2c6TpCJBacS6WPSY3MK7qdffNkyGi3cYi4maCiD2jAnPfPXHGzrhna
0Qc0VQ9kkghO3xU/KydNf8U9ZI1X/+mrlBbyHxNjw/QZ2RTn5jqo297CDqw6Frzeh2wzR9Qm1yy8
6RhVLSYiB5sjuCWxhhlsyMQBTAoj0OQ0F2pbokIYPF4gQjdeEmbcaOUVwBeCJr8n7KgLsjh6kqae
92YfESbZvGEmb0hkVRekgSplhj+Zox25z6QYQpdM+IRbLXN/uCuZpc37KZghK4rWMFLkvso5n9EM
yFlXQfabevZGoAj8AtBvVAzwhzmUO9/95zBNFIPcvk3k8ShVZMvRg7+DhHPQtD+uAXOrQEp8byBL
lAjSIbvOwTZbb9ZS6smher3wViqo+tKVy0YWsCbn7fvdCiDI/UWoHs3A/XVB340TUzwM6whZKE0J
/lNNAF8rrYqxA/DLbJzBWkW43ytRDb9mXp7J7imTjfx/pecpKR0Xp6IOXH7ApDcndNeVpviKrPAZ
8k99YDUefhEXWllYaPzymXqAOlamBrRqtRvw3OnewyekJ5AYdnatDu4E05sUdtBdzvTD4S5doxRV
C1vJjbj9Hd4Douq1LWV4mctWRpVLpw8Qg73RL49zNCfYsHm6wW+xqY8ussoL1cWnpL7FYoShNsrf
Wg2i2K4BC+aSppP4e83dGy+WBZcRYVEvmKddaujpe5/MetTAyWDXBolu/LipEL3jKwVX9oPF3t1a
ZUJ8kmIMbu09Oa8l6YnQDzurXDGbS7YKfrg11jm+srdBovn6mtCe5J+Z6YUFwnr5YEwtfWoTYA5S
szhZ4fcuO8CjNECbbfjV7RD1q34mMAwPBq2MRcDYU6ywAcV7jIVqkboLEgDoqcv1VU207yqTBHFE
riQyssVgPJo5GJflri5/PutmDla+0OwIT4BulGOmTkSAdlB4Etdv5uR9tljpIL9rSb7+0imxRTEZ
dSd6jA01V4pCfWJrcdSbIm4OjmeNpXzLpUA7ce97zDx8S4VmHMLvRlzeRXkQgOOwhvYha1JWPnnQ
dDCjB4yNrlaRKr3tifQoYeD6C0S2x+Yf2n92y+FmBzRfk1pluRKCZ4h5JpNfuI6BhF8GDBYnYU9H
sRuf55ptGmR7QfKpRYJyHUXh+CsFIlh3PtL6NHNk2+m1oNoCvMhNMQNTnoRe+J/lD2IC/5Hp1h9w
AQmISTBCEckyKDvxCxfmvSwrRYpD4bUoUV1T4CJAp0qq1njYMNmQoGqyYmoLIW8D3RLHlBTn057K
JIeKECdhS+XCpusYpKkbq7y3mFkJX3NYF3MZou7Sb9xs4nnnu9iQiQ3ucZesqlOZRb+umrTjIPlA
uCYkJEyMfVRSiGOUKCv/jVac9VSjnoG+IaB8GXzN5nfznSkn1LDEyVHBZ51kEfRkfWeDSHqZ2nWI
o2QxPU3uNlVINfcztJjZ9dFG8p+vMf60QogGSbctWqL89LMs/3teV52k18vQo+bN3qPCJRgZid1U
ej37odu3uexe7Vs/nBLcNZhTFc9nmcqHjdSxTniGPSKLZDLYR1sIM1mWLe4eC1MFq/J9P9o+Q9+k
Yw6oYJ3GUulVRi3hBnCWfKkKzzZj9/kLzDR+SiaGgaWfsECJD89EDucAt/mAyqAPbxnXIKd+dDMe
n2RpWkRuByaY/QPeEEQnuemeGCE3I11MYh9vp9a1cBy66gvZ5Ta3MRVgYPaD6THdsUi6S0b+VKVD
0U4+MEG1MNTfxZZWdwjUUmQHVFByyjlhU2HbVEaXhgZ8A/TokgHw8zQSSowMsIT67uSvKQpV5dUw
kcBdAPLAoOlUuXWT6UnhlvMRHVsZehmDNNwozpKDw1FqR9DE2y+aslb8JyI2KGGOaX7y7y8BOKGK
TkDzuyM0HAEA5umxt7gX1/DJLazNiF2ZYHF5v4vDi/FCt34WoJnunptQ2ryYJZ675OGq66Q6mOzm
5UIGDR7abcC2JmZc0/6IIy/mFWJCzhR6081uZOF9lJnmRgLW0I4+Zb923LqYY0fj90QVT2zyaHea
LKvNuo9PMMW/8elBKaGE5M5T1eVDqiMg0A3VDV2VHSZxYQ8MOvolDBMo+6arq05/XeowmJUYhww1
zKlctCCyingRqt3zbTESEI9KMWpaQcuDmwHFwTkEkgXX1n/25+n2Ijnkzd6X3285AtnmGZIfQNBB
6OJQfA1KsPMimc3W6XRr7wChJsuil5XrimmPnuDp0dUOBB4tKf5BStMCXtMczwq/z6991cewFmsR
HNz6Se2/AnJwMO68oyKINfkymgIfQS6SeFMyiEyvthtElAFcY8jVmO2b8+nuHlVP9XLCel5qL0GP
9u66liNMPE2mnXj1G2YGM7Jj6v34XnGqRdV1BNKSW3TmRJAbsg6COGBPFczq1P2HlQ8zg9EG/a1B
1EnsRLtbOyucX3F7hEIFq5z1UfXd4eB4fLMIz5N+Z0Gm4wUIE3rXC93t7MnHaDJZZa2XPROUHc0+
nB3rfbESoLYpurROeOBs9zmpjy8idRfuGcSGGBSsQA1L5cnIC05OgrzF74YPvCW22CiiBJY0YN13
025mPrGWsqBiItz8brAeS1yGT0TBuqumHlkvjOl3l/63LB/y+HXT73OIGt5NiC1YJb5iQ0BHZh5p
WthJKvzxfeh2rCAk8Xmx2IF/ACA6TZDgGxi0mQE1TVFtm4w8UUBa+oSGOmK2D2wMnxB4W3qrkLuL
roox36jpducpmmeI6LRaWiW70CUGJa7oODjX1BzyKYm/rIfe56TPlUOdbi8xaYR9Wqy5nYdOgc12
2LB4FfO75ytWdMIJQdRMSjqv10pWw9x9EnIMWglxYihOHqR6W5brjBpwWSljm4QnpSGc3l9FtjbE
NTAjbLsm3TTxMP7P9wrU7Az27+zkIHkZCCghQ7n3jd/g0IvGXoh9fRB+k3cPkKJxQ6LTv7w8A9fL
C3sgAA6xWYukCc9L4SFw0W2pcoYej5rYLaDstbj2YP3/BrPzGnS5gVgJ5eVwqeEnhWwpOfkrBT/t
uo3+0vNWYQ3tqHeMJE9bp5A4XFwWbCVgtrtv2s7fhidtby7T10CSC7xaZrK9hK2og3D+kWHOgq+q
F2s1pQr6G4DjTdT3EDA+gjmsmfTa0Wxiz9CzRumZfmwwFEFkt6VKWlZXvaMiHmvtce9x+5slRJsv
6pE7udMhR0pvOCgXa7RLZ+ioMmjJqjaQhub4WviZ43iGpBVnp2yLwsx/0qBMoTU2N0unmd7gAD6W
fNGLRqSYkWXbcx18V+JEc2L8OK0pIme1deKpHPvNwIMSWM6sfoo5rWCvuh/e7T4SeQicKZdPaRui
GpfC5sohz3WB8bTDVh5vlf15Ym61LFtxyqDFNkhHfyxvCs7G5AsAWB4DPtVyqPIFdyIL+swuuFxL
m4Z8r4WbLU3iQnUDL2DvXgkYjIJMdtB3+ZN4Dg+eAF6a3hDBrXNcwsamWjnMMxK7db4hM98lfoNU
5FwlVFuw20fkf4CKwcfiiwH+GLNa223bPALrosJXw7d6MSlXmMguxJemuBEnQcdVsCNmF8v5rJ67
5gmM4fMOQHjG4mHi9VORPHvIw65uRuuPrYqUHB/clPP/ixsPjI75VHg4vzrqnnYibg/LXX3nvdY/
tFfbZywPPkQeozfqJC5vjQqzv6ImI6psYmJJ0VN1bdzG8x2uiXUaE9e9wR/16YPWW9xgvpNZ3RSg
xeIR51EIG/stikfKitYrwT0akVyX+T6gU5QccJxigvJ65M21u1PAVD7PaZb/wPnrzVFGG078hxmE
01vR6chRnUMyV9ytncDq3o/yabPe2RjKq8UuuFNukJCq0AEccdgapOQrkR7Ar963SnBREI+lmfmI
f+QhvlU2GAX/YGkgfl7Zl76RZ88t8LyuoKF4QyISyUbffT1kgYE5qf5FqAVx4wLJAflxFplndv23
BYUbyNH9ET6NQ+X1mX2VOgSuHI6TtoxjdBDt98nPxJsfNdrqfBzd3idAG6fifNNYKXMQ8fh2vtFr
WJ7UMzRsALT1m6wRwYueCYfhiw934poJIPf8IRz89nX0dWVBaJKmCcGdM+iLaNre1q5G7pBfr2AN
TpnqLEmiBXn4vZ+Hv3lwR9y/qpGeKyF6ZRO6NTxHG1bjQcM/utMddn34sCiw9bq9ph09cm2zGm2/
gyl0iS2HCDtcm7N/So4zC8Yc//662DvOJqYIAgPovS5KFWsVFY5JvAG+PZla2mBOl3wB3VICawJK
kF+uY4KDl4EWzcW3sTO5N3JDkpZjsMclOkB96v08vYgUFAvztG8aMKoVgmDQAVxPpzA43YGX1TK2
5SwFWiOVyrL1rFp1k7znhHiNlkl05E5n5RXCeDq7uDyN/UIXI1iGQor2Duq4MUWJtWpxqULUSJYt
zWkbCu8FlDeDsPhgLUo2KMz84agBreZ5p8qc47HDOMorTCfYgLiXdi8L3gV3Fc6QZ4EpMWDN9A/9
hBymWJt775RO2lwX9DwVG5kxel0AR+UXkCEUp/3wpA6jArCSECCt+T4acM1NnceT0bSx0OoOPgzN
sW0podRKr9OoqJhOi2Wm7mEnf1TM63K/TTt8nt5kngfR7ZjXujaWhRt645unUP6YuWV+T2ek65T7
jinek7q6Dt5+VOQYQa2ihU4WCchs5KOWYysDNs+jZjZCdIyoibzhaQs7WIPrLQ3BHJ9xBCnXDAho
CToNRjqTTYr90xMR5PsRSZNszbmteLg0bQzxX5LQftN22HTxngugGucY8Z2retc4hp5o5h3zUUla
qmDNPmmf3Txn3UPn214C/gdwQ/HBA2XGXFqsYLkklV9aWKXcsfj0Xw99RBFB483ozvidLwbR+MJQ
onc0m0BJz8+tu2u6gRK0AdmRBgqKfHF9ciqd41fWgJuoN5E5aGfjVAUmdBVjVo04hXs866/t883u
azTcVWtcIYQbc/y97RA/+oaG3RpanAs2iPcMCbAC9nBFPk6jPL7OrJi22/z06iqbpLbhaep8zRJX
V4eZ/YXvRBDOIvnBjXF7X9V6dNX9Py1/mR76P5e7qkW35fQxA6QuUG/9zpxkRuwKwESGyQoWaC7d
x3dk2AAT5e9rLRK2a4EmAsiVpgs7A4aYQ2Cd8Hl1n4hAg5RU6qxPuuIhj5RbzFTvI3DagtbSDh3G
bweqT0QVHZejtNUN2iAWq794lLiq6WkIJ3e5nMh1T4WHGpipb7kZPlDUgWBwcxA65h7rAO+eSNmd
Ji9qP3SsnXLNKaSnyGjSIG1MZkleNFDZcHG7v9OdO5VcBnmkXZdruGcwxaWlXFzzSg1c5cktG/Zb
fF5/5dR3xSZe6NmxesVXnRiOSGM46pMphdDXa5oKnr96AE5QbO7MVsWhFLXBJ+CEEnEJaSW7hHah
1+0qDevakjf+pZPhQYfuOj2UFu7FGeLzri83yl4S4Ofm+JUFirqim2WJR08IxVauatLKnnD1uss4
G186kUHqXV0ZXd8lDEDLFsz6BXwpHizZJwKSSwHzqAr0vdEnSeUUgSgQuS5sjLTHDPb9Epw0X7SF
q+iZ3uMlMXFGYA0mOCT/1Qzd24OalsXG5bXDAvPHRsx6z2MXg9o4WZYr5N5DMraP/dNdV/xfgF0T
Yoj9R7WVQe76aqtmTkhjgnJM75/08zwop3jwhIo1BWz1wrEiMipRQ5YxpN+FfBMOLdDBkPLDKxTd
LPET4je0IsDsKCfDY+wX0h1NiPh8R3F7oh9KzMBiBFF1EZym/iu3+joxNoeswwcUCqNjdwXeFDCv
bCLiRlrUcfY8UMcwa0GjZ/wchWNyeqy7hQ/IKEQAYCPMKmWFLC950A2fVD7keFmPFkdyyHSFEZzD
yk31n5iDt8QrdCUvPNHN+IwCgBh80IPhaY0ZUHxWOH9h2Mgtm374tRBwMlBOEuhOAqf6mRJLm0eA
gwXHJhSSipY4ccJm/GLIfcO7Q1AIEL3ElGdbCdU4e2wPmXV+oEznSZHocb/P4ay+YWziCHYAHK3f
KcUeehykuJLxCkinLkxTiPJJnvEwkBuKxFX/SB/RjnTS5OE04855h9t1Lh+9MYsPvkl+DFpMVlEL
fcbjgLBORGU2VeOc+a1NwWYNDDOn5H7PGY+jgyquO2nnxxZPNfFhw8sjgXbFqyMdi/3N71rnmc52
hfWgZviayPJ/zLR3sujj3Boq5LEm0deghEgnfv53xo+Kjh4ld65GPflZwR4ZHiOR38Qa5wY9fmJK
H0sFM01u3lM8/o1/Po6yEZ6Vt126nV6xfa8SjXcK+N8eBKleEOvKu2TXXf6C+JCbhTGhNnCQSZ2U
6dkcAbunY14/m23dSkqH8UQOaoZ7As3nbRGlNayELuQ+PXNhOEXIWv8hbg5vK7qdutuvMSrOt76P
GVJcHIpxoh8iCYjGNsoR7Zod4JM11oiWJ3vokcxFOYJPiBzhJpMwDUrJ88Mq+On97CeWHWWDNv0w
tdFD1SHQEwqdd2IDEqhtuBJyA7nPFueZEMaibLqWyQLzv3MW8HSoGOKdVi9J0/qEeIBVf88qAe5Y
pjN0PFot7QkXJoiQGskJGeBxiqUXdM7rfaFdNcLgU92weeHb4c+rTVXApimiFn0FEQIah770/eUT
LZZTNASL/ZNaVPfuDqKlCkItH+H7vaxW5LDY3YiWmdqhkpqECV7TususMiHUauoJOKGjlZRdY1TQ
eLUwO9xM3LaBJZQrIBeO+G6FL+98MFbGMDQDva62rwtudUZCES6JowCxCrxturVYl7ELcDoqOu8I
XufBuRjJBeetHVAaxTnrQIPyJnCmTEIe6zY4x3m43lAvYHPxUih5AOWpn1ADNcQi5XxswuPniTjK
gle8Bt4DB0kqCPh4vzXvPQs9xkCwm108Pu3heTe5SnrkSu/IGCD86j7cUYpBXJjPfMS+WC9OlmWS
2lClYzVLpHBP3bmd0rXnysBFQly9oGOohpx0RPAOfzcpwTgriDk/Ju1rAhp/k5Wpc5IRRi5lnkps
OOfcM0H8pZ70wM8iBO4DCFOCq2/b6A7OZwgVozaAOu7Q5bjMRDLjtiu2SY0nu/IzLE81jxFe3LPh
nDgBWKy+4IFeb34tv3DOrO5Uf189OsYCPb/zNI7HtUYnAAcxGUlwHGyL1S4/Iucs95edZn0j0mAW
+KHAH2RSUB45djTHT/80kUvrlGk90c5k4zeYjjplRevWAxy9KApfzQwf9qKwcV2Fq8IFGvepP132
+j8+uViLIU40oF75sVeFCc7Sg29AliArbSoI33m49QxInMBp9KHSB6zz4EBLmjixCyye9211h6TZ
z0KFp7NPxTyoTW/eYvmE0luCX5eaSCO+B4XsvpUP3fkBiKqUjAedBKorquEr9NxWTQtX+ySfRGUK
SBBLprivcIizAKqgihe+bbTp9h+R0Ago0yF8a8iFDat0l3PcclgIGzopgXjsz3Ml2kJiBVmdEqPX
IkN4GcvX2Ry9hDopvWFaNMxEOv79od5Xinq/b/EQ8CalUNrHpY8oAbREagsShpNH5XHbPxKTRy3y
rY6fJKNuC7dxijotQ5dmmFeiARzKkaTS7aTGCVzOAsRLg92E0q9eLxMA0DsHDCRVHgCzJXU/1we5
Mzi4sKj3gBc3rcXIm2O9yE8h1jKnkz0wMQEd+ZLC+3vQrjUyc++MD24mkZDYC87Htz3IiqRMb5Kt
0TNqnqujSrwvzsvE7t5tXIhWjECxd+banLVnw/EvA30EnaydgvvgXt2LlPPFyclCJ10O4iBGpq/r
HHkXjoWS2PrYbhW4UfccN/qRLhiwxWdxozwtA6c1jGKoglxohzOwUCl/i6MtC4bE+m5o7KbAbZSl
ZQzAX79Rl1qhaEL69DGHblAi7D7V81Jkv01VnS3bBvDVoRtHbk7BYMdumxGDLY2fC8Qij6kwmFd8
eO1dVRmEsoHlCz9bFQqs9NZKXR2ZYa6GCP6ijui0eY/xj8Jw5NViAfqIsagq4/KjXfQhYOTLX5jW
AtjCQEe4+JY2doDT55inkpUgHK9sm0m1WDsUaIq1YyrbPjBBj/e7/hjTZyeoXX3fdqQYvOxcBWOO
BkOgxqxdgU6n1E4tQFMjs6AKEXY13smlB7u+6C4mbOwPrAQb+3XUZjDnYwKGMGRDcXiJLU3uZ+tB
kGOyWuNQuZ4koR8sI/wIqCDKMiC8RtGClOgW3mFqaFJpdw7mHwk4Tcg9S4wx4yzlNpDXixOYWyTk
H+a4uG+PYacd2lJaBfc9eNt9HIFzuZdU7qNWwvNbbH2bsiyAWCYbm3E6YsRDEiUe3++0xIXIvWoA
qHC84PUrbbGfNHPwDKIk582JIJr+mttY537yirJMSZkBG+n4k9I8hjROxfdCjTU4DFhKq4qjD19c
5X/lTOuMHG461hKIEa30rtdlYdMK3Y3iBIg6YQ8tA/szu1cNymPCuPccdh81ejAo9fEl9xJZO1f7
Kd+xXYbQOcBxCypEy+KsYJPW3YpaA372SqldTu3CtVlpLlocuOntrJvnYl9oS5qBJukJTo880GKz
uQqeQ1MNiM9qp59JlPPyRR4cSfoOSgYOeaDvie/IWKLsl/DDR8DWTeUwH/hX8nsyrA1Xc9nVT55l
Hu/7HsUmQvKyjLRRERrzdxVWbVPrZtXWzK2ues9DQCGipf2cLsyor+Jh1zP2rOA+SEEOFizNU6jO
q+UTFXuOE4srcFy2Ul0sR84JCfVlggzU1esbhcGcRA9H66WFs3GFFvrYiH34hBsZzFKZ9qHXTCLB
nQc2Gaek1MKQqE0dlfGnnoDd7cgB9q/F4sOCFdZDjthPKcZNE5XYKfsjTsIDclS/PT9XhuCLTrex
+/dhPDKkLNtngJGJN2cRDTfYfKQA5rlCCrXiu36hy3T75XcUUfqxRMlmo9Z/JD69hJJbx23CDk5C
Xt6bhWfFiT47f285RXQvEZePygu4jVe/vXNhu4UJjkGVg8Xl3fAWSsAKfAuw/Ou7ofpmsX0Jyy0k
lrFeTE5LJugm4HKJlYPpV80K0PwFqXOwBvNyP2I/3BK1TIaJE3/+0nO2J0Jp7cHBGH5dzNnXsPGD
Ko9Vx+fjXdk7LEzJ9GGMAv/aW3N0DCh8nTeRQbekN8mwJJraBj4BlK7LzwSGqQe5GbrqHFjvwCWz
rJsfToErGLLzPAL3A7aL0NiMtVVBWWRHDKgjfCl4jZTOqy5mvn30suby5LltBfrBVnox5UDbS8yG
8cUFlZtMTknDCAN/99O4SjvX/ia2h7HLn547x1a4nprnYn9EKtjLgSPhLmWnWZKhzUGrN1wld4in
kil/ndLXdLmZBanOiFolN+KgBMrOIGHROJYijuLwAPN+juwvY1ZGLLhDHV3JLorVnQ71iV2q5txO
h1/wKR6ZNtb7BnSJbOHe/A1PenxRY9hAHstsLIO+gE94+E9YUYT0KjM+2MzqJHAW4zRsvKk+29wa
B6WBnY8P1gWYRlFMVRd2nZITkj0H8Mdj8MTiCb3jnFXcyR4BqLmHfIfm47Gk66A9K49Qnmz3R3oh
xrzHzAY8NlSMnk5aslQfwP9eE6y2hJ5hcGYrytutzh1ZWmQ0UcDNzEnuBpacpt+x0+FOgHAxjbGa
cUS2ZSpztBvu5h/f3UmhIASSnCvLm2PyZsI5HaEdSMMFcnzk/G6t1Gg9CEVGkg0+66cUUXIvA9+i
pPEd1UMokMJPu/jBydYGxezKgtdXDHxE0VhIxM/dmC1FM+5jx//GF+wX64h6/IlPJJbd8/nGH8PZ
RJ1rMdDpVV96dumQBR82LRvW/Mpi2/5EkfN627iDFRMqEpY6pug4aRvfGmbE6fwrSUfm56yEY2Mc
SC7r+Ew2lOH5WnjpPxETY39OU0Wt60bptIRtk15YmR5ys//V+vrB/XHi6iBLRUsFye+cXR96w2dP
oy6aFwFa/den6WgDXb0KyyfV0EjVgGlMOpn+fFf1qQW/Q2sYD8DeA0XIyGRKN0cBI44/Yn5g26oh
RL8B7c53uFJa/dsoQZLTfcCSgHIjGuEWp6B8xkvt2zSR0CnkHYwVrwcfvYLEyox/JYj5fkd1PqDj
n1BupnxZRNWmNV2sJ/Pxw7f8ByDfxKrNox4vvfUqJLbfz0ErUFiInvMtuvZyZJaElS+gUhiQEbyJ
rFCJziXjrxRB1DK1iWQk1jPhn8HYnilhkjnX/SrF/X9totPzKlwF8iLEAt3WZO0t9+Zj6ABehgT7
SVq5JVUQUOmjWlRLRcDvcQZIOLsR7kOnLKRM3mYYTqstlPIY4W8FR3hoRaUEF2nwYJJ67FVEnd4L
diADRN5jGg28+YM3aYHntc387nrdzAdH0vpAUobNQj7Km9DA/HM/UahVSoDtifau40S6jcbVj7AW
ZTixneNhoDnSRb4joUpT3o6Xk+Zehhr/yl0VLguvMn2CfSvbRzsoqC8tQV3Opu2m3mpo5D/AdqBk
zkavXMJDD7UiJZE4ey+EZyy12MaNDqjNJg5Dx0IvKUA3xt5nb6NIEBCh8+MqPFxooK9Q7CMLHqK+
benzESfMXUJGgJpKMC6/l5qPYWU1p+zCkOV+PxmKayxD5WLiqbXGQcQm0U+ybt4mLYngWQJxc/eE
lM2DGWfcTFfU//sG5D9wrJTjT//tUetfLgp+mwGqzv5wwuV50siGjDlQVqo5HqZl75vY+dC5aXSI
cyqhN+Qc9PwmfYXaPRaoKUwxhPS5em2g0fBZJfPL2Kw7DCkju8JUBBYDuw5s5E7tpB9as2+bBu3B
2aHNApD6E2xhYJNZoJ7CRraJkvP2HvFRMb1J5NYiSrsdFxH8rOzJwN3td6w0NbEsO8BHK25341I0
y9CE9w6TGGGoTKuvPm1j8VfOsrPFlIgH8La6syexNVgJdyD5qaWCipN9tiXsvRMxpgBOTbLSXZ09
MCxW8ORE5OodTLxBsGpzc263PvXuVT9sSBATyhvfKkN01PlufRbSXE5wvdFUnUVp8zwjueUiqPGO
IPU+g0erwDH5nTe76YjWLuqZ+DfWDlqG99NIjgoElFQKPksvbEjxp8wtysIlKyuRBKHbdiZfZS6r
tl/Oik9CH9/l+YTGKOSW6xko3xlC1BqPVVPwrHSluG6ffu9Vs1AunxXYYfgyix2ddbIvbBZSb4lz
jhIUhWmRXvvzpK6lG75Z2Bb4fUYYJ49CPtq6DxaMYX0bp7yPEh84Qqtm8mjN5SbduUg5N4bxCiDj
ZLr1o4tPB1175ugNUU7NSdnrhZTz4dEzXo52KcPhBlohx9c91jzJSTY4Z5x9IW1a4UEY6Y3BIxEb
NEAQoKW8Rkf5zXcdIgbazbt0+iAbuZ3gR8AF4yyGQuH8x0tvqtvYZUShkNIAQ6V/O08POwUyCOd0
vZMIgGxzo/7+W7GI1/qPa+027dUmKcAYruQhuKMPVqSWjorQYbsdVeIe59UtmDNdc+O/Y3ZriLpA
9H3VLH2hEU9AAu1NcxWnAk7tq2xIbVlkm1OrQRFPcgQYLmUmpfdvbsUCM3fgeWhIGNd2nP3IxWpT
9gb2KUVh/JLiAXaQEVhM8qOe15PFedfUz9kIpc8PnWsBGxARNIOAht6mnxcljxRbITMBwcwnr2fY
9zJAh+Lc1/qI3+lhXI8h8CmqaxMyTPGXyBxNz+3HQep6NiMDV5cUQd/APqtb7kydWDgUOH2KM0lV
idlBxsy9lCz1EGvIhygLWQ1asFtzKgMQep76bqeprhkY30xBrGS/JZ+aW9K/PS3guu7hL9vpyFR7
kl4xc13SuwvI1pY2Jxvv8JSDFT+rWJSdteel0VvDyARaOE5f3w2gDSnjWPuMYXEJ+/yNLXrqIWNO
dwQoIEoI9ZIEKTJOBqPs8GxhqVaeiTXA1Fb4SOJBRJW4Y0vm/jjzyFPoQOvIaKg/KX/YXhXgtlcR
GR7NVTh5xnmgRIQzqlsdI7E75/dKJAfeyKZsuugK8ooTx2Z0SDLQf4aqqz9XhvtTZG6Pw07qWTYT
kFvN54C0Fj9Y+sPk5qvnAItwoeeelw3Ok1N8P7SnugRSD23hXmJm3gp6vCzpXQ9uIcC3CZepa5QK
t0iXLvtDvo4H0WnN3M+QHmUO4a1frLbe7v4x3+VJSExfLEx9cdKR9POrpRR0/gg8ADyKN26CCNWT
GliyXih4RCZAogb6AA1mQB5JY8c13Bqefh2+G6/KgMqMFnMwd7P/HxSihyUUnZ0/lFYBc6C9ALLj
WhIoP74jlXqj4IXi6d5X2egADY1CcE8huwrHQK+TbAjQf1R50p5QsleeMq/HmGslZ3psEmWWPI6r
qpxjmCsQCWBHY6Gclcz1T3SbJDVBNDBy4c4/SYYe0fBisghQB+iFa27Yf9+hMLHI2ZcQS3vhpjm2
Fv1Pg5nZa+sg55cefWMUBnIZv//dk5dQ5bHweimRSSWvbqGK+K/zVQrnNMrb1+oBawGF6+DtvrV1
0xZQPp7r8evjZQNnW7stGmBreJ7Bo7eye2I1QfGDtJMxdUL2/8i7u2YJSiTkTFPMxvpfS573MYGC
SA3E/arERBXwrBOglfHO3RKmPhHB4XhRIk4N1hFS1ZOsBNYJBWyY1JCrUZ1EoVpaGYoAFzd+C655
P+NMVKtEHDEQ7kpu+KmO+SNTmXe215hvNaj9axtK7cm/cwRV2KZ1zMnuQYStykqygS2fvGdjOJd9
9Nloi/8q0XrmIadU7TXiHJFQO+lBFhLlGErXXQMhpRuy/NELKvQqUz326Niol+dcLtArR4EDmWrL
O09UgRl9VF8vdtpCBEjnCHyG6uUldbQmkUJFPqcTonDrLABDA9dsjdYz0Fiw4/cnSUEMMpavc2Kt
QGUF5FRWPsK+Ut/gJdEyItbu9iDRHHU79xcnxqTtIEtzxFRTnwhxVvHAKlbuxpSDoXIe7g3h4iTj
HgEL5RwrNtycRzF40Pg1DcdsoIlhqJ/aud2cTAz+ss+YSF8PAPtuZC6uShM8ZwhzRCVdrCyySRyq
tfmYN6IJqdNqaHNUsc0alGuK+1D0OnGTllvCv7J2jGlLw3h9SlyU7M3oFLlpYtlOfyFLRnbTWCbc
ZBXaxSUbYLDnseCGilq/6TRgnCVg7YvdwKhSuopXe+Hn0QwgMX1W5mqrWvv9N3XkJxgi+MwVmErV
TBlZoODJ+BAnll133lftQL01kF0/5fC9GhYDYriPcQd3dekJfFNTvoX1Hr0YtRy5YWmF3THZETQ4
jMHKIUZMRu5APMxnIXFL8f4OL8PBzpt5vQf8Ik9ifAdtdTjh3txht0U8L5aMzcYWPjSqf/RcjJDG
Z9PpkOaJDYOO0CF3CFLpTmDEcwtGnW2gLtjljK7L9AvUngcs6Lf/dviOOuSzyym1zKurQaBVnqna
wVlFEDpDrGjwZlSLWygbV4UZ9ni1yfwmeaqlDFThmyt+Yy2LRs+cN1MGRZBjT04mfA/0xG88Ujr6
bH0aNhI8youW7O1zfySWamBDS1Y0VHsT0iJBsnKgeLXyyjCrJAznyuSQnNFZeBLKfNJfpYwjBprL
bfL7UFJf87yNQ9y81FoZy5f9kzGy0J4z3Bkh37EjDcglxrcfikbJrBeCpG3oCBBm1QDrXgvDx7Sw
lx2H9RRX/irugMMwbdzxk8td6kszsXvFW7CdcH8Z9Gu3rlMpvhDPOYym6karaINQhaWA0+4PzUx2
vGMjVVQFQnKDmM4XLqLA3aiPWfVBFjWo349uYRO2SajayWPwcaCts1qDXn2ivBSaGaxHAkPyrIAI
REnFC0nj7pq64Nd5StdovzHN8eR1fZFW4JzHqbs6Gbk4Go5KeHZ08QmvIgGI1STTwKX/QlKupCup
0EQ4SeTKBIaq4FcTnrCf2796XQtqWApKtK7C6/AOWOdexDXsu5Sq1/Vx9ojLfRaBTD4zcocmRa3g
sDw9DqBhKxiuqOiTtv8tVzB4J9m2kiSkQnd/n8i9RUAHYctDjgpCwJSvS6Tu6+IzINl0GPOPz4Pj
1VvF7B5F+XUYDBeRCvxUGucGnLw5ICXtHGn3PUluP3Bpti0WOw1hvZgf/ardlD71Z4pl1J9wd6s1
A72c9DFen3UwwlilniWvGjDeHj4IdePzaE5LQN/MaT4ahKZTBtFNfNiNytEIyC4ioLORhcJYQ1Zp
cNmk4vlhziqwTnRE4COeAcny86PmqP+sjmywzBEyy0u5kJxDgOBKBzAAgNO8FYZBuLgEShJl4gsA
yTTUcyBXpghMsSyejjNQU3tUDyrRzTDuCBUyfryHX7o7c+1eJpdFT2em/i+8K67P/oupnPNSMrjY
QG0YDBPUZNsP6iiNK5Z0YffRkww4QGCLNXLsSpbCMkWAqPRGtrY5LLaH/BFEGXsE1FW7MQDJkLRY
/f8c87ma6YQQ4VYdt3QIGbI3VUJIExlZUYqJdyDcKXo80FSiWv+cdXgWWGPIgPZuNqvP/0YCXcJb
DpWVCcV545TQ/mveZ8XBygDXVn2r3yYjuPWU+Gate6fh3jedM8wkKGL/hZD8SJmRF2wNqzCYpBYl
vkLvnS6qD+PB9JlJUo2QXxHnYdvOjTnWslMsbYjLEM1zXhgwTQwWQtV1xR+ZmnK6vVtXnyDN9nf3
4Z7EgsqXZ/gHzRsf+QVmDvg08yEze3S/dg8PPv4Cng9iZZWBeuwysM3ST+nG+33wGtJm8NgC6bH9
Y2KVR09QF5NpE1dcHczy9d/mrwGgl1dS15NYGtmDAc0MHb3/WweYPR6A3MkRxGfkY27adSVsNYLH
YIOowuIg7L2apywEs/G7V3a0XcM4d6kQt5E43pebiR1KZDmkHQQK2KNFe0PRBT5LY0bS5WLVxA43
ch7j4L47x2y2wz7DQrD6aB3jaIk1NoCeUBNf75d8fjRX0iSAVpzUNU7L4fAmei+/suulygwzoMbG
hYhOo3RuYXz3ILekG4KKwD+n+F0uA+M1l2DgM2ni5DshgIDqvyGCUncI5VqBwWhfo6FsSqycmz6B
2/L36ToOJLBnaV7c8E2eQdTru9QkCIj1tvqM14LbbggGET9Y4NDuWuDDUKldbTBeEIrhKXZsXrBj
6mJzG06IqHEbkymCWjucDQCGXjUcHskJB6qg7JzqSaDuO5HvtJvHahvLYMN4AgnI8NnS02ZB+P5f
mTTwlpKM1dUJz+2eguACQiGPhqdInk7BhdWcvtxtjbPje78nbuEU8HDFFMnJ+SxXQy2CshBd+QV8
VziObYEVf18eTtPrrZRZt1AUokPWHxWDAohZITMRW7SJddP3zAOVBXbwSZSpO2y4Vpr4wHOm87qY
i+hZ3kGIVllPrpEQtRfw+WTw25ppAc3FcXkXrQYv9LSblRIsCdQqhMMSTWxp7a+DFILP45A0GfvU
/FiL/DQra8+p+C4C2fv4Zdu5VafegT3HK49PEV+4Amz+0lMwwddHm4KHvAJAH6E5guMCT+/DYsTF
W42bJ8+OmOxSXwt4Abygva2DXf9AH4/dDnCmg6nKdNjMBJ7Wf6wDZdOzEKjB0wqznK53qsxxiBKc
uYB1qkugEU+BWNe+gH4zon3botXL86JQ/mGJhXMzgRsSKNidndDLeuo2/DmnN7HVpWCZsPUzGo1K
YyTl2a40dvKp4yR4hKS8VoH8P24+cviRpw/G2yjWI739AZ1Y6hb7wY6w7jsQkXkM/RsGoB7IYaMI
6Rdh9kLDc7vnTtnI7839k73buea+cWAsAXsdLhCaM462mc//0CS4Gnm8lxTu0l6fYLLDEx1CFBtT
eMiKHpnXIIK/AseGGgCfZAl2OovAw2VBBupihSQa3H03B0Gk4I2PLItkdDSMrACHKEiCjj4/yByk
KlD3i4LlseiTKUXFByICc8cAF9t5S9sKx7Qp+jmPye1dusWAqoa5/gBdCG4xwR7MZNjBQszDL8lK
1vphKlYc33HENv+0O+PYL6J2qGpFyZd46FkUUnbhg77pNMhlfPP14mhZwgPefteE8NRsHc52YvGT
neTTyoDuJOI6cnKKoUHgNnicngOzeXl3h5bpo3sGrxsLTkp/KWBzFnTuFi3owUTvM+UEnNPWMAVi
39fJuNNs+fg/XnBJIBYgp3/NwmKVihVgDJYIQJzCYu6hMSMqYPjig7VzRjASP0svU+/VKnB6nWLZ
0U6AX42+vqaF3dB/sFBxly2jlONtNefvRUh6pjI4I+4i2DzMw05A8Zn3lmcbRw0gBORSuqVCdVHu
6XXlINZLFOJUwH5E/+yeXoJNbi2LEKlYim6qiO2D/seVeoUDzvunulAO2L9Z/1oFBsEG0iCyLVIa
XIpF2RjAp3ERPtoPoEgRy+lulBTkCmjAHUezJJKB0xgtjaVt76njO/HVgPWRmUKkvDD4pp1Hc0ep
g2zs7Blx/7X47ggHoguJBOHRd+QOYmQxjtB9ULFtv3gnjst1V2ZtiaCkszxrCXJjkxZZ8UNz8pOY
6oFkqo+hEFjuXLgs2N7v7i93bh4nsh8AjasN8qe3Vn8lft+Ar+TmR58UKeyEWsflUKXQd0DgDtUe
RAcD6XuVuKa9oxOrVLk7dMastikkHtOYgGe+7X+F9u7+F2s4tFvECuLDZGZF16Ow2XzxVAp/Pha9
c6dcYn95bKQyvOQ9BmxtAu6xw+xuzNnbK3ekjs/pehtbTITmak0B6zHEzjQV8mHsRqloFE7PXq6q
U5iF+vn1P1VEfOr1/pvtoDXYZhm0h2EWaG6cdvlQRFvKc3qDzXK+RiUdkhZdaYgxbWsDKI/0gGOu
FYxNbuxBv2eRtPhhHN06p3jIoljZhAUySiU5yIBVLiFoqd32TFm+prLc1Dnvl3NuX11H6itzHfmM
B4V4GIDw6rCWcgezShs9yJNwDaxsQ85W5o+99F7nmP/0nA/qxFI7Iaxbym5hpQdjMMwebWEae+OK
SxZfv0oVDka0avkhlznIaMvWLuSwBx+ZX4nqStNj5TZ2vy/16irw78ra9J5ve6g5F5AMo+UdtGmS
E1x/NJrgQzYVswdOr8HRWvVKCfHaVbQNHnT8kBP7TTqpk6OgfDqVrc1ijs6wT5b0Sxgajip7Va28
C33wwO9tll73bQZTkpbzc1uldy5oFwdgEf0i5zCHRJqD+qvFi97nhMlH9tlQiQKbT/c0rq46Bc0J
xjD/wjSbq5aB8ZBCHXEKTkjXo0No/6rBpuQ+/jEY7y94sDwwRkKGdD76QpddxGPNoBNXUnGLCTAE
FPA29F98X1d0hq+OE/TeQSLDjYUOprBe6ajtgb50NghR5+DddSbk8UZJtH2hkm1GDC81bOQEFXRZ
GK3VObvCdxRsL86HDDXIBsf30ddfDM2pTrbH3w8BlT06aMr9WL/il+j7NgPzxgVV+zdh2UW3Evx3
SKaRIpGEiFpI4+mK4VApncXitpFbzYqR+nUN13yKMJuufN7bQd0+kmLcd0SYeXlCX6Zz/qOQOhAq
ylamPEwm7U6Q2VYK4OLQhoSI2ysGXz0tZck/5gTGlF6JE/L2T1tXlCitlTcAnmBvifdHdkurL0BP
lUNPnvbOUzq1ygFsxqpzaKzyE0O7eJbGeE7Ad6+fHRpt3CdoNgurhUfj2vcgfsJQ0WFTnmVUVlEV
5F38uOVp47TVVDDYi/LrelRT4dZgHfgThdET72KpL3NhO0yBibzP4rZ3wUKiAOIzm4jqOY9ZDPBV
e5FytN5w2wEuts6xsEr6DKJb+dpEbZSU0RT5fdPhsfdYeDL0vJS18cSQ3F+RWfo785WtDLCTeFT/
u3Dx9OAzG0P4cM+BbIs2rYlYaI32i/+j6LN44lgV7vYJnIIGtNpx5frIwyz7f69S2pVZDqEkQdtb
yXE3Knxn3L/Un/T1Ubn4XmWYabtxOG7IrBb/vXVeGWhD4Yhh90NbNvzd+LLAggD1dB2IkvFRJieb
KZ1MnBZUeNB/RfuqBMwS/GaTWSrhkHfkwB6AD52yt2zKfA3Pcx1oPuFgd3mCZ8lchiMgheRI2fzY
ioMEpm1F+4KID7nyhyStQCiOt7LdiMs2w+Fo83SGFtc6K5QjBz/CPvmorC20yIINYqPyNnkgDahn
sVXR6Qqh5G4XEeToWeMkWrmEzLMcvXQUxq5DUFHIy5jljU7/Yu/lxQ+7VcOWa7Vqx11rANP4IXaV
lgacEwYvwdlaJZ2lTFZsk4MkpghFzVDXV5Vl0Vp0M68uNp/5mfKHr+VtpK6mho3xlzheFr8Cy1YI
u6IeqgVq1XtzrFKIc9f/WYIr0EAhr28J1BkbUpPEorfxinRFWs3PJxZ9wooFpAQ818sxLcU672Qc
66JBiNOb6QiJxK2EGNBbt76EHFiu0wa85fd62ywEqcOjo2SUyvT8BIx0VvTKudftYhSJWcP1Psz1
lJPUa7Mu6rm0oIV4I8Bhh5TLGCdtjlyZPcLSAL4jbkYGi+cVb6bWremL6vaA1mAIhe3yuoIS2Bep
XycKu0oZp85QYqdoL+x5XsOjuwyff+cUTaS87q3951GPDq82Bx42DI9r0Vt5JPrUCYHEH+LhnLDa
IAbsI0iCBd6bB2YcyLb9Gf1Z4VEH1QEZRv4vfuEMqFJR4GzAEQV3yw+wR7pRnNrwd+JbGvJp816Z
xmZMSJf5JeeydMlK2sfSNEyfrGLXyEUBhkwmM3G2XIh77Kh/RBPOkJ4YAZ62t8liFvn0i+i5yZGs
8JLviDR8kOgM68DBv2Z5r5mPYehRBvhKFZDZsCf8N0Zuja4n0gpYXo2pIlrhjg7244KP5U3WFU1C
N5r/cq61eWwpd+LN+Ffqclw+6q/6jzB7Dlnomuomo7BqQaMHCPYl2WrTVa8KQ3ue41ln/2BbPCRm
cQAdfP4ybT7dNkopDr/IeAqBXIk3aTcYVMWL/gNtxGVEzh0V9W7L8J7TQE8c1D/YnZ4nivFKpgon
N0cuBJRmiwz3300Hln39PkOULeBXkYA92ZtFRCRVxT5j8h7xPUTcRpXtCqeBfgLAeCNDMKYCaLGr
9hxuKUYyNckau2u9IZ+6IbjZXn8sNDycIDMa9X6kvp+yR/qQIgL3N7GZbmUz02ozTf+QsFnOkGYR
t3IXmwAtdKzq2CIk1ssSc/AdWwRMie5gZBr+U967AocqFTn/0EoMY5ckq7qNyuDUbtvdmJsJ3b56
loxKBBJfY3xS7tfH06rveWwEeTKE4j8JzY0+rLSDOulYc97uj4cDpBgRil8xEfhEM6mhE07i2Lln
DVGpqdCijr6ovEsHuQ/pXZIGBXX+zCWbvfXgK6tf0FPBJsfbvYfBZCMyB1LU7/8SkDnkokbUYR+o
WcSRPk+bchMcEa6vsi29af4aKi8twZx5GDh6IHAl7wW2yzGVI1SpAuO8IQzjyBgX2ZluTGmzXN8+
X8Wcn7hbisUtAf/mMCLfyngB+3XsHTSvTeTgjooIFYliYlsLCUFC9Q94BkWGfnIWBiq0IAgeeDRK
d+jsS6rfr2EtUUCjKLQLrsC8zJJpT4hx9xoJcV8RSevUWIzjjgtXyXxILbP0brL4PtbmPMQ9koQ+
CsH0piPzQ6MXKLsaOIRSH/wXc0M7HR/jRCIe/a9USNb1eLAxfkztrFdnkSwOxP+dL1aJ8cADwBeu
JGCf9x5ZCADiwWabYLTZUl+oJJBBRWJAjES/fMY7YOQ4yB/h+prqDN+O2tAG/aQP60IiaF5Db3Hy
yOxdLe4AN32HA5Eopi82RnWl122TIpxICD0hqsu7bbaKfgx++CCNQTgkmnG4MqMXGi1mTzmSrMsN
F2B6APNRckfClcfzqtugeuARhzLC8fcsHlYPUj6m+vywyxoswbWUk6VegsTef8HukycvTC3DPf3J
7Jhl5d03Q0N03pQ+AtW10LSqCdR34LKTaBFnwUe8wmxSYbWwIMJvNMDegD04z6CFV3tedDMdt1/Q
wHcV8aG1enRQFCCuOrZUnPrX94BOvE4P92s9/BTqGObU4TRt+3fRziRcWtZfWkkXVhzH9UUgE2p7
58FDXSGccb4HegzR+LfqBXoKRwCD74jGOf7iVf8ELjSoBg5T3KpdbUt5hoFCu1YXj5ovBFUMYcfq
nPQ2cNJOPN9BEiELHXfLPqUBnuhQImDgEEzQd6DuNF9gXyGFomtodfZup2jwk93t7nW6oYMmNx2O
ldEIF2ELwIe5QTyCCKLmZT839NGbQcF6iINzsxZk98RN9RI5Ib9wslf005PvryKYoCUo3ZjLRXIc
x8qEVxvsn9RhPplvjQAuMHSpl6y0zWvU09XvpJy/PLzcP+5DdNqLqL8igdxIK+Mh6t2P3FxCbz4G
9bK26AmRz9y9yFXK/WQCrYgx023ZpdG/zYgQubjJy5OpZdvcxfCESLtFxeSQuCIeniAJeaGlqqFu
6EKVv8+6MhyGXXLARiOewZqgEOo0fanJkpjO/xRuFPk5N4Pp5JuY8HXZ74c1UY/MKT3Yp+mrMgQi
DH2H4YPQPGn8UpMl9+jnLfkXoRwS9BsD9r03PeA/HG6F8dW9H8obxNxZ2kI47Q/c25j40R8u93db
cjy3IeNUpAjgPiiuDuwUoAixw8rmSZSQfTdSnpIJezJ3+j8gnqE406nZeOIbELy5mtrqUOywAdXB
BqrbmJBnWph7Z1qbmqjfpyDUzzEwjuFcOKJhNymprSFvkOm/W05umOEcB7uT0XCiNUXq6mUdOAO0
++3POSRGkb1G3fwbM7jqFbjdxwurrYwERgRPtd6LLbX5MPS2PyKuPq1U2TqoLh2Obtsdqd6m+fhG
ocg/Ze1khTkHf0MAFKYwd2xOAI/8/sGgQPvJERekaxmBDmxDq94eVku7uUHzT8NijiwCnbOFKxEd
oZA5V1gdypyAhXS5Nu/JbLdghHbfw2I9NGltL3mhO4AL/1y2qX9eZnSWdieFPtNISTayNKMeosvI
zoAnYx3+Rp4v8J9GJDFR7V8IzWO8y37wuWnTs7nYJmTZ7V0Up2BpUyZ4I0EKiHyTjtAMG3qHmx3j
JaPu8pIMpwfmEieRrbhUb5y7kf8+z5ivtDTan+rSpclLvvLrp40OqtzbPeLZwEXIATkFEzv6YVsU
p6wtvq3MGYtx4PbUuUdkgKqeAnNrOraKnhDdOzpvjfifZCiLebwRSELKqo08mLgS72gGqTg8ouao
TqV3ISC0xPrazOkuTuT8jLc3W3gPQNFJXo2DWIcKdxwvGn025+Vd3pDw9xOUgelQam5qYQYMAepg
ibXD8HDz6jVeNHvV/1fiWeDAi3d+LcaBOU0SSjmWUfYsg8GkKtD41l28PfSvgXHG9q9kXWWkcA0O
FDb5OyahsTM+r3Op2yOqHZJb9JjYkHZtmoxu4p8yZbsGqsIImiwlYEjPNrZRK/ZWM3sE3ewQwZqV
nIJQkL2hh7wGD+8gHgGMNwnKeCaJiRktjQzLjDI3zUbbmnsmfJE3WnekujKQTvtsm+v5eRb/vwPp
SbMzAtSCkj30N1tNykEH1GjQ4La5RPfjVz4Fx1uHOz+FlnvwohjtsUe+K0hTCCNQ7Vzzz2Elhpxq
uUo0SORdDzl6u74Kfdlq7fE0TlIiVSBjtLJbY2tiEvMfb7Npbw02X8h1pHkbzpRr1rp8/DNpCnWh
0TQBK50bKNxzdS+1pw+7C/Ofup6rlxB9ccU1r5OUey7MsLNmOUzuqK9E2A4/eIyNv4SiAfl+tY2K
VAZQ2OSlhriF2rtvSRfXG/9qx/VzhWezKaYUXmoAog7DX+86Hru9eQfm926s0YnZ/3y80UNNy401
3e0ZUcbDJ+BcCR0amOO99/i6pHgMIEKidpUU3ljgVI3QWtsXCorUKG4dibqQ5bZOA1CngdHg9pkR
wnxu5ZPdQUy3Tq+rmNnImf03ih0eN65goBJOilD10qv89k1BqWYov9NNDUtNZyaRbGnhyAFrdUWM
qIvYOvOTj0HMH3CCW0ZFH8RoVvWAAffN2o2KjY5z5VeuHqj4b8b8zqUX6kWaBTs5wKhzSf7DJV7e
TFTRu+5zzXbKTtzl6Gqw4BUQhFXOb94875OMV1a6CYYxIv8vSTF65o6/u4RXC2rzh85yHhmmUaDj
VP+xSAYW0j7XmN9ekehIC3pbdN2QSunyYc4WEGE59vYCo5fUV5tP7AIFYNo2t+xGWNBVHhOFoZW5
mBG0P636TsowUEHqZ9AF2FFS4Fm6/OPBOK/LYG36POkh5YQQkmMAKMnoYY1hWzoZMXttnX3YTr2r
MguJ12ig9/sQmBmMJ8vVXKnLZ6byubYdDx4pDuDuf0nYNrgLtE0lor4+rrXiZ5t1o56I1YNyKIwi
lS4F7EvyZKSaUYkDM+L02v9dc/8PNKHYZuBLbuJdZGJO9v3OXvrTrz8qdrOBBJGPArKsYje9wPpN
IBklivmvyN2bXb16hSqLTcrkjDgs8eqoluEsmXXKo7ZQPi/wROAI7AERJymOE7+UVbBW/NeWKLN1
VZ5+nW/GD5EVmGSwpNhyZC4jYHCiVKzamn8RW32jieeF0WVyTBu/CfXQ5wvpY0NME3FJmL3l0g3L
5VmhvUuddtYpnVCixm1p/m5C3W3JQ7MMVX5oOxlQYQU4TyWjpE/8bqQ48pLfV8j1vJnYH2iA89fU
edT22YJfqxJAFgTrvczihRunCcMX9vVmEH9s3+HaS96iDQz6InRDfY8Pe5O9gUFQiiyolKm/8Srd
2snEMLJgUp1EkFn2Yn4RpUO90QNaHTc/rSXoVVz6c0gwUgPacdiJCyvGSygglePiH4U/iYkvsB+X
J5xJWZL+hHIQTyVOd6it8IAd8y3hOAL1Eiok8DWwV7FwBJByq5HGLmWzpL7/JdyPA8ais5TmM9vQ
YtbFaY0/q7Ljshw+X7s9cXs33RXNh0l9/Qr3vXaT5IanSGvbSajNSeTa0djs0stkNlMsmHMQ9bd8
Zf3hHXkfQxMddqtaIAaKz81L8zJHQ6VAjSgiED1vTKHwdibs+WHaScNqA4OLZPDcuDYHVI4wyuBy
TmukFVB7TImmVnFndZd46178o4DbCPaNiAknZk3LC4z8eiK8vsJ8m7OIpvvjJ/E0f5eSZhPmkXcA
gyW5D/tq7t2dEHJLxmGNAW3FrNH1k2s3MAsQGzuIrUvOEmUnCJPcWN11XT2AbS0N1pGf5zW3sqoO
I3fC+rVfZLJTjDRliP8cO3NBYA78xGNWpbJEQ/kdLkW1javJ4YVb18zw0ZgzlUsuWnf3n2y7/kDf
+p5iYKEC2hcyhxM36JIdMgthcDyvGckifsNvisT6VbzpP/n13S/KLpeBv5UMMGdLJIzKiScYtrgX
tNWsGQH7cykWLFymENG0ZALAdWeJiIU2O4g59ouMlbm5YCg0DR7eJLFc+2ZoX8uoR4/Z38wFz06D
o2wcs/OCYRqIz4hTJke/oF9vb1dKTAilqxiwYYg9OQcQcKxH4jo/uoT7O88+YgfFCKKvCjR1HPP/
yaUM19uG8CHJ4pZrPuDx5K+aQtba2zzVKV99SQOm705ajY0TOmCYNKEtv+FazgE6IQSOkDpTIPbm
5sO/qMr1asN5Uuvrj5Ngys+lL1/nOTmx9VtRrjXLkeGL4PcKEaPa0D4XqQJzgammXMZGItvbqfQG
nwDjFZxitFqP0rG62H9nS9vToT4yhtMsDObzNLQCDxj/q+th4+Akb+aHsE0qN5eJfC32Mx79m61h
rmO0AX/Q0V3h+gniZ2rmPik7uOl2uUJphCuNwpW10BmA2zI1HN1cChdf9CeutwVFuAyeg3dVkWJp
S2yKLn//4Z1F1yTNiltt+uCzwrAg/zmXezwWTN2Ds+X6aQawKCcSCQJAZuf5CXcapk9eXdus7uUK
QCeax2b3z1JFFr5sdIH6o2F4VM58ZPDc78g6g7I9ubvVGJWpfoE/gRczRNqcCB4X7SepzoBRumQt
/xyAUqNRIdrT41Tjy7uVqLZzPghhWtwatKq1Xu4ik+XWyHu+N/0W8OgBv3mzlODeeUamGNUBSywP
/Py0NrFxQdl61YbN9cnZ2jPGdw6/Povz/neOWGhVEP9BSVFmi161A3qZ4c0ObtS8YhzHUqS6DAV4
lIkpfuwb5JTvA//HOP7rD9TnscEt3MUTkd1HdK+jMDSVhudjQoGziyuhq7O4iBcFOev77V7f/gC2
4QYTyJD4gbpG3SfEKLbQpHIMc+La+PQRold9J1jKvpW1JzQKtx+daHVGCce4uHgV0VtiN9zBt0xg
Kxwlw4BUT70LEH2cY+YNSoP2A9/a6YQ+ha9lJcALP84a/ooBjHKTDSPJ4v4T9OZIJebuBzkD+saZ
AmggcWB5mQF10C4UiAdke0XpUD+ibeIOdRddzGXFAI0WpVrXwSKKJcK/u4qHOtob5dLBZpsjvXOu
NuvJxditgUJj1KA7xLKV8xo0MnefB4gXg7YfioNb0V6BRJCiyUx8ZHt854bzjKL80+NgZ8TsGm48
krrRLpusNnY9wQQuws4vVrKwxoz5LZXqjUfeqvEY5jHQbAwCFj3hkYYeMyLphAn0DjQ3zXIWKe2/
zNw3qZPKzk1lg1JCxhhfCZebh8OQxZsiINkD+kMTgv1f0S80H9juiEHwgk6GSc+r1IApxGtI8nne
IGivHmC0wj0/8taxvHuVLjZOEsVCL9R6DnhVdSQsUo260zEEgFRpePmuRVFvGNDjMTfO7fPcYLGZ
nn3lYSXIHz5kZc5XKR8VKzW8I/Cqt5W9mCPtv+N8u/9pice9WhRyeZKGReEaOJH4sIK7qr7K+IxX
fJaT4fkXbDhBdB28dGevyliV7FX5qslEzohORZzt+giz/updEdp35NvIGwvzj5KIqA/pgamhrJ25
pP6kh3VFEAftn4X32aguqjIGVtcZJYc9dYvWk0b/GGxlj1PKktz4JTIYEJ9IDQh6ql6S1o+veFWI
+HBnLCFw1AsxkF40xstysuJ+WQ4EX6OHLPmcPRqFcrhy8rMEt7/Ko6FtTm5wSv3hbMiLMVwkxMuc
YdlN0oedkC2tUWlcBLb1WgCZmpNlIfLhbXtldwYjzOeL0vNlDzWE4/LLx6ossxTRqOsYXQjWMsvB
5HfXj1mfxURCh/bnktLL6wvuSGGgzdGxC3wW2EmDSlkWOOmv2MJRFCW8nD/430XfynQBCe3DcTYC
dQmPUoTTxovBxHnqfxo0bUVtgPmnLSa0Z6XAh7kv+xYHkWMfMPiLF8ud0FvdHfEkBrakYWBfcSG7
MYm5bHdRCkxLnHx1pZGdNTEkvAMtTMDoYc0/G5OmZ41WEh5bOlo/S4aBVKZszfXuCqGMjm7+kclw
TWA/DXqff8yJWUwOUdapD+RAk2iSmgN1NPizlwqY+l1Hxr+MjejglyYpLveyn9vcUwSa2nl2AORo
sfJILY70qKHq5kWNqpFrbV94DQbUE8TvAJdDDN9Ae/J0idPwNp9hN9zYcVHEbLhCxXD5OlsqjTF4
+ACRJ66QbqdRrYuHdUv5y2UhkbSc6tPRQdY+DoZ6k6OV+wsG62lbXsrEr+P+5URBqk1wXNrlgT5G
fuwCsFpOIwQfRjBbCce9arEozUSlpPsVuphOELEWIOmCkKFFsakoT51zAZCdo5eoofk/Qt6nnD3h
sHSILlkv0zkE/nfPcT8jKByQijE4ijjHo5bOl25RXKAtznKNxZHGhARdF0/gixTxm5NF2WSR2GYI
cBq64OYbvK4HZ07GHnx1kKYOAN7Gv9TviyKsteECkQBnOz6b9B76uMPYjgynDpp0O28dgTqgP4+n
T8rXY1OvxJKQPkVnzFYpFw3BjrLRuSdTU2vYT3G7vh0zvcAJiizCp/Ij9P/ORjqdPDaCG2vMt93f
VmwaJ5oTzHqlkgtm5f2AAGGHK6YqITsNb8XD9EcXlGP0D//S94/nNXe8aTFguoHCnOSGq+YvCDDW
XGFPZPyWs+XHXtdfaTBpe26xe7Rafo0tCS5P82DAJlDaO4rkUt124gd1LS0dIMxTl45hOVT8n9zV
+OtrjLqpILEZjULPYN8wSXhT7A/JdyWNKzp1iHfdW96FfO2TKmlJyofxvz1hDxSWpN6OQKtEAyrS
F2CS77npdjaD20e8ayAkIQBJKhKuIKUN8v8xSqEtsH2hZVte7tdh8fa/Ny57mWYICWMFkMda3tSD
Eo5uH1F/2GVGSPF+5aUuJTjMCOEkh1yCvfE9hj2o0HJ+a3p0iWhrTizxs0jExlGobTeWt5QqZcnw
TlCVL1rbjVDQIK56frxf7kVQ/qhEJj41XjaXYkFYkDVBwPkgGdfz82Jpr5/GDyjC+tANrmXE1LKB
QaXv2n7eP+jJDStEWpJClLmRvUr7olqempI8DeaDkpimD66AAGv/R1jUFyUwezDrRx9+ItQWboip
CmND2fVzanOQXdd2ZCj0vfUMZS67D1udn4kdMxvXNUFgJNZkvdqJE5yYZ5zbEAdwe1gOWGqZ/7Vv
/YwynBKPrfJo3+BPYItcXrj/DA41YJED/exu+rdMhMgoMDpQ2CzQnDZZG8Z6+ba6zI7w0eDZ0LBW
kq6eBLXWEDg2THC7mPkHAixBAxHpd0Jh6bm23XE+Fw4h0Zzy+l/KExqNF5y5OPDxP9jk/3Tqej33
MfJlAp2FvvAXFsssEC2JibLvW+h/pFStkLWFEKcxMJTtzVPchMpytZV8+3cN0BB0U4bVmP1mzCwN
HzST4KpwhYJRARmhvhd5vMPM81eDbQoAKJVquhpVgFsBgbATT3NJPcVX+YhTzsjCmM0pIuA9dPqY
3snsPgyVwUpevP7u5lklP3e3C8tpb9lxPQv/25JFcUSNHM1bSl98XdprXXyI1Ntll8H8sw1NwMRO
ndCXcp6rmjHQ5v+zx4PXlcmqjrFVX4Vhv9Cqf5UJsZ9XWcLNVAAQpfEYW2bHS6Tn4ck9T05mbgIi
3BF+8CHEm3YdwWgwExGTPcx37xmKw5AncofYEy4UBEk1hfJ+oB6CKMD7yqT4Hj1/pMb8AljzAJw+
5Bh2/bie56K29kI34XVphsvtm6rjMbKrU7AVx15Mt2O3E9LRyiZtcEUkRB9nVxeQgWFZXfyR1549
FCHI+wDb8/xcVKG3mnbQxBB1sPE0NK4l3h4pVkdKXss0ecnrmxfXnqXFantPhYZjgDXkY0JOobbp
6SEPg8Zb2SxPKe7o8y6kXSMej0ej4PKeWHEUwVtAKo3HgG8vG+yu2zdrCylMf86smyUQzt1qz3Wh
fnVxm/N0TSixBPPfxRWpXaVvQnWlpNZ5r/sMBdLcPR+bFMZjntNa8IffE+xKYMlOS72A/Zl8ybIu
MGFrgpP2DZ5XpYtjTNy2unTynwQ+JTvxnIrBt/+UoaSWLTXLen58zg2p60sPfn4UhTsms3jtj4kj
YN4xKWBmvl5E5ra5/Jt0QW0oLGRvkXykluv5mHLLNgD8SNVKg9Xb0KKOV2FnzHGNTUFwfDDXjgr+
lMDBPw3ju5ZYiAJwQ2RD3XV6iedycfyiLBMVOzBQQb9KiE3A/9fm6m+yfjVXWbn6JxdH3Uv8wPIM
qWEHnHQtUcgwKId/U6qpeoaeRjhZQXsqnPKfksOuZGiZrHgc7PG3QUE5vdktKxViywxmR8YuHqUQ
+avAh+vZAyws09hDnkLHs0CHiH7qTFhkz98OfxXD5HO1eFLgFsMWwQ0SgEJPX+ZBhbkRZw63lPeh
bTZ7hATGuih7YyH2oEXyBXHTG/01YDVQSYMQ3EGv5pq+WSKMOdK2C0Jtkdg54MyEvj2EhZGJZOdn
CfEEUL7Nf31u14Sqx2sA4SXQCV5sT9Q96p8u4hwRguiK8geK3/4TB4C7pWAmDsjg7QW7Uv0S/bY/
NK9VtL9lRDzF+7GjvJmZ5y/0DUXNYvwIeNoc5QqGqV2R5fosDzgGYOAEht5vjgGAD8jPeftQoPbw
Jb1SWrtfK87LXd9s0Z/jrkW8+Dy1QpXOiFtARh5PRS1Obg1BVRVqGgDmmFj3+OWYZpR/6pWepipD
7X5qqdh66D9f9U2A8UtarY48AqaxXNdlfF/gV44rIBt9pU5fpQW0t8gJ6ULVogyssN5xlRc/Eik0
IIhEmbWPdxcrBMHnWhMCtqTe52fpA5PrlWOIFm+jpiUTS80Fq0AzNXHqdewx4ieH4yWaeICLp+db
lCZQ6cCkiqydwEEMKZLX3VU7kX6Frkx+s/gpNFiItv0AN/Go+85dl7rJXQPDu7Q95pDPGkhaG+Y8
78qxawW7jg8s4c7jtBR4Dxq9qJWPVUZhD26qDA4hxuRMcIyfpJIVWhcN9TOi/5zxRnlZzpYI/vQr
nKCAIjQP1wmMipRdJwaPb2AP66J7Y7kHwlvI7sw/b7KwNC/JmfsU5IWj8gH5h5PsgmT6a/8DNK0j
xvGDPcZ7hXAi8E37C6ep1qbyqql8rsDlMtXmbUmR5nfW2QkRiOjhfuREAVgMGmD4mQrPezOHtUw1
LUviDMBSPV+NicAsCj0yuysRLByx22aitxj/IHO6UPvWAitncEwUAvmHxve1VP2spX/t2JppG4Lx
ELihZm6HHUYYrrf9w6sdQ5zTiQ9GqxXd8wy+sf82bQIqdXfmu5pGg0+4LGKaHTjLN04YOHzriyes
Ji6cy0DulIVIAvo1cJd3GSaG/Q5GM6T9CyaJV3OzJPogbT/AmQhsQhvpidIFdOvCzmB2KZvySXqR
IPt1JEhmc7J8cxrbk6pZwhX9/BaZfN3Xtvm5Cak/sLLYQM8s3ccbhfdRFKBsbZQ67Ze2CGKrZeFA
iKIUYG0mw/kFN2ucPAwHOimWRySw38RdAlepWNrlQpaW/ZeWjnSY5hTkoA6yXJXweCzqGVa6E0DS
ubrlHujb6LLceMMEMkTkp6MLqxEN7jM3t1sN6tOXz4nlE2WoS18HW31oMTPcMFMDmLi4h4BXw+CH
lTnt1V9I9AvuZqTG13fQ27AyypP+/eFJzIQm5qgYdzp6+b/ZKLu+9/gbdvjzB1JW0rNuk2Y/E20B
f0ZYi+uzSXuNH2NQIW5f/WlcTvAFZk328kze9BQiYbVa5zhl78WQqoip2Ohn6OWHP1DfOzbUXHTp
nSvPSAxL6WG9Uf7p4KfHquri+VWjmaXlaaXiBG9DvBAicE7DulExUoNy4HUd3C9om3y6z/r4R/Gj
Ab6xelaKbP5qOAigZhZikVqkuzxIaz0iNy+ulzg9Qq1D8tDDsPbtjErC1z2Igr79z4+d/sNX2h38
ksBZFAfmZbhjnTCkeOz/VsLBz5dyRoKMjJUpUbkXCs2Mi/pW5N/lp+Q2hXjYYix20Kw1pJVuDaTD
J/l4g6bvenDP0zb4h9TtqROLnR97E/5YsMYahUAgvLENABI/nE5p2msoG0L+mC9OBtueGjNw0jgl
VCmbOi7CM3M62jHZlw9z7AgM3e43sPD20o/I4unNPM167i8drogXWqy5SljN6PioJHDDp7ndqdFl
pU9LY2SJR2N9+PQYA3N/yBlHQ0njfTf4lVR8Lm0LOG4jQkB6ckIEYnRxqUJz0u29GaVwFq9lnQxg
6lxK6rgfyRmCcWrGlHiaB7f3fWeqmCmLjZa1V1iiDRD/JNlsMittXrdxSWIwfh88YAuxkk8yQ1S8
7GZwOBgHyvw4R9VokQlm2w42nxQ/NNYHReeu4ewotSd1lCTI8cGjvNCqX19SRYSVvEpj7a4wg04a
Od0G3ipYmFcQL9gc3nVjF9cbu2KxZEe41Ac4LoR9Q0aSXlR6AnOXOQUeLE2Q/NAIJMtZL44Adian
0YlyW3NJInpI4/dHVnANAZxT5mB083mWrR9bLUYw39suKqYeEohtP0Su3Nm1I4NCoGL2rmPVGiXH
bt7h7kH9XmLkz0n45VOwMGVZ6cdznYAtY+1dDLduFGbjh+p8YdK5xczIaK6zrndgPD7RKd3XhgBC
HNh34QPs7oomCsctLgpg7LaRZZPlzf7JgRqegXqjU0lzr5G4BJyUwgahCEXiwrmvQOmSWk0yMkCg
YdBSmq0+bjSFXNeFr5jDoda3U4hBA+/WBdT008sKdddnOmefdfn8EDsn2AM2kol+2ptasUhFKzUy
g1RHb69GhDj5Wtwq7/KBVqUsIAj+3eKmL/5paD6z+JdGkfwmdaECSewT04KI1wAZYY36NswjyTkc
M5Pqw2/lChuxfHlT2X9Mvc3ju5Jp7SkZqz5oDFTSS7TQKwQ+O7PJhtD4pEryo/vkB5p45xbd0TfI
zkehGAr4YlHRTy8UkDXdkBEC3pBluP1s+xNj5roN8A7dKXsbhH7PxZ/kBoTlgoFvgtRNN6plBLGp
QJwcfynyBkZOxGCPAyraUcKdjvYKQ6QY3apKdCcfznPds+xyNgvSCBG1ZSBLE+zGUfgDE2ZGcsrj
ewYzI4K5sPdHVIBZzayJ/miW2D89l3sS+h6+imn9SCqeKODNOhTtj0Gu1rOBLMa06AgWbIAXV9E0
RcSDinrtIqVqs9vDgpRnyUR6CL5VQ9b53ouFl9UoxBBXZvlUS+fOmw8zi8cY+QwnCZrnvWpkVGBv
YO4mjaRejuB/pZZaX2yYg+NO/DZB4zXjlp+b06+VTQbU8mETWU4IZ3DQ1UFM1A/uqC/DFQKArw/L
n/Nv9qKmQzdaYf0fOPP3Y5MrpgTV5SRxCbFKz9iaxPZi+sxlj4wUdVjyVk+/yvLJ+c7/3NCCpp0Q
qv14tF7W11W83jxmsKsjkjEIdfTjUCUwPbkEkqa593HdmrFzYUZ+x5ZhlsLAc/iLUCrdGrrx57F2
ZFH4KOl6PaK3PpQRrC5GnnKX2lcWlWs5sNWlGwSqYAvCd5VYTlmrn9GX5XByDFvLwYK1yJqoHVfv
jsJ7xVm7Ryo2Aj6+IQ0kr7MIVHjPcWfVJLNFYG3unEVKXG1ClN0+tdJBRGECvJOWmXBe0YFiFONr
8pdP/K2l6+pu0Uj1viQmnJVxAPrjnsXpfn+T+/r873aJ/4ndhoL4h/3LLg/qjjVb0sndfT7tvIY4
FFGKCM8vKcIkw8Cv21OIDAmegLLO1fIDVNUIhm2wIgT1EQojW3Z3X1byyGgGbG641kZDgoea5aYd
1NDkDW3i530U+Eo0q4Bhh4a8BJt7G3BwhYxgwEsUaxHXqGpYy5oH9i4MI4AGZVLUSNGrsU6BSlJm
fVemAlMVtZk7YnpNUwsYXMiqeFxBHw14ZfYmPxS2ix4YjRIzbBxgEVHvEbTqKO2Zx0dFwE3c5bk6
IuL5nIWogUz+n5o6OFW0XVrK+FtLV+I7KfTWdMasw1UUc7miUOzMZEOU5dvVIjl/OvVT9+jydq+p
utEAz2EuPe2D0/XQwg8hOwv42lHMjuTlIPmIUoncv+6f1M5ReHtErsNhpiaznU+6bCavhoc6fSjP
JUpBuLX34rarF0XrIo1ooU0Y15YE4XzvGP6ma+tB4sol73H2nrQOfIlI6CcDZfcqybzEXILJE/jK
VjjmD3Gv0gIWmuQkf8rvy0mA34ym1aHw9cRTT6aBiHRYHpMc/rKRebDIGEj8vseNvWFnszzC90EZ
WIPIoyG8gEnNNKXh7i9Gr0IMTA0Ly7fLMcMLdP6/S3Gcr/5Jq6b8Tjq7FrHv7ddnfIADezJRb+NQ
vtjMBPBqO7gtJVp/j2+ybF4Gf/3U9Iv9XDXniKbJ8wvJLlUrxZx7WOE36izowjqmPhBteBgg0TbF
9RsTrS+h7zWcA/IdcImWBCCR48q38TBvj1g3PPBl3kHNocns7Xnbgy803Hf7vorJ4DRM2LemomLo
cn5YOyDGFm0bKmP566sz+++4/lGZoYnQ3KUXl+fm/+oG12516DzZa8uoJddndpXRSrjgXs1ey8Ml
cWH0DZFUCQlOY06MMgqEREgMbpYbWMgH8TC1y0l+ZcMtKZX2EPNqFaUfnJl7w1ACQaVQHWCRZoya
8Pppi9UgnPLYw2f17mCYbjM2LeK82QJVMYZ1AuBQybPrrBajjBtaPtT3Kwt4DvpsCz1rmEz4oavA
aEblAZgRvr0gJxHJQHdfIdJZ4Pgg8XsgZJyqQdYu+2J+UJq3irqYZUPGQClEfhXaGvKc3wi9lS+O
ZKO7rKCNNBPUwhkDqYDMpCNXibnxI7DBP/+VLwpKIwKLB3rDjVU67Q8sNXdCyZ/ydVIv9py0W27A
PCHPKDCIP2ELg4pWChgGpUZ5p62rgaPzL6k1mlPMz/AqQJ5oaox1XTf4t7mGacef99NwKmLkzOwg
I5RIShnzljY9YIuCXUYRgPDEkd1j1wunuuyE0NUu6M8iSMiKt7MPSL2CwMQ8ikZVB1kHNHxfw3L5
+EmFXv2jb7KdJ03T6NCn+emJ4bBZqujs9me1LUmrDN3Pc8yUG+BNz54RdYuTFoPHxjHoq8eShhVH
oIR2upRNCanLc0wSxjzxJh8iF+oTEG01ffmxerLo23ujuhBQgZkfCamecaSh1Th/cxyQ84fcWYng
absNfpgGr+7BoVIz3olygH33quUKc2x2q2VwnBYyUEJVNf1caRlZPDnwpvipQnWH6jfD4af2cOpe
vlKlFdhLdlnT1B1Tjg/UNfvZc46wnCzqMuZeSUvhHetW9pboPY2A94jPUe6ZqxB06oqPOI28dQfH
frWzO29r72aGGM14AoYRdALtte/sp4kmkiXEX/y+W4x8pzW4JA/hELEBhbSHXmGHj7mhCMgOlO+l
XcfoAMkR62Oxbz5LUGRoOqA6iqfdktCgwaJ65LJrbEg96+rv36V1r6yCmBkhvrLJNWqglss5FCBh
vKeP9ixjYc0j+WihoAfiOa3RdWalan6+ozG7nZQvOYY8K4x8iBprnU1wZKwWQFQAgQdD3eEJpYI7
tKSfPfNj3Y5BYTuD8aCCfc8KvHCeWiZ8B1xFDcFv12oPoIDyc+c03mwVKSKuBBTSq/NGOVyO3WYs
GQ16NEtoUVz32QkjlzKWjTs7CEYkohwWI9WNqgP7TJrl5ltK161g/s84q36GRaUF0xq6UD5Q6a/e
OxQZG/L7YSQhfzSu+/1DSFldgDHCRUcGDIT/rPCCmn5lrSqT0o0PmIv9gv4lkaWmOLrlbd3F1xru
zAAxDaAYQYPKjLu39LZC83bHY9WvVLg6mE2+kk32YM984ohLMQNS+GHqLutEVnSAUv1yAagTeLdz
CLRA7AarJSyEIHyGAKQ8J7hmZdG5B5f7KuNCyvoVhenjORpItjqOny3IQhYA9U++T02HMaD/+Yv5
eqUaXpeonvvTqZu25Qqbxnz6YAojA4w8Qk7tSTYKe8Q0CKP75XpH3z6hhBQjm42JFpa4UPPaDe8z
SHDrOCRcEDIsLOypNAs7lxVzGZCzuygr5oGtQMYraQUvLYjRwd6kApT7xIowjjq4bjYgdk9EjgF0
5H/SetUT1d+07ECEswgn3uoWKg3IWdtqJgEVeb/d2haRY6oCjmIZr5av3Rk5RR7LteGFaUu+/nQA
L3rm+2YCRFhz8cpldpXfPfBi4Wt0VKC+GHUx0aZ3tnrOyBZGEwlUI+4+TOt4pAn6q6En4aKTPQHo
sM2mZOfk97cAk/XWW9Hj62ouvdTjL1yBOHuSa/AMVYx/JsWMugrIqmrqk2c0Cm9yfpGWGoIfDebB
5UkLkix5jhWBcLQ3IZaKZ4Qtf1jm8GtH8jjxJkz7gU3LngS+DufqYEl8oxktykVqbFj8jN2+kZJ5
zzwhaE/nUuB1NiLXczC2Ieb/E5HKiugiQKNHfxCjwB1+g8vuFdzcCPsVU2/pcTJAbtXlmNL/1evV
mzNpy2D17JuoeMhMW0i2jmPLaKMQQ5EqXIIwlirhmQCzzH5nkPagJDUQBZT+ZzVX/u4Kqice7fc8
Ib5g0kV7o/3XoctUdpTZu4du7YsVImlG0VQVPFiJgOFgyvRC0xMw16fB40IcKDZDKKcix5BBrYg9
MyPr91pPrN7hv22/7A//yarRaXEnPSoJPfy9g4ylXX9eNIWo3x4MNidhP0fNkvH9IKB9lTDobZ7z
vUzScCNfjF5RHRSjJoqZzj/6xb/Lxu0KL2pI+pMwFlSORWKL8k9TW3we9ylb4JtQ1Gq4dJpeGAhM
hMDxhJggxz40VVQOQrRxRb0oI4xCyqBaTxil4e6B6vpmvLod6TS7c4JDGjavvjy3U5GFr+KoekFE
vWFe9ZQtt5+HnsBhrSBWCkqV0hGRneQ7SaJUUwMLAuLrp0A1+SnRC9CW7KR3JXNbbN1qUb2Bv8NY
K+W3bJBUp705ICaFDK8CSVkeOZT3KbOp0/hGCoQhJkAc5gI9FxzX6/qlF2MqhbyGK5JtOPrR1FNC
pPktQvQOujJqlhIZBnFLvcCO3nko1TIQ5NcC+f6mFatb8R/sjzzR3eEjOuJvbEnJQLtoiAzwA7rV
kC7mc8u2WJm53POYybSiQr0T51lSgjX/heUmqDfClJgGmyKt4Rr61swnLC/SnAynm1fEkl7l8u4r
WmAK0xbGI0Irhzgw0nXW0zxLdy2svho9DcVT13lsHRm88ERheNNN/6xq8Q5XC357BmV2shMonBUq
fjdGHzdSkXn25bqmtFgE5VKGpBihzflWaBAURyo4M8a+8U8MUGdig/A+eBLJNlPKqUMOdvBG1glw
Ii3Z38f/e0ZtjxUWidM6+3SijvrbPascLhqO5MPYM+IfJTP5U/jUen5xvkVwnLVdxkTzUeRVQMO8
JboDoVDHBRmX85e5tEywhdw21kbwyKsRCcaw2ND/fNqrqnBi3oXZiHdQj7RjE0yfXyeNiLNxcXJj
g66HEVybcMtyqQRLvqaM/60u7ongSBSK0Oqbhyl3P/YMyEwjbGeA9B+TP/UXbge3j4Q47b8p4tu8
nIZ9t70jz88a0rv1/bdpR8UQLSJpNvjx1G982zDqnTKUWthXFneUZZwG8sxiGPxIm6jFkNc8EBMS
lsg0RAwPgpgkFFGrvn0SfUwcwMG5faSFUr+RX3K0xVykvNfFnaCqL53A3+CDbqvQPP//kCvhzz6p
mm1E2Z3jczXlVLuCHOHijHdXJouJCnkaeEnoLq94ei0Wl87CEGp+kpXvwsqiM3K7jhYv1p6X4Uzv
+bkZk5ooGEQdxF7pB+U2Z9TEy80rlrp8Hb/MuQNL25X0Ia2tCglXq4JSHT8N+B6ZRKvp8LYcRqK8
L5gqRokSETs7JdFE1bqLolLASbsCp49ilWqSIhy42PNPqZoK7R2pgwQ6ICDQmiPmzkzX6cR0XOfk
9aX13kxIVlJvWhC/AAwMJx7lUpcCr0aRwtVeAYHj0WThIOKQFp85n889a5zd2HTn/yeLOzdl6ZHN
vgo5X6lD5z7F8FxdOyFFpoIlwiVc/bStB78vcdvHnk72cl34SwMVddgw9WFlFaMYtTLDIFJtfbiS
4M9rSMp5OuIY9T3N61IGVvjOW99VRs7Gx2S+ACV0h8rHwIL55v7xSSTs76kt9JAD3CwcaTsurSPX
zJGA4QfExTWVcKOYnDwE4Uofl2NVfNPqb6eduJdS6P079Z0n6ZxkxbjZWV+0pd3M6GQfe7mLfMCb
N2bG3YzKii/7PSCtVGrT8uJpGlFm3tSnbcKktL7Mqiy7Sb8LcZDMG8TH5c40WAbXKDc4VOw6SOXd
dTq3mrFiSK3XeVSWbUaA3dvGpvrncyT9BERILzIbdzmYRr/d85F2ivrOsCrbWP0PdUcjxsT8pk7k
+V1fhI0wFFVYO9FHSDUc9644dVsUTHyieBFyaFCA2r/obHXHLgWHJZlMDCGKIMxTM1eb7kQCkn6h
W7847t0WG05IW2LxGjqJkYW+C6KXkl7IUzBswvhdVK19dZrMT17IfSlXmyOqvZT3pf3aOHQ0LKG3
21xslo1QEUu+slYlXLZhJTHFcXaxxkIGYZLwaAb3PTJS186LTv30IIQpadjfmwlsDht0hMPcpBUy
PmKGpZGGa9UHQMpFc3LYoFnJWi+pwPFKEbX9T3i0obnB/oc2C+oxnvkKCteOCak1mUqUIz6RMRaX
/DA3c95pBFh/QwbIynfqBI87RiXx/ggldEec3CHD1+Fu3Y53FcDh2Fu7wgSHq40xqr4wOyx3BX8D
pew4b92SRV+ilysbTLYqi2/Cgznj4EvP7XEM41tyU1nbI+tmfuyaxhhR1PeHOHMa430Krm2MPxZP
z1CJEdx9LxTPJflhDkNJmg5BUCCQ6ccsKYOfVNTNLbAISXk/bp/09uNwyoZWdbFeEQLAgONTH4OQ
2+ibj+0ZOHiTh24xJULwP+f6hfevwDIHCa2nPaBBaOmTG4viIiQE/DJhlYfPj924QqV1juok7mOl
KkSMiIq+2quVS3ZapwNg0h0r1Q955MyuXvxDGGs2kQvYysiwu8rmiuYYWqULulZzLTfVCp9AlN7d
BGbf8Ohexu6hz52zq0ymjSj/ISzfHcEvaQK3VZd2JFNyEcSVWsRrQRTxXB6uKX8ODf8fZB7Z40KF
ik12BoOIOkC1CXwsxTXSALSNtjqoDhHE8JlyQm6x/d9ZQknpAiHoSDdTyUErxiB5nRhrGLM5UtQM
hw/FYYIaRg8PiCcGD3l3F01n2BG3/DGujEpD4kjRqTf1ToMgdnQIZUkGnZ/utd7KqI3n8PEwp+2N
3R7+KFhtbLfsOLpQyr6ittPOh5uI4I0fZvvoArNagwMsJ/N8heVYST6f8ovBGcNivtpOupJ+KAH3
9yLBSAMNg2LDanmizc+zW09I8+pNk3Fd4qrcDyiaQQCeSzo20WINmYeBsKC+rWFvaQnNWkNl0iyA
mKG/uKF+vTLD10xw6GHuSR2y1/WSQ5EnUVrpjKKW5FpkBr5URScbhNL2AH9DjzwG0QK6UrfOCbWT
Q488CCqNZn9CtEr+VmF8DVgIgUDxpNkKMuY6Pdz9whXBQcXyTJrT7/0N+LZYZagDRibiFYxJKPUC
vLeaUth3Ez8rQ5YBU/TYHq99ccH+v4RrtSJChCwMQCyWa0eBw1Z4w5x2zXNFJtypM4XrAnU/AtF1
YI1TKo2PYyjm+FVwgkOUA0BJfDslOPA7UeN6I56r655nbb2FHFqRQo0pdzSw24FjoH98ImWqAEwR
2jRKJymk4ZwGWZqTd8PFrAoRHwVJ/SPWjq3SyMpVUnovq5DbDXFYq/g9v73llrCmly343rr2TpF2
fgQ/fkhTVzxcTkqr3bQ2/AXdvhd7jPASzNiorXE9JAe5OUke4yP+oY3IK6TRvqxHxNwwzlJatUTJ
wc523hUvHJQaKeapXVyMo7+N1+OMcHJXg0BqhilUSoa6tJ73wREQytWqrsB3GOLhh4mUOzm1dQc+
/H7JUA6cS8HP82uMBe3ERdXkE7vteb4s3Qc6bAZZct8XIghMihR3dKe0kEyJiaGCtWqtcNsBUSWp
pgMcJQaUqmB64qKLJkcvnGlJ16BDE+E4GizOuoj2qoL+00SXogIe7fdG7+KTS1zOzrxBa0kC/QTB
0Tl5jT3Fc5A6ElAxh7vXjj6CS3hM/diLpe4mkQl5xUl35+EBrNiP3sginV+Wtq0FBnVpAvaLoC3Y
VJzwxUfgDFG1ZvsDGI0avjDNyME1Xrs8DhyLacI5OyVrfMqwUOPVJvZj9g+3QSHIeHVTjw17Jhcc
Qk0lEKTVtzoIb8vhu92J6qnoHV2paQVCKEWLDJS2VSP6d/6REwCa/gCBWMzy0WEEtECBBACOTq4b
BL/TwhiW3C2CQXRg1omM73Vs2FQ546dD+ca53ROu2VCCncwq4s23Hs4m/vr49ZX6ModWplb1mrfI
NU3IdmJjPrDnOLZTkvsauNWEs8bSNuDipzERRM5SkrJDRNH3aKQO+DFot16x+2QdSzxguSRCvXum
Jpll/pZCSE9ey+JwDOKzZaH2zsRbiFSa6SsUKYVXw/7kvlK3g3aHxB98bk38hz6drCsxCMw2ZUrI
eBixzt0b5Iua+PjQt3AsjqWiO5lHU5VbmHstCPK11sExEOuctQ2zoTjapn2lWdpx6zJ3nlk9O3Qh
BsjpLXcvWKlEhyvQCZ8Co63ImpKf/U4eF7H9IeNKBCp2MxfcQEYxqO8up7MXZ16cSsKKOl7GFPVu
TYfKW1PjDkpI65oe/ui2qHzzq/rfRKmow7rjhUmg65ffBhXblRHTxtI/cE1wkeuvser5CPgVtPsM
7yHe/wa3ZVOYKpkWW5lCsuvY7zF6qrHSREdaiKuflzP1o9Dvz0JkGahGYJybxjCBY2LQ/kNKR7YG
Ts49/0A9lw+SzLfENnO02W4NG/qF8ON0XV6J0MdqL6YnBu/9kRrLWwdzDixlQtNRGtKtAWTU4HxO
N6HNNt9tJ4pH9piSU6HvUE0KSssAWHuwMYkDtkCAPaw9Ja8z9NFHLqAB5mMmJC7Cfxg7fhh4fRad
lyMVcLDe0GK1BkIbRi9npOmcYXvSOBJ9wS1dxoFB2SVCvCtapP8kF3eGsEKgs0GO/G1XQTE+eZGH
Mc/wKycU/bBKvYDPBlAfX/yyp7mQmAJo9pY8Q1X2ZO6aso5c1YIMslF+NxhUpciYC6rrI145NYp0
DY/sl4PRr2aKf1F6mTZf7ftT01aRDCmTB0kHejRtmG+aAIoow+OZg5VelUbHA7DW0Zgdyx7bov+D
TBg8IHDK1VpX8yQawv7a3Nh956ZHzS6uVg2PqBKcLt1YWo0S/xxT8IRK1C3+PE6orRtW3O7Wc5em
aUAWW9NUwEtLi2TKQujNoc5bwqgzc1uHKmmyLzyJ//qsjFr3c04C1BukCtO4TK6fbWw7V7OY7PoY
1SR2TD+Qev111rQu/ndAA1fakTY8XI3Ttd0dTLAXQSIDVzd77ZTr5YrjCye3eH/hZjjZATkOVx0K
zh7gKtiULWrw1RHx02g7mf1pK1fWSgo4qAgSTd+Zn2sHb+KJksJLtF7Oop+cjQj+oXqmOohp6kCs
zCE3vnk46EshJw9C33Fg2By/kdiLQZUv8Fjc0eOVmBg+RSgyozJfPrDJMQahUG3auh4bvQ2UXHPI
FsaWMt9//jjoFFqWL21D2btxlhHPbIjpCjSLseXEWebvHGebn0G+gM4SBZsTyWRMBymPOObOLXwn
HMCRNCzBtjH5VcSGYncJAE2pPQzVx7j3iZffzgAj2Qzz6/R5tUQLgTsrcOX11SpDmFyyU3OuagIZ
LHZoeFTdjGhDCVDUq8b0UQBDOWqskfm15G5d/IzV/w+IkYxBge/evVmWp75+k5+Kp4rEuK2a4zjS
cfzRVZBdgx8WZ55IEba5XzU1XpsiQIO5Cjx2gaPcH0hvIcg3YOBlSbRefRHPMnpNnuLoj3jJHCiO
FKbP1K+BrVtQU4ZNT/psQ1e1sZvX3U+bCiY4e1BrUEIZKrTxey3FNaBtHs8ndiuY1msJ9j1pIuMY
H2rbAcYajgdH+hRVinKu+zUFbu0O9uyUXC49jY8NtxrlBwMDWSeQyAgGoo/CJ0U8zoS+EpyW8O1C
jAbAmfq0Vt127Vuws+sbScFp8h8aRtbSpiPk3E+8Ecdvdm+FVv9R6aEbJL4uKgvHzyn4wFCNxteX
FH05eU35ed3AGkRii5U3mT5cmHdOoWe0+uvfNvo//dpE0AXAnAY9ACfdTtOGkOIsStwpZTqdwvhn
L06hK51V2wk3+do8SDmAtT2sdflux/I1WSDOj21MA50Od2W9RIQCylSziQ/Vxt/Q8gte1LD6/cgX
yxokl5bc9HIj3l3l7Zfde34axaqzLg0o8bL2QDFunmh+p2+6+Gsag0HKDEKQGqW7bFJIX8WBcGU4
iHQrQw7i+uqj4vTNrNA2NxhfqjaKB855QTbt1jnK5wPZ2rkjiMnKtsPLQXscYdy1KHMuQ9SMNCJf
8wvZ325HeSKwDp5hBA7o9coAgMUcTiTD06y9ZKExA1lBShBb+7uJJvvk+xtXscf2xg4WB1NiAHg/
blM+V5JjiwMMCd/KFCBwlYaNba74zqwEbVjHwybx57oywGRnIkVZP0jDz29xHuBsyemyv9omGn8c
B1ft/7WhmUb9fLEG+BJiU+tmEr/Z3L6zxCI1LUeHFi954UOksMOg/UvkRw7EMaH8yDlSYFga9Cts
T04HPM79FLICQtZWaoUP6+gASC9lvGFDr/Hm+XejUGGfIrrKDLzpIabi/q5b4IL5Jvp/6PLE5yQ9
CJnqfCtDeNZ7mnIJLhYy5PXY+hDtFe/Epnk+EUj6QLAxh3b8PKuRKMzm9K58sxQUm3ZdmTfJl9p3
jzSwvTVN923n+bHtwxhKRtKhsCLqxfjS2SlXprHopCLQbgiku+YbEEyYL4zDIAO2xNB2iqbQTYli
hB5kpVY5vUgNmAXA7J/ZFxHYxklsyS9TaxvFRjI0N+v+nu3W207iuNZDFeDMD2eyDuOPd7VTqwQ0
xZQYOvtDMEJRQJBCwCR3OSP0WZWtAQZX46bUG+VGnvUTcFMxq56Pt05kjUjg5k9LQ+g22e5aLuhd
aPurzvr5IFqWcKe/hZQOzm8FdyfoG+25vIpgMsOl1ql13Xss1DhedEiFI+scaDfPQ4RMbrQ3HeH5
fgbr0XaqckKq+5aLdcS7pWCSlXGCrWVatrfcsQtPRNdkzagkTKgv+JtALTEtQ7o1aygg2EHDsrcL
PWi0gceoRfVIxL/JKQcni0idfClWdv3W0C96x9V+Oz3DywY/vdKCiiF3KTieiZR3cBym8JRpj0qj
6pa6P0h2HLrNSzLfiQjS2I0omWkoBEb4PB0E3Lg8Ep0BDSIOFirS6RWuWQYZryPMtupnxmp8SHQN
sHI+bgQNrFaUojGQQsXxw4VK+5OB8RIcTPofH882OB3jYCh7lDactz4app3HYcxrpi5UHjj/Iu2K
5mWVModNLqwjY5wEKAbp/qDdScPQVhQ90X7D0kFSy2ejVuTc4bhD/e0jIh+XsLw2E53a34V2XTUF
zuyyaRnHbNhvdiBT19fMpfIjaB0ToagjgnchnDCjDRyojEdpSz65SYBqxu64jLN+ulR36dcDiTz/
yhRPiaG+lCB63N1GEm1/0HIOEsr1yEpNsX8le02LLSuVC0pTX+hgZSeIXvQfp0uETDCkAOd5w1if
l3Ig7zGAwZohqNKK6KQb1doPxvsGXwSqkjVOWg21Gi9de03vfconhduIg6cnWHFxNv7yvuWW5qf7
R6J4LWvJPFU3wqyV0L1AmXWbmLas50GhpUB4eBDI131IdkGeLTjltF06ZMK5Q3ka1uFNBjHVbylG
eBOB7JS8d8vF/Zir76KbTTBxMC0g9nKQb77QylAXVL+xSbleW91dVKY/JBbHpRjhLbBoEC3bmK1d
lRVfoSadL5WX7/Hp4J9ekXn1Wx4/iTx03cCgW1PBuOTdplK+w7E40gJd3NfbzL3xFdHKw+ysB274
IbSxD7jMYWNHaBRycSP+Ymo+EKXeyAGvp/glfqV0zWrs9JYAwihD1hFvvTMTcqN8lYk+jYFF8Tu2
Wbkkm7bcmc7vpGy5+bjkUX2yFpBc6y/9dJ69HeJlinuXENfjYGDoaJed63HbtQM8VuLAUzPen4v5
aoao53yEA+2CJDUrF1bAvbzKOIrDeLEnidJXFrZeYfTeUWdt8kHhveBKrM4CUsO6P7137pUP8vie
YcdscHzXmhvY1fi9KUiFI3PR407qvyy3aPz2Szinc5391Fvw41+OtuxZ92pyC16ApNdqKobmvBkQ
/dzi9yBJPam6ypSqJDHBymCo+KjvOni+y2ZediDdQQ95ltCXWdwYSUuUkkxFmCsRJLKYlfB3q0QO
o1vtDmCkAq0AS3DVy/CTdF1Qmy+JydggOaOYmFt0RxJb0Vtjb0O7QpqAkJKnkreXGxTsU7elbTcB
3hNbD9OwJdtLSmz4GDyh0r9+HfaYvqHOMDwMgZyWqCdwJoDfAGEdUgfL0vOlkNTnqTOD2W5CImcb
LwNCkmP//PxN/ljde1LKM55Kx71ip1IlsxRMsjJdrtg/srMVxdh74OFEKvmxiPHJoSLxYuR1TOjd
EUKZXOHVTFLO69Z1R9kVMICYva7si6ympR6e1Km9+fO6R7NaWkSdOQ3giZYLIcjsapER52t1BsEC
w2mxa3QWriCySMyaey2lFBo9FuHzwAU5TQfndkfBBH9JSLfpb/C4XHcVWcJmCdJEA+FF+QqM5HeP
mHs8SAT/iK7Jza817wNswCRwjk+zYuiokMg1RqtE8F6ZpV2rj246PORHlI8gGTFSTtxCwtMeSq5e
1zVHKb47IV0Li6hWV0mZE1CHLZuTliDu+nZ2vadtI0gvVdh8Gh5ijHtBBVhx7XYzrmXdyZqAuA9k
uh+64sFSYzY8M1i6/g1OJr9sriAiAH6VAt3uJrjJKJNVVv40pUTvpgBNY647jgV4S4v0C36CrJd8
BqJPw9jOejglGc10dlGI826TbuQ/c+eGMf6HDpMcZajTdbSpcKwTd/ZdVvhqRl3R+ZEVbpHm6jDU
L6Ws3KxiaU6S2W3+sloypmHioor5IJoJRqi7eI+vh5lUG17IrdAvscPEX4Hxtr3ePYpulKByw6dy
lTAMh0ch6gYksqQT7THN0U5TkA9yfdBAW3d6zcCmNNxQGuyD40P8OlIkgNB12hc9/EI6EhR4cOWx
ddynEKxPdRa77UfvzIQJnzlxR01oPgsfhBEld8g6q+idVXiGb06JiOgqiihsOaRGYhZyAoye+R9y
/s7KdfLUH5sbEaTFjffsvqCbXkL2NlmXdl77O+2GAfgNnMqaZWqdaa2/KKRKrm5KqvPO7LE4aw8+
xMcjdLKi7y4cqCv0kBU42zBmG2Wqxo1E1K9+OY15KZN6x0EllWCrah+4bY/leDd4TISL+7AZW1L1
QGAouwbY9sw3GpdLcBtGPaDSTRKSqKezCdZsxIuOnnkFMfWy6isBzqQ5TVxpkxYeqBrLpU3DZmEB
eba1JQjHT0qQYNmuzI4125/cGbtFoQQlAjRw+9Msx2Fb3THEUWgHNQ1yT6BgHT9CdCALF+vbQrUV
BEpZCXFWASGc1YtckukGyI52MYzmqVuDnDCVfdTM3X0jVDv8SXLrku6fiBU2ieakvoylmRe4ld6Q
T2noEHFEslYXQrzcAvdSGfY4oDwk50BDeN6+SPtKrPT8sphHU2Am0Auo3N//U2NHRHE+MdOCRstY
zybbQ4N4kPc5pdeElTQXvfLyQbX31iXLroTT3ZC/dfU3CpLT+Ae/Vd6jv8PaQFWdxVwfRkIpEb9I
bgMm07m+b3mrVMtrDPI8l/0INL1kQxotUMHn7r6rPPAWSdZsoDibAzO6FWy2F+IlUSZ3N851FArs
wrWYAlkAIy/8ofu7BXGrfcuRza7ULhsu2/L03xEY2++LtGERcoKdlXFn09bBao+RsUakeNoKRVp5
H1QttL6riEpnov8ITvAxlNTVLnQwhgI+Qpsb8Dw+k2m5/1/iF93EtAcE2vRneCJNePSqePhnubr2
ADahTDTxk0mJI2PZLGZAPOT5e8ManoGxeNgeu9vBTMOmADnQWdzpzLA4RnPRyvGu04P4D4D8SOVp
CvQBe4yC5rbyS00JiDT0GXTQHandFdINslyJYVvT/HMG4deRDWeS7teEstElq4R4GlveY427GX6Q
4jQdKWWZHcahK8u5g+XNfDVHz/yeEckTLUQlrkBEY1sa9Mm9th4i1MJGVlvwJiOxmw93zbLRuP+E
v7LkWjBWE+WfmkCzLbfS1ieNe+mV2WlpTF0wNun8P1+Jh2k31B95xKzJVwE2St2SMgFCn0x91iCR
TzyHpp0QdZ80MqY9OBjqes6Nzuqzp9M2yWaXkq/oE0WrGuh6xNw4VCwHqast5l+CoCNjewlenzke
Y0HEQMoFBT7IXWx6Gnv9XNfr8JywoLEGqgGo+OSVlIVGzPvGYiED9D2PAN643dkx8hkLQBPzX2yE
2po+M0HKs+6ZvJd4pOnoB0ybEf3OfNlO8p+fXPradOvzqVQTiRtHWxPlF5sJKIvuOks5O4/bRryr
YJ64BpiN+r2AFaEl+Sr4xNegTkpFV8wDKIuVXFbyW2U9WMzCYeb6WWjEtr+K8/4pbj1j2vNfHCf6
XhP4Xh/uF2eM5l9o2udIDrXoarEy14iPWoghTb5axrQgUCb0ThXr7mjfkVn13Q/dKFm+10Jyojx1
KnrWTWN1ak4Bmt+1Tt8y2MRsBpjqFRYXvZX0SUH/JYHbacY1pA7edu6tkHmqQVs3z10WO+DAVnSB
TBv+YJvRtnOjboFDoFmjANLYe6TII2VfcF+xV+7epW+OPATGfTzbVW49Ale1v4xwzq9xz5vw0hPq
XHOD0yhEYpg/KLZ9am3A70IQxCF3LJ0trsFyMGTXq6epOfjS7C5ktZl2oFtZcdO4uafMg+g+mVmY
nShMOeqiIdJQjwCA5RMruyI3RoKKpf3VzjZZT1Hgaef70cS5HnKsN74jpPNuFNXTl1FMG+ynwl6P
RNPXZvWWbpWeiy9qp9wMCcmceMSTrTQs/oFEzq2vfdbZw17ZDdNcxy1sjabnIhxyLm1w88oxfTkT
IcfRS8HuExRZm9Qa705lQvsiEqYVK7prtb+WdIeImpoepxmDl2GLiZiBKDAYSIyNftJUI6w37NDQ
IFJX7xu6VW7ozjsRODuMW75Uc4qcpK0Kv72r2ffCfc7vjz7B53wXbjHxENM4NnkWXnfIv8Kf/cWy
Wv9vWTUwZIsAR8UkVOcPmJgfl+aaj/x0Jbq0D4UFnn0ycO83Y5XlJhLqfBbEdJ9flcn9RyZBUqaU
xhvO4X4uS7lrgghy9fHFungY0GkTFvOmcpp8nAkeE4AUAEKFfj609C1z+yzVkS9wKrW7hOHB+M+y
RUytmvmz0jeEYMRWBYvoDLVOs3oStHBK//VWjcNf7sH9mcHBjQ/76NdwqYldACSgnu0vDTzOg5Gd
tDdBCkXr9UyPqxaFX02vhk+WQbncgpVImEb4XGZtzE5OOIhvJqLjzXx1MhBhw7kvbYp39Cp0B90H
WA5Ct6Yib/EqbGXFxnZhpilbiMUyvqIJbKXzuBOXjD6j1iSly+0JGXQQ6uShk8o9ezQUb8kQrydt
JYEqSQeri6lVkLIK9Hu2lv2/arcQBO5WH2YJjKhY0qi5Z7puP8jT0B5rFUBgkfXXe5uA+pxRKRW4
IZXLk7vGrpD6abbGAjU7X15lAfeSclzHIgKChjNtpwK9UkqjNAMYP7a7Ub91reajQT0uvFOZxPZE
m8WMwzfoMEiXIZiaxryZ+mm24GVpRjyS9aIYnpWiBVlUtGPiIRXPifmrKWYsAU8gTgAzEn3oTDw2
fim8cmrcgGhLy+sJmiVGhWdHGS/pValaih10WZCFpTBBtnYIA/gqwXAEzyKQFDx48KxntW+cPHbm
LNjLqDwRGK4w3WcGIYpnniskavg6QvrGmTcB62mgHrVCHIJZkVbSBQ6a7Yl5CwP/oVk9Wbb8Gems
nWqffJWwRzYYTwMOw1ifdzwdkMhPzkn1fibY7oor3H5ER5w4DXWtp7BPgyeOTGzJhzJ8nstG11hc
RxrfNPkVFjxmTuY6pvljZX23Wh9wtAZaApb6GAdi4lg9t98KVaVOrdQOZpLH9DuKK5mxs4A6cWwz
LJjFcPtSvyDZ0Gn0IREYb/ijk0nPr8qVXkecrO6xYhQjHaPLqMy074I1I8uzAu7BtfT8oLxqKKYi
Xcw3ZNjq2yirYCrV9OipE9JzTOPlhsXX4xDAHPgHhVEBFZ1P+xUo6hRyClZo3baFVpPz46v7j5Mw
+b0Q6aFD+ZBAjg0LYyi3NCdM33OGdrhZTRzVxVRsK0UzljSG/8jj0ZwXDpOMsTPaLpUfhsg/yLKa
v4C3JV64sEsf7g7N5cuqeiCwnU6bqs65pnd36nlkhWU+V7OPPZyFl1M2Z3M0APsXmEP1EKgNoH3Q
1y2S3TCuRBksuXmmrlbVjToEqHVXDxdDNHZrzoe3szgoTMRMECNksFJbXWg5hPipcpf1NYHe5jg0
0dQ0t1pOtYl0NEysj7S3apzdLuyRL3baxjJKyAudbYbqbN4nqNelsHye0vmokhrmNj+A/Qq3uoSK
poQbEYaXbuojqhBJFF1FSfaGt0uoqzCN2Jv6nTD0KRB/NDC4DVN0mKrYqEh2WOtmpEveKoDYeeMH
HNIqT41EpKXILZEirNPjPWQJ8YH+6K58ZcDUL6/JYu0pH5ZuJOzche+mhOysz0zh9AGi3SCxvhzP
DTaLNzAszUC1wOdaOY5g5d/AGWJNHA5P+rDCpUau1USRn1IlhTn7ZnZH0Em5VTHoUtJN8xGdbM3Z
GziWsr8nnaGda/zySBimNFSBg5NjOkAqdhdEiiwUY5L7hza6rZdSBlhNCBqBBT5T+uNJdKCsjeD1
UvHDnytuvwrjA/PG4DkRbFlSIQOB+H0kM9Rp4p2NwElyNclptNN1KTnhqkbV9+t2FieBAawB5LAv
0jMuHukNvpGkXQmRqzlh2LXUNArEWAQvgCdVvmvzbkxHpIR02/iFGdI4WnRa++2Sz/vC7nZbYAX1
f5JNYF0WzwpUCQE7Y34ffLmgPTXNidDjawYUIUpueJTnNnFAe73Eca+HlfOOiJuFacDTf/LpRCn+
GO8PbEZVeY2GZzH8v2Vk0LxKwAnw8iVk1JaC3TAhpi/hGGIY1ORAs389eRMnM6Fbcsrfu06Sh084
JyszV5ayxmOIqvk9fahGIPUij0ZREHtfiOLpi9c3k8Is1XG4nJhH1/AgRLBrd7E5nQR4VagZqdOX
rRxtJf/DRnRigF1sj3gE/mLcmzqV3/V+1aE8RjBX2VBQFExobLYx6GAeoJNcc/BpcED4SusC4D7B
xDfQixSAB95na1hz2C/E6vdFCBj2Vo6EKe1af6Hojj686cS88QaUu7EPSWdq+/2d4RIKrH6TTrVe
e3ul8/6Gdn37/xIuxmM9yYPs0KW+gHuYPtj97JtTXIC7fuKa8yFEPxNuju58TBNxFaPahy1fPzIL
QN9P4Q2CfCPJ/LU/Xb86XsAfxPPHvMm7IizAb4HElBY6dl8em116Gb+WgreNggCBGr3de8fCIjEq
2+K2YOn/XN882FEDjkZlfjaG1zxVj2lj2AIO58c896Xg5WmR/OsXDjg/pN3QamTPeF6kauzFDEOb
G1+YbJzAN5j0h2CESh0cSv7zge6ruzrEfB3Uz345tS2FOU3IuEbdzD7k+UR9fjVv7iiEs3+BdX9r
tCRd86Ug9GWXeNXtCaPA/dt5+9mgNicIQzT96cTXAITf0MnZHNaAyP4mC6UsslPmeziL2/dzmD4b
v7TNpe76n1vnB+E0TyV9iZG3BxHnpqAd4OXaE7ug7w9MpiUmp+5wo/L8W4rMptfpACObPEb3wXwh
oXsj8D98/E9/tVNBcADpMtj2g6aNa4StYcXzuSViV67BKJASYBYMnLYVjnkN92HCTRoyU+0HccfF
fTpVuMU6pM7wCaFTxHmrIsBV9anVDtgckI+gOPNu51x8rPOrSfJ0OTkX5yNcQKyV5Vj5qb1mjrHL
sB7m3UbqTMN8KlhdxKzWnSkAonzemCw+6LRDAgfShYyiiOzohqd89fJpkeC6Zf6DTBl7n+Hx7XWk
mDcdcdGMIsKcxA0KJmDCsY9HM72D9yUNK6RWitp2+TCryioE3oFbAt/bqh1/4OJQkgAWezXS3Klh
4dX4M1FslxL4QwESiyAvQ24S6WBy48Qf+Y1wV+wOjyy9vC575/wuCo+zf/VXQdcvD3Jw/wJnTtGn
1xoq1ayfKHxig6o5fYRksT/3xUfqFUzUCz4hbhWkHrx4O3EBaM4BJmZ4cyEjqTgK9Uvy7vbnVSQX
60h1aOnMvHfSP04ACOy1yI4VL58ffjX3NUFpP+7rSTPlmTJVD5wLtQP9IRon4Kb8hyYOZ2LwaFDW
wGF9iDW6p8Me2oTWkajjkIzvuDnzJ0LPWO6456ezm5268+qLihsO09Ng+pyV4SR01921g1FePslO
mfSKNu9uCgTcgglnM0lUeboukeGYHcv8dqOWwdf0g37YwRG42bQXfWpFS36DQbMziDpuxwcJyIQy
+mLjYoqyJ8Q81Ptr0Bjt3FSqvxVCky2cHQmpLhMWZWFMGZMqn1dMf1tPx6jGr9m9HNz05IEWHHL7
8KbyBPxbi3BEkolCdUww6yQM8t5/eWpEpmFKkC3rK2lfYmwJLDKSXNxEwRDNijyBgC6P7PrEE74A
p9Kx/LWBBCOCTFjLpNzqkGpu2zt+7QGqbuGcjeYKSKsFeiyR1K0sIE4T7exKk6Kwoi7zI6gH7jDe
Xn66OGaY1opowYKAmY7aJnIn+jpiBaiSJwhmySLLcyLftXvZAh/10jKId0SzL+VZ2E5JdCGjqxQz
t2OGGSN6TlZH3DSd7Tw2WTKZ3K9JOghPtvYS/URoe4LUOUSVp7oeJLNzBPDH+u9ZXyYwzChyeu1S
vbNvAXOFpr0g0M2AGjO3MDTUlVJJvDOlkNauyjTKeiPUmwUxk6A6ofyBEVT61SczwtmfWCqI6Egz
kidOrt2y9SEE94IUYi/7XJTZy8slxrUD4Dwln5EpROzb6BflqTWMWVhPPDE6bfMNNhUsLHEsD5Rx
w3Aq196LWs6lnEoLjL3N7H/KkeK2TZrxdoNEj8gpKfBg1m2CKOqHY5jDrLDoj7rRlToVcFf6p+/J
pQYPIe7KaPaUO+xzFopaQO2mJ67Aq4BmeFJw7j1FVQOPe/02HxDRkxrQfSMt8sZKxSxeqwNDU7vQ
mLfxtXVHFPp1OXgh5GnNUVn2l9iOsOht0ameF/96y+oyKpK5Q6yMUKnJBqsBMyJd9MeQpiUW49Ry
ikUJAYDZEko0WsooTF6f45Edud6N4YnT+uTFQRRJim0QoTjGef/cr2ATPNDbIKVoF1QKJe/1xvtN
qwhxTeOJqsMYKhIEKNX0EgkZGEaHattW5retMNdd1h7zQ2ocQCLXwvvbwNcC2oyAeyDAajVKnqej
tfNLqw4CoWx1+hhGjan4DS81S+XUW/ar2hvxEadx8pAYwqyaVaaxdf1SjweqOcruvaEpBH+cTbzB
ve9HhMP1CwnunZLG1BR54UOXmud+K7hU8sOHA9/6wPiWXQn/tB4jP/iNSS/d8S8v66GmXOwlUnVw
YOe/H4iZoqvt9PIKvLnnylyw0vuGEp2E+ogPb2cMX2rwwA5JPEgLaNg1+aLXmWp0CK4eEvqULomK
esTmfxXCHE5Is83k6FKcAu9MlPDMOzCFgB7JcFF4D6ia9JeCmehSIU8w0WOgRjABDTYaWTyED8bv
opetVxy9w+Rog3d205cG8ms/YEQsDuK7URtXnr3RFjsf76pU9Ke/rinuIRQFw432H3bC5ag4JLC4
5eJs4vAJJtLu74cEF2wOxinpJ1ALKearFn9uLx+BMAB8Zx3zkQPvUaJTx4iWN+lAk+WOQn0ap4Kp
dRk/DktJZpV0teFmPlz+Va0l4Rh9Rs8BW5l8HbfSnKxyoPYQcwm/avmPSkPe84Pq6Bx/QevxSRoM
qdSAxR6ap9c0CYT6VIFVdCVZt80On2U8U3nTPDCdrp4vJhq5C0/BJ9X9vQBkjrVUhsKWxknWF21b
uGzvqYojlz95eWe1u7woxFSwC/7hfMAkMYl2IvC1DAIz1og56R1x/PJHb63MOQrNSxMmP63kM6z4
pddX5j3Ar/81R1XSPPueIpIpkG81JDc/GhOB9ft7C3aTMN+4BnkDTHvtQmR7GMKvMM6uava+8GE2
8etQW6lh9RkHBi6hQfZxMQptMxpEXQNxWpQjyKgwGVVZMswnokxO7BW65EXa/wCsahSGSqYfqBUt
V0VGXqdMkuchjkkRMiLE+iLmo3bYey+Gsp/+UhtdA86lr+0oIK0NEs7vtq62np7xMtFGPaimYeam
9Dfpn58XkMdjOupWDDkU5A3M7119OAYcqe1HmkLiQghznbtUDcZLT+aOm22tP3+CuxYZjRya5LsS
bTf2/xu23FMBWUtVMvzFWPe2VEW/K4XPlaCW+xMGONXI9v2IPopNdI9I+LyOjw9slFIs5+MYZ4of
u3tihx3FRzohqO0DRMzpaWnaqN1D86bEYfeIpSoLHRYthUoJT2JhJ9KfTCqlBwv5WkiB6ugaXS5t
0CHhaqxJjySD0KhgIsrWq4sZjVSom74i63gkkX+E4c2yPL2CXLdKjLz69Mf4MiNX8juy0owZgA64
veuKVaFnrgv6bHOrhCPkbAVfjCS+sVP8vnjmLsrr5h405/LSZBcsqX00X9RpCf+xJkZpXbI/STZv
CZpuKmNKI14sckk2fRYajNAZYVgOB2tx3dhsBM1+14ZLl4xX9lS+/WmzI8ldvrxuykz4z+byvMAC
mM6/8OLpbyR7xTLrmW0Dv7UaR2QVbPWL7Qtd5Jp3IWiZ47XJ9HAjWj9dcUdFWr6MGdfW3pBrpGMD
Pllk6iBb5coOKcbqEqA6tz0mvhQJmbfDsoEkGLA3eh+OOPYVmRC1u+15sLQd5HkL5T9LnyijhrDc
kdPM5K5Eh1THzpLXdNT5Wg+ff4XVQNoyhgh0eHCD1ykZg3ucQN76jBkqT4OMdPvaaS8Cs4kqvq0l
GqN0GmkSvSvpx8Nc/Ffo20cqcm99yGq8AbO93SZ5bvxjv+gzCyQXx13YZqyZyMNvrErAkcHvjEnm
QDPVIMDJ1o7hV7b71Ega55c+0KvHegVV2CBniUBK1Ndtvu2SMwroDFwzvhX2oZK39xkfGJi8Z1+L
xMYKQKxjEuBYitq97IHb34TJAxUbfOad1RGouUKAGKMmKz1ckCXWBuU32cCSny0rFG7dcYcNBDaj
Wz8hcPGqMZomDA9rNprxdoYoZ0YDk1lUe8sQtPKVj8E5ArcGeGw4OUEK/0o+xiDmd4EaN1A+f9l1
qg3Dv0wW7AzK06D7o8FNHV0sZ3AP6G7ClRDmas999LzbdDMBzP8oz04TrBYYmqd6ew1WpjbjdGBh
KIYYkgYnqdcZhbvp7BQKUak+xqzcnUw0LHfW8Pb7X2AVmwpbMKx1rdpoFZpJp1/qdDcMC6e0UFfs
1995v43P+TsKCGScBGBNZ4thcXAxQ2HbiGLfX/Bz50jDx/QWgX8DEvgpiV3ocCUTcxzyud23B7ol
DDyQbRCliWX06QiRyjMLgMc8XphfsE95dz6qA4xDQNMaen317NkI38Y+vkD7rwhpxKCtJHZJ/OXJ
Q0Fw7kh+C59TyerW4M8vmwOozWSdfvZHjUifchmJHOmGIFgpZ8mQesFyG7SthXP4daOq3N6z78EC
1Z/zUNi0M6kgbDZBFxizQtGQVNmPkIrzqH9A8J/9Rc9bTIxgco+FLzQW2cjrSzqEqkZm3BoJJ7sG
uIqls6bm72c+NGyvIkzVaLE8b/jmaOubf0Wc/RYpodYpJUtFVg0Oq/gitw2vdvhkVahLcHQyinqV
M86N6qq/WEcqus/7Sifu5kuKYeWidfFvKldK0WfdQ/c4z3hsPS463TifONXcW6x3s0T7sT3pur2Q
wElkmiBApY13IZxKmQrD4VDxQ78UWOyDRpNKuFOqmS0DFO94U0UNDwz2FXieOHN4aXabhLn8dFw6
QS6yFUyuerWq382aXZg6lwzuEHtge9NqeJ3QQOxWERe0KHxMx/raM8x0o1zI0sO9XYt2PnGFWMBi
2/mv+3OTupUnp/qEn0GD6K7rotKBmgk68O7oFRVEHnEHhzcbtBYZxtm7pXCchnKkDU5zLiPTuS17
c+5XFQgFNmb4C4b1zkEKuUQefIy91EL/E/bQlg5Tbxz/iIxDjrqdNOX/YpRFh9UaK2JNPKvGxZ8V
Q09ij+K1wt0OKXkqgJaYTMGfr0V4J+BrmTq5O/Rt4o51CdtW/ZAQao5dgjzK6KR6rYJBva/QJLre
Nk+V2Y5F60DTf3RzURW03L3Z3fGOHKGtVyYucPB8NS/R7k2mg6F6LeH1OqwvrTXuvwVviJSq81jz
ppN5hhULdaNOi9eOv91raX3PdeiktrFiKS7lNlrMjbQso9SdqhKRrDZPDIImym0V/XbEL1/U9Uj0
ZaW+uPAA1FhhR2lTTBHoKi4cWTcAlEKK12Sa1qUTQ635y6wnQEdTep06OXdI0JSylH5pLngfD+uy
R0jRxFtSDbD9/pZMbl/QULal9rjUWqSRzIHdNyPzY4W4ebe3T/myEDT40W7Mnj7daYBwdwCu5Upj
fF9sXnNzFt778Sl+M3ZJ3SifWwYwkFfwWXXGUgEP+b59odhJsjraxscxahWlqwHHM0SpvUJgxHQA
80GZf8iG5M2vCo/nGe1SSnuPu6Y255qNtYh42hr4ObvXYfTl0oJOkRLB//aEjn9WWHXisNCUhoqc
sgiYRdjDZFhzfx6pelxl+Dii5sZXgu+eDiuHdhKzqQ4HWlrtsrRi4uKTtnQGXZZpxCzRTljTd5Ze
+e5Eqz5UtG8ojt1e6Wz2qPcmx7A2t/Jl41Uh2jxdozcnG0aDZV8pSckBN3uZ0mBVjMO3GAXkCA/j
BvSnmVlqRN6r1bImN5qNQNjSf6n3YrRFmfdRJ74XGd3xeGM5boHfkJI77wt+Y3KwiB7/ze9FYZt6
J2U21B399RUUwe8pOr7yruiwF7G3n+2WNw/0PXbC8ntlqhGn+uHyeMuIlJD/kdQWVpCQvPit5XjE
2g2QjW8UYjrGcdV5LgO+oA4VglIVbfsqDDCeqM59pBOCaGSkDqJ2iLJyJigsim2hNYirR/gDKD9A
1AQjU+Sdn8AloLS7KIvg5HEZ94eUEMFmL1c0Y0dlXwoawQaT/jRbn6YKZWcVT4D8antprRNWqfCp
XmID2YNdoetxZtR1QjSXs1f3DUHZqeP1SeZqlp4DnOIc3GO+zkBWHnZvBWcsbTQqqCxeUxkPkU5m
uAuTinInBoK1vvpjK6ufVMvqC91L1W+kbZbHxMONVMGSyYeuh5E1avelCxOuRYlMha3VCcaumgxU
NLukfJ1kL5PrD06YeFm+/+bcpaOd30o35s1S3QMyJwdOOqk9j8/aE4TIb9ZQ59JkzJRaTudPIXPC
aDlm68EHiV82tHKMjF8YMgpqWgoFmfFaL2GNKEKMLXRGj5hH9FULGOlqGAzR+qvkKzW9JtWtstQT
60nfxtAnMsnFOwUpIzEWtLPJnLAAew8Setuv8M/tnhn9BXIU9EC5VOZOM6sCE0ckX4hYstqwUGip
kS4pCICqoPpfSOLP42Cbtx+EygN4OE2MFvdPn/EIsWVYfoSD3MJSCTaN82aZJLlbvThpEAkZ8H9h
JwTjYTlsxrbmLtfut6gomcJTIZ6oSF+t1OTP/gwPFuk+XXP1EBE4wWvObeispg1b7AIBwjFuQUWs
5myLTsdGQ5OZwnAqMHjHCG0KiFmSe66eOm022fPb329dwRk11tCGaeCrG8Jlo0cpGwytQpi4NUzC
2G4eKts9fdxhY/PXXPcpESw7pp4VbhF459kyMBbR6//dx7Js2jBXLHOXLcyf7CST0uoC9JCciJGd
iMXgfJwblVAFADVidHwYTsnPYqeW8rrbMcLq0sS/mtTqgmyuUp7v/eGnhGtzXxYlow9vQs1sWpsL
kZ0LZb5qQGt6l8qIgKrT7qLhzliewvSL3dG/zlxPTsINI9tY4pPxiE5UWC3F/+tioUAiLcyDQuxW
Txv8//qHVyOPVqZuAkZ498/9GkR8mlhtVTUugjrmfWY/xxw7vnHjIty175i/4P23YoE9sZi8JdJv
8u+4tLtte+1YYhkJ6ljPSR3oMiBg1dSrNN4V8i8If0ERB9xOGcrow7QO+fg32THxrwz9z49cijSG
U2JlWdvOxl936taAvdhrUWOITcX3Lkkbss3NUsaRY7beBHooEkz5CbQ/ylL0/Y9MhIgZk8QU07Q+
7VyfEqjynbI32P11EZpEy60a3porZJoiZoPbJTj0kcnZBc11DuXZb6bUMziWvSJwMSishfvI2L9U
s/xQTDHSmk9UOE0fuS1IW08WJH4IqUWVW19Ttct+sca2ZB3hqmBSMs7WRgC8+zeP51O18b1ggvN9
4KVn4s4rZnqIgAWQwOkQ+tQIWXX6ADduK1QfYpCe5yN+E2Rk2z7sKto+MIEkHXRiaXK+5MJRGzz/
/ZnUuz1I9j/efe/GAizRUYr0H7f1c/FSZQH56Vsu6v6/N9v8RgkdmmF/4uyAqJxaPeSnivMOcRGB
V3VTPW2RoNsHPoHu25EcM04L58HB/TdFNdBmqaVlna91eGAAFZhEI6VPWe/VqjxmQDd1GPy/SKJc
OX/rqa/QDii+Aq/LIAvijLz6YzKnP+UnhI0QcnkCyiUCpHY7sEgz66L3lKYAxZXUU9ZqR1kJHXzu
j3EcYP5VyBd9KDUj068jDjYPEx7369cAYeglJw65vmdjJXK25zS64ToYbBDlPO56fUhi3O45ZgZl
01oBv2s/DyQlrt2CdWggQsOIF4GGP1FTnMIp21/WhhXlPg8lsWyIqWc/p4CaeMZlrafmRa1Msxeg
zsddkPvnYw1zosDtI/4GaWE2wezJfn56R8JJsxUh9GXFKhk32f+WJewgGhEpGR+8PWQtWjxm9/Zx
lkFlI8ManzsWn47Kxpe3NmsBvY4du5dIMznM7Ga8y4DUp8WsXulUbJ38vn1AFgL5QGDKzK2B3B1K
pqZHczw2fCdZY1ums6C5S2gy7ZQUv6lBlvQT9Sn4shnup6qu8I7MzMtDYU1DhaiaFshnWQV+5Pyg
uLnzfIYTNeXi0bAYWgEuDB2tnYiBK9ei/an2i/zw680SmhdoRj3cxJaTw98nl29qzcedukSU/3j8
/FSRlLe6889lygT8zJpOEr0FVUs9Dmzj2KiVQY3R5W+95xdA/Ew1Wldf/EOIJr9oX5GLmbNiwWhx
zgw0I1fjEMxCHhC00xFS9eGjd6Q4t+s5cf3dVkmZAvVIwSDimqZRXCO2MR2XqW+xI6BLX6BgPgqN
CrzXVBj1L6k2+qb6GR5vTYwu5M+4rxhBPOalMYAdqOnT5U5m4O4lQZNCuGQ6s7c9Pb+hPOwzzRsI
PIcOA/f8XrvXBGZo9GLSiszsu1jnjDMXySDFsaFJ2w2O0PdG655n7GlZl0ffpvZC7WTZGRIykR2u
l/VbG8NpjPNojTzJT06uOnKzUnHBU2QV+1wU8XoyM343l5jW3F+MgYXvKUuty2SOwHx4VJP2lphW
EXAt5acLDpTBJK6/RXxu4EY5h/yr2oAdLCtr5DVU/yEXyKg5OnNEN194HraH1IDkiPvJ25cFeGUf
fo8nCyrOwn8pXdKnF+U/51N0CbsKANBzZ1GVEUqB2NAV5l9GVF26Cdk/cdxwTdpAVEUCnC9eH6J0
wqRh+45GV4zrzVt30/jZT9f5IAe7gCy6Vib2JVZsJybK0GOLyFxQi4YW1yR3CPO046wMfqRwW8lt
LGWPecAy0MXSXo7RNbuHCV80oRucVldm6H5MSiOnO1/DCOgO9XU7VFHxGAxYo3cP2Gi4nPhc7lUp
pCcWcBcpA3hX89FjbcEbUllSfgHlLK+yT+Ts6FhfnUBL6b+Qt9N1XI+RiZ9GFSSSkAWTvNR4NSTo
5sC0fSnNB92thJ51DoGrx43MUGrXg8MIKMAXIZEPMcBRh533BhZVmVx2xdxv7p1ys2LzlyCb6KJJ
9PWPBPl05LyVRGsv2x7gn3WLXXJaiczzxXE+ddUjw/dUZ1e4vKs0YN20XEU3zTF1kDbQo9z7h1hI
p5W82X8F8xKNX1MqwIyYwbCl2OzxWyHsY8zanPf2Gh/xh+dogg4026DJgChbLiTYQYHl0ycF7DAU
UIKt7iP7yfL6OjT/z65kHxMhZGbto4WQEuwiBfGoyQL7k5QNIQEoXcbc0bW9SyPnDAzu9ijKNQuA
FATcpYw3fQWV9kdl4gcNiWbpmWt28/gvQ16G3AJWkAo9X6DEXNEg+uUHrN0Te5zlaVMsDnRS3JW3
ZlGXUNL2EimeF1FZWvoSQmOGq/1bCGC7+QJL3iwklEOaUJ3TJQUD7S9ka+vVbQSlENmV12ciWqeS
IEZLDgLIvCuTtGeYEFxxc0ZUesUvIi3QvuAggNjZbMzXmPOFdNPDJKdIoORPs60w52U51B29KvmH
DOFM5SJbIZCqSA/ihj8uW+VhysF/2r8f9oE5Dy/Nk/IBsCiOpt5yI1oNLH9eP7vC+dQ4JBvjMp5U
P/4x2Wr2np1eja+T0cYaTH5Z5Viup2WSmrr9VgW86m+ZCb2pMVW++ZYxIgWsEn15hyHdBqWjCnQB
NyNZPaSnYu1777rnd7ivF+RzLkA5fI2ePQzIrCaESIyXbPkwJGSR2amZlpn6FfZR61CVoli/idzN
vdN/w9d5uml9weksK8ABGhu1vFHKb9hQUyRedg7uQoLV4bsuTrrRHIDC3QqagETy+Rk4ucemomrg
oonpTnnyY2sW7/nu8TvM1CfCTGcADsClZI1wcPRARuj7mldwCoJ73gDMBsqd3p7gBBxFUboIZ3nB
zV5FUfj/tzQSDyVcECR0eEmz72olIuErotsKUDdGdQ5T6nnnWaXXdk80IMAeTH2eTz8o5GnbsqWb
QsSNE/2r9u+B798sWDIAhRHW7UJl4qNOmAC1255SJ66C472jXnoTxkgelyxca1IHMVx6xoT/gjey
oIZ8v6BBPoIUZNkrTM//gsdOWG6gP0urjYNmjUp9Sa0zJLskjUqa93amv5qGD/xetkNpIayRKWyw
z6iTFn07Tq4HXtbO0lDGOOIe4wpA2jBfZWNXdFem7j0jYZ4x6nFhiGRSwua4AqYHBiGwu/Lu4ZQA
n/IWASUscVA+KFeodlhoDivjqrBlmBnBKrdywIreZKmk8f9J74d3EkpkBUlced25U7MaO+8Canno
vyge+zHkp2Mgjs8EyumlcH+qbQAk6s+1zB8RBurjRSnPK8abtZQda5RSZP9OjnQUCsezTnRsh+Or
zBDXlv8GpLeBWe3lQUWkaNQm7qJTxhrvf8fTQYovK8LhkpPf6zDxJRkXP4tRmVPhY56BcktPBxnb
mgJEDovPMq+xzUfKsI1V36c5qqTVKthkaQ71sxtarl4CBYZhCCSxYBeuVZ628MJSFkFE8H8np4Ii
TP65CvVKzV5xcpreYvQlIsOOrhDPZolQZgJtyjkzoT+j3TwHnJy13RdJKhfRFoyn8oBoVeiLv9D/
3tQu/D6bcA78+bGnYtIQQ1CIfQNJN5eKCzvRglFEdJof1q+1u3fAfOCZvrLo8la4e7XXd40726K7
n5IfrCERgvJJYjdZc9IchZVozBYKp/GKYH0qvfA+W785PIPOhuUz/f6b/hIqPdRuoCX7drmjS+Zg
3NMT4xhVv/pmr94z9DiIpDRD/Pj2l0mYhv37rnj+7RMzeaWM+V5vC4DM6EgJ5ZqlE3qDNJO/1JM7
c1pslCdITEd+uTGbYArZfpfRs8543qPSmxdtAYCMGw9sr/8+4dAVaA4d9PCTo4DHIxvQHm1Zw9+o
FYvsFZLBL3En7CfdBQuHXmJnyDwLWVdqm+I1srgpX0Zr3s2HwwY6zpoJmX/b6QwmLYPNvMKmlqsY
kUZHj+6HFsrcrms+MDDw3G4HH3hHyXsTtBnwm5IL8hVdz914VtVESB1LpF1y7Rpje6RlIvwHrR6m
qsD/bU5X17j18AltfZW4Fy8tVoJJa7tyotiDG6Gl5lVQqa1/KpxGBI7sTf5fffSukKJ/GJxAYGCS
ymUPlvl56zxK3DdqZUy+UlQ4JUCXtmEq9RtHjWDLElv/LvkzkxspxjiWWDvfNTowx3fZQcZaNJsM
JeZzVD12+a69o7V1WLcPjdgltXoUIVp11pVRVJny2gPkP1SegW8MpobDSXiLKwoFSyZ25mPjhexk
deEO7lXilNhxfwrie6ttpWRah7ZS/W7AgzvccW69AkPfzvx11XpzhGRLwjxd70QePKDXSmOwmjw2
asAY6h9JP1yOHesMP5oJOgdNrmVwQwZqs07PMogsSBBVgFRrFN7C8iJf7OqADjRzUMsgmkOgZ+xP
d3fNz0uNBMUrNM2mQSwtvjPwFiynfDa17nTg8AdNFCectoEIRF0L85rnoaoaPGoAcT/XI73OH57g
xP9Dl7n7yxKfXZ/v8DjDDH7uY1OUSiVDFDsam6oZticQLSOUOOj+vSr296hqkj07ZG4PnH/eukH/
/woEhEydMpTsAR1rOQT6d08xzJ1O4Vfz7fr7zmoRwTwNaC3fmebJ4Wz7TjZnHvcQdoRIVGnQiXpj
I1jay4+F+bdFsE9Z2jzJqjZZrKUziBzl7R3y3mIb31Rhh7vyW4dS1mp0ZBXeCdr4olSdHFR0YRP0
1pq9TN2Xa7i8deZoL/Pk0XtqCAm/Y5N0eXoAq5Ej3anBNEir/dwqyrMO0OtYK77bfANFeHLcW89U
c/aTVE5zVjE3BtgLLYpk5h0zIfcjM8kBm4+yYYRgsH8HuS22oL/epoH1OFn9n62sYZxtGFNjeYdN
6QdJOd5PPtfRjICXQFBkJnfg8uWTyF3gRqRQkDKsb247qg+UCCmAAyg4vxFt/xoRfKMzReeSgjbt
DYff3inulFl4aW06JQfmxuB2Mj4v2S80XqkWAWLtsOdxBIaI2ugCs9VDfTcyEp11k6wMreEgTaQe
4cEbAs/sbQJefNQ+w8942TOIyYdBiEAAuzCeOS2t/Evf+epYkJstX41pYHeHwt+ZKmogOfAJBby8
bKTaGCgLMRe5VgAwcdMPyQBs76j2hEzOl5VMPd8Dc3+lKw6I0oIrG5HQ46X3HlQQfsZ8NImStrvq
Rtq17aZ5e0XULBxQjGXEjqPITnldkEoqNRmtOktZeNC4IoDhQGz7LxXbnLA1rDvvGlrltK3+dNcC
jxw9Ruz2dUREBxFnjNc9f0NLPhtLG2CYvxtLHt3oH0zSUYDMiaMNVLE4jHpSRUcQDV6XWGYo6/qw
r6EwzIbsHcILPTeCKIB0YrSsIrIH6tGoW9wX5A/vxBaypWWwAM2WXDgAUK7X1XkZ30uGwM4aGcw6
e+KkYhvzIQb4Eh1eisBvDwXK37zP4TWPuR9lEnBAEdqkbLz2P0u0IWzuhg8y5sAMG7ltuBsuD4tg
C3KRzAPw7VGXuEmgJlygU68fddq6ReU1tPE/45cL8lvkjlgazjZE5BLyGoq47Cg9tcyBAqjOf9zT
xepoVxKxWi5PPwmK5UNnp4j8JJi0o1fuYqWrgRX6w+2UWxT0hHqhBNwwqeugK6Cumdn64bWwA3uW
pnYVtQ8N6MgxEl5/u59KKfEe3O7I1Sb++1Q4XMf1BT41LJxsW5Ym5rPN+BodpgTj8IXFGVF6pR86
awvXFmuiVhZqjclvUv4/2sX0msvSBmjAn87IEgKag083Wb3DE7PcO0IsOaYWnfpKqFAY6uhTr94h
NLGF3MI7KVEgANn1QCbEcXcPA305C4LHlmwTAsyrsP4EeJCqWAZ6FWDmYO+YdKtl9q3PGDu8nRyU
+pZKO0iDJR7WsSWsNN9kMlq9L1xZq8zSO8jNN74P8opsE/oY6AzGDQNeDj5SuHmel1Xqo3VwENPx
OfGXenwYV/wlb40e5uZrfTTiOoVIkXzlzDz6Kqtp4BTPux+JenSNGtC9FxSTRjZ5bJOAOGo9YQdh
5qHq3+5jA2SKS1ysZQU7dZQdz4nDW8sxQmlVaQyr7j3aIf2lAqc8QimGxaev+0PUtRrqyOC1Ux0C
gv71plvkdwj7LSjFANmXt8SqSYDSWadVWAW3PFajqP2BDCidLRwn8QumbEXE0A3xDUwWhLpiOqZe
ZIN2QYBl3/PIu1lfs/dFH9IdOEngDligmwy0wdWTdnVzahTjIWlFsWgSKHWuSh97LPCFFjLD+g2x
KzrBQZCAnYoB6Vt1x4U3oHC0jUBx7JW45i8KOLv30W7dVGOMlVQaAJDyYDIWSr2VYTAmgMsLe1cQ
1BGUFo15FrI9AUOB5elopwmU0GyFj6ZNAeTjzReB42gCS6eT4Dqvzsdqxqd4EGx0+3NK8FgkI7dU
rj7RKhBrhedapETsO7llCZ0xmY2Ai5uxH/RTyr8lq6A4sxWM1KFgx7bexb2hmqPWnUvTSSS55mtH
rXsTEo6Q4f88MdMUn5a/kkD+iHkrF/YRvzRxCfSUQ2yy0alaqPz6/9IbQyzpmUWqY/kqehpjp+Kn
IcZ8S6NIMPGIEnYnw9F/KpNSPEuGPfJ6EsseKrSFzXYAuTXsH6HUp24YeHP6KCPO1oipxHtdYKJ6
uq3Z59CI416xN4SaUvHbhhFHbg3DAK3OWzcvS/0+/XS+DSFfoq/4aZDkBRMJYmnSlnp1xFMlAY9T
e/mnnRq17mRQJOSXtP7atybLJSlVcX8F0TfYfELBa7MS+Jty/HECNc0Zcsgf14HRAwoOd0zL5QLM
glA0dkFP5LhtTqilulUGUEyA8uIqbngGK4d/bM1X7Dye2ArcdUX7ydsa3JN0f0xKPpo/J8jlMz1k
KMZpeBREwKNNcrl/77EBl7Xh7nBE3/GU6vXG3nz2hT71D3k/Qa22SuhLnWGgoV8Xy90Q85Ekvgm4
hNon2Kudx/xITSzkuR7A2WyEHktIJiRgIYYwX8qEQ45bw4cB5TYWe0BKN62SKhEH+IdeO4zsmFy2
id1pktZQGKmB3Fb0QVQDtbmlmnjOM/dlWZPBy5rV4LejmvWqFfSsyLYsL9Eqk/XB+MyWgTPwb78X
VER5l9Zg11Pb1QlhX3V6YOJce/5a/EH73P279AEK74dVFo3y5UjIyCDe1AqXgKhA/oXjbmnVzleX
sbzABlxiC+hGCNHgPZNUOuhnnHW63XJsoegHUxPRUbio+PVab4xXCrqFmPkvJX5hiaBfu1e26m4z
3s7YQk3ZiaWgRprXgEvCh3BvXe2gAdPIJMnSXqvbzLQC9bsIJGx+QYgnvmQPubAqsw881HPj0t5q
tzkFYNcsstRP9W1WykkUNLDtVz1x16XbEBvGXV5fvn5LxLKkYT3hP+qKBBsx5ezMA2tteicXaj90
i8fMgiXND+aY/oH2v7PC7AkfeXQr2OrXm/pB/amY/G+HGgpIqaKm/o9On5alGsZ5D1JaAQ0oIK8E
Mg/L4kxD6voqCY2+uOB3BiRh+rrKl178HA2sVfIW2R8jY6TLfwLjTd6Tmzxxd8R9UP8ts/9cmYRA
gG+9b/vLryZlj2F5DsNY/C9W7EYp6iukISuhB/5fokAl6mL5PSO4ufkS39hLMhv5BR+9FokHaXM8
WBXXte/en6yX7hg2KeSCCRjYalqE+dfvjEFfiKObMJsgYE83vLeLq+QWbTbF/Sj2r1+SHyq+RtGk
5CPLtopph3foFTgMCqxrNPn4TKlIzwqKeZJ2+knwCFY6AnqRTUF3SHklAZg3x/D8FiPJU6bgp5HM
wt5EQf8eS0pY7eG4LAwMP2dLIRBcrBg+WWEyeAcRqUh6XTLIKg3u21Gl/o7OdDwO85r9TFiFSAOq
3d3be1a2mRQHfTvcdBWw5d+5Vb1ZstvcwQrc4CavydM/QcymqBB923MWPGKy4TkKw0zKxzQvU9+9
GrhvEOY0QmzkEOYRvTgjov0GCZA1yOuwC5eH+ZPa6R/9ymsGiIL9TaoA6NXEw/7aAwBit3hYyNvj
eKO11dMxDWW0bjMhJa736+1NwPR6G0XvFpjsj3nrc958vHkt0ausnbC6y2aqYppM9VIme2hmpMY/
PUGmGWv1jx1reTS0/DuVcarDRE+UJgPmSmpNVAXTYLiow9FFsNgNwu5CgSemIlZrCAlXJmhrKhBe
OkZf/osJePYwxPOUZjFa6ApC1FbFpAzAt9UbNtsUmGigC8jlZj35yzTiHF6hE8rs8wF2VIIptHmA
qv2oOjBcjgHcYQezSC+6dbPryYLj4U1tk1XwETF+BMLUIN0jmX1kQ4LVGuR8h6ISeDVbw+ECAkcY
k4ATeRyfYbsivnUcd6Jk69gphwvjuxaDbp2uMTe/0wIY+l20blRDVmfb4P635NAUQlhcEc89flAB
GexXDMKDrQ79Ugw4O5+F0NMN+WmvcM9fKAoZIqTooSx6Piy3lZCcD34T3bP7saQeu8nuR7u687qw
mhQbLod8HohXPNqWi7lnG26EAGLBWBi1PJXiA+a6wrL47JrO4gTNN+pznhPWfS2957poDkSAKbQH
6HK/sFuVdVDokIGFGOHi/NXxZ3rSDH3zVHQ6McsgS+orgRZ5HuFgmu3DkvPCaELEGkXTZz99IFaj
ZHUPPAbgtdd8Bwc22WRExCXe0pX2ElLjTTsg2afStaTFL/9Tp7jE7bhmeOvsL0q9NT2doxcW5bkT
trI/5iZygB5NOxCiYZlWkdE2MymxzB4i9hKyl8YYWW6UtCzfpZwDFvxA6O4b57FDtivA09926noR
Zco9OCfWcIKBMZvuMVFN5T6j55Z65/RMhPOWDepknDGEU76Yn9katAx0LFDCuk+eV/ZPYv1Jixl/
og+Jzh9L+GPWjbPvDSUC5+CXaWyyokvHaNdHdwudn6+7Ilhk/FL8eSte3r+tIHTkSzXM2wkpzETj
8snztoxqo76FgZOxbUVu3dVCmA/hQrElGIiYfMDXepdHXu5nupgZBWR4Ojz4EdwDnubiHG5i1hCR
Y8Uaz5k3PP3XlwnNkK8goxfPFcc9ap+Wv6hSqbQMVnlIhGya07JkX8ihR1FKMLQgT3l6NR0Fbjnc
H9LWEBrNz6OyyZUBR0eG7UDs7RhiK11bDHrgd1Y2nQtqfOBrhYHSqFOsTXLDw0mgJGOsN4erGWsB
A4M1GKMrS76PQIghTaDWd5EWeJ7xWEhzQ/rD5JRPgsxTOAQusJKFXmyP4fN2YyGbZIvdtbiVKbV0
+9ipDU1aGf9QTrzX7h66U2M7MLMs9P3tFEJ4mOqpDLzeUlb6G/kKMBBpYuWme+HOfiDh6Y1mhBKH
JkrkE8D/J2fMDCxzj72EWdzEsD6TTWFurITbBCsYm0s7h36QLl7s0+ap7/sA8HA2FZmG7mdN6N+y
XhnJR09ApJ+zdDI9qIka9PBmKDQpSA62lht0cKqivKk1Nh+l6su3y98AebXXQum3ZNSTGq6qtIzD
ohFx5xBQUqS5MgtV4aKRuRZ40QVlzL5/J3Eg3mkvi7yExaCw2DmYd/C0Zzml+cl0jeYREcRQBK7s
fplVZWAlB56bZn9h3GWyUwSpMIM1zLm+omkLRvUJOxflfO49nDdkJCD+aZJCAxXVlzT2+vxs0u7i
gfqiMsWiXEvA5urblEvKemwYOU3tleou8KhGZURWlKoe33+BIk1slQT7Z/IsK59PX/0Cgxbuoj/z
Wc0Pt9f94NaCueVbjyc/smM+IYuk4xq78pHshp6rQ96Vn3DRqpGbiK5vYN+ZntInMKgpsTynzq0C
HIgmi4jYYACxdWK7fin1l6rKMVae4EIC6qL1cmMys0aPM2c9UvsGtQHsup+cXOS+CPcJG4DQ/Kgw
oDgL0mNUdiag+S3RZbiuXanl85ym/RQAEBta5me3J2cXxGdW3V2ZWpeGqEmKWldk/DudGgGFJmB0
L4PwwIi0Tc2ujIT+/DaDodd/wEGyFYcMb7Mldrm3l/LyA8ZVwPSfNTAdIjFrxGr4bYLez99t5RKz
ve8rz1TS+9aTyGSha3qPuv0nAsx10KF9YMpl9zMo3z/UMmT/0CC16J0f8hKa573sl3fha6oURZUN
HyoIcdAEQ4z8QZ1W6VN0hYvSxobkY8fIx6N0vmrYpwfUb94x11hK+k6gj2WlFvO7433IdcMqT664
kGOB9Ckt9MAV1BYi+mBM6/iUddDOaxAuZXiQsBnW1BeSzpXvbskZTxtIO93yoDFGCHutjO8W5/zC
Yek4Kj3mfNjArZiUW5NhtmeDGGv1/U5FVQik/0lyJ0Edl1gcP81y6QE4DbvdFWBPQhFjG8stEyF6
pwxmwMwr7hsXYDHaA15EoAOEyMGvrs+whMCT6p6hWU0XiBD/iNRLX74biusG/SswYMVRju5eE4vn
oXOzueUXYzeOYj7H69q3jsVp984dquR1vw3haawbLWNccJE2k5rGvaMyNqwQQY37hrj7abw6FUJ/
BGK9NTmwSSvFcyTOiOeIetrJjaRD5JwhRMq2GAsop8bMs707KstTFfnfV3cWQqNd7R3km322hfu5
7M84gxpDWmzz7aBXMuBMnOQuk6YYMJgENxDQT0ZQtdEYhGnBu8NO0i1o1VX8J7YItZotw3GmhHLy
7ADC+sGtn9yyEe4kkJK1Dj2fhalISnFfMdR/m0iu+TNx5qrS8MzLk+c77SOAvViPEM0ajhaQk2Q+
L8u59mnsxKD03cjQalPkTvd4bduHfKDYC+u28yU1qWzeS3Fo8R+/CjE9SQjh3ov/qzod79aFAsFE
5WNzn71yquqY0sH3u/akP0pEmf1CECvXnqesaNsgENVisj1Tf8eur7y9ETte/gmAVNFb5gp0cuuT
dZWO6BSEQVHpv8+GbjLrRKBy7OCVgSKGvd7bHOvpvKDXgrNindVzplpQDuH8BViiy7yRTC/kiqMM
WUFNQ/ZQ/qtfAKiK+EIQZRVfF3Dly+hIfAlcVbjW6WYzm4sxnCU4HHP+TPJGzSIR8/b3TkMV0B2p
iYO+HOdXNzT3nSrf1yAVrz2QaqpA/t2EOy6cqgUiyH/ODh8lXneTcXLy4uxV2wgIXBQQAFUV7Cn6
CezW2tMc0++pABc8Axh6J/j+95kJA5nWaNtVgFPedXcSvGvcqRPfeVSZBy+qcX8guo7VtujIbrJT
uhZztuPOL7dLk6OhSFIwSKi5OUihX3iS0fB1xL13EbuqCjfxO6938IgRA8/TWfEUU0rjgXZloGtW
UlZ+v2ZqRSd2S5NVdO2wRxvJZiOHelLKd7+nTV5DTodrgtnOd3/4W0S/PAOVGdd1TRADXnaGEpjl
4qPnR7RntDAi7SyIUINxqkKkrdqUGO/U4yqu6vCG7nFowIor7lHGv/EsE2pt8CfupVtWqsFkXSwa
oRleNNfkTB33ujvWSJ74aJkn/5ssOIcYM57Tdz+A2BBSufd8HdMRfCfyXNxyruXlZ+rVsZL/hJGs
ElW4NJf99b3ZA98EIcLCthf5u8hTrhq09Vb5OhKc64f9fMuy8xzyXNbeQodGIMGCvJfgybFDU9Uv
hJRTeQ3paiTqOoINOmtJYA4254FULHRmi6pTxShDcTv6n1TXBwGP1UnV3X2YWd4hnvSJCaOyclMw
8NhQNyZDFoK40xM1ChtNLNTdVv+TPd39m4fvn94HyZywzDo7PZeVTUvv9Y6c18ITiBYBX5f1Pm+8
OGBGmhw4faosaA6VtSeEKgoOwgGgIFgDplKf041kd8YzMNGvs8xxhhliYnJPxAy+B4jzK7pKbqJh
Eqmlv0/6GZwDwll78RlGMRHbI5MFqDl+naDYoxgU0oXqYhRTlk/msCu/ECk7dIjTIFTDofenxYUt
O8nJddMDN528THfPzdSc8jJKUofUxPTWv1QSV4F8/ub0uwPyPR4OYRK0jFDr/FKinAg8gwvXk4tO
nCWXOXKupOVMFWxBtrtNpYeNyrIC2X9nuSx6bqZl82sYaDVqcFisK4kLYcetslRLcf+dfFPMU9w1
wpHyb2PS+C0tDGUCgzfM8MDtIgWVlZHzKbJgZU9Z80jM9AnoeyCUF/hdFKMFOe8JrGywr2xCCnlL
Bal+Pww6s/DTA4oHCAyI2ZrDObcxyTo1uXqcZufqFdCoO9RWVDAJBAAbibW0pBT9B7YUy+/mCnze
vd0g+6Tg9EMvEyd/DsSY4d3FWE0hZGk5Mzjeh6YnDlcQ3mYBf4CQAQXqRpfy0niXT1df2EKuLU18
u4nvL1xJigMwKnU0yCEZ/y4Qj4co9XMACNRG5BoAUmjINNrm/9sAHRQT2CrSVxfW/UaSS/8zih3W
B8wbm4ENGkYa2cT9ue3pjC/H0dLwJMRsHwe3fzbWtXeOSO75LFVSE43zNBHi1D8OMYJvzZdXZp1T
qsLJ/hmRA0rcQ9xnkJEkWXb51lryllx+JeaOj0aoJQFnJ/A+qROxTeh/jAgZxUI2V8mLqHNusiHi
lBvib7bGet/xgL1hre4/FJG5mk4A06ikr9Qz32U3w83HymqrSBhnKrnts+gtdihxy4HZvS27KGO+
slt1d2NhYK0Ph3BYHE+X0xlzTTbHTm3Qg/qhI6gZRD8acovbdUPhg1Glz0lGlXAcPHvRxxAlipHb
f2kn5HZb7vlj5MAj6nFRhmmiXGBjrYWrOT884RIowi67CUpa7CECXVPD4u7l2RUXILuc+M89uFtQ
PrM6sY8HzBu31iKWs8NnVNNR3Eg+TDGGoXXSHmvJLwzoaBiSI0uzTwOEQ/j+nitvbmi3KWbT4w/0
1Rm3DtGq4q79cCZfgeoGkyCl8QpY4Dq/RxiF8rAVIR8WupgdcdTYaXMiLvuSxZEp1Fs8COr+222s
TlKT7IdSxhDJ3RZq/dohZuWNYI5ALzJsejKCF4QZ5gT5EFAfMD3qhtDOGHUZ+K9InB0Z4WHSvlaV
+p6d0QEH4krTE8Tf8FPGo8hyE9VikeqvBLyAWJsXBU2Xm61BiIYX/r9BVp6OiqEvg5nxJnlCv1Mv
jZ30dNiXdDqef3bmc/wKoCpCMoPKPGp4SEqFj+/Yl9L8EB88yRlmtlst+gACLKDQa+mR7G6kN0Do
KFc5aGEEGGwUC6qUlRV765tU1H5WOrESlBBHBt+qB93H5IvlNKVZJgDvaodQ9+M3xsqHPPMV+hG0
BJYRnZ08Q+ZBwJ2ykwYQVvqwptzAxyIUK1nmlXUW1YBCWMsthnnrG06j48nUTTjksxnlgF11Tdcw
smD/OLfLyOiACilq4IOkQRWHqEdJ7yTGf7AvVZGN0DTTJbdZQUu4UmODmI/GDuEmv7ipQD/iRm7i
oMnL+qlOkC2MJ/PbaqRvUM/my6g2NaNkJKpN6jEbK+F8kTkHq79jFzG/brRH9joe2Fe5uUe3YfmA
ZbO4V5Nn9oBLLQVmGINI3b1tu2GrfSx2q2J5vEbyHWrxaNMzB/uXIVIhZ/8aXDaTqX+mRBeJ4wej
zuGSnl8aFaA/7OSCqRR0DiZ9iRBF5lGU4bZ8WKUdcKeU2Lnq86rTkZBheVHExGG16PCfPZWdUMEA
19XvQVJPbRUtVpJY6U8HF0j5jSa71CsVni7kuk18DDWhnRKGWRRdjrxXI5rvxE7UUL0XSlaiyvl8
CFC8TSscJBfjNkVlHS2GX6iF03qS8kMwfiC+UTEFBdVRgieamO2yowPk5hw1gY/mn6YhRRz8ufO4
D3lXcY1CP3l0ytXZr3gjg47ooucyESmmqOqag+izZNhi1ElzdKJik/tZx1jmFY+SiG7OMmSvFfgS
4vevao6fFYqwRLyse9TfaX0xAFk2wjlhrtcoHIyhE3CCdu3dGkENyLZ8SE5DDrIv1zwwBD4X52yn
KubyUJ0RaX6Xy2V0+Ag7zcTjJ377Vp5F2/gWpP3djUVW6cZ0PlFao/LEKdoHNiowfqMbYP/z/UoW
d8BXWc7ltOPWYCa3H5FVgiq3chy+jPANIUoJ2Wf0L8mpfgqdzX/9JywUpDb/g3dJsHDHtLFcrd6b
gduO3tEk5yR/sLG0JH6D71t9kLZiQ1vjJSXziVEBw09YFeut802CyAcNxfdetRGJlWauGpyjfU4q
g8XZub+Qbmd8115sOCmDlSs/56pKXr67nGMB7oQ/2A+/axJOLNU/rt6/yyirrFut28jtoGXZRgvw
FB7ejKLkuMPst3CT8QhMQrOLeBbLOm9K1rrC6Ju9YpfmBZS08ISItJ/WL+ccpGwOBmM0wqN41RhH
lH6QAVJKeS0Cw/XEB8WALSHSWlxPjXJXczcQf3h4+c6WqJEKq2TENhuw6G6Ak9ySDNMqacSFj7hf
jNm67Y0qRDdMHjJPxeHuSmfAYdG5MaU/ccn8DyjjMwRHm52OFNNR1f8szepWc6VZwRvWl2TFP4KH
jNZykGFn8wAvPDgXvc74d5exAdGNZWTwcpyzSCT5shvnQ23iX6V/oXVh/fm2mniCe1S1pMFP/j1R
i9S93plDx71MvCwZ5qQ9jj3tA985e7XnbVEShAus8Kho6GKqNsvjEqZcJgBq7SnBSIIcwO5xeknc
BfaTOvgpG5UC5fhXFCPeC4R7BN+KypsaRkpUNnhakIKUyGn9L4SrylucywD2gH8QjyN1fsuOFR1a
anNpCMcOt23ObaUGTXaG65uKTM97slVjdiH1f/d4RCUPYQ0k6UAL2xd8RzvQVTe506HoEz8W0Y8U
GcFmwmxYbhk4e4WUXgspTdJZFTtZxj2D+RF9aXxxj4UZaB2y6Rxb0Okl5M6XNlZ/V7YwEUK1fqBM
85XtCFQKtsB+58Z0um5Mxf8N7aiVWjHZqLhO2ZufPUBz/JCetKh8Uw8fORaHX34KZanpdneqwAsN
PihsFJYEke/ktHlhIrSy1YKoZRW7CDRt43+/P8+BY82VRAvUNgWBroZSRHNKDNMNV7PPez7QUfrd
Yf8bMmUBlOaRbXMoGOPlAr+OsedSKBQNAP/A3XAE4Nwj7rDMrm9/MJNMikJe1v+dvRJwo0ZYu198
tgilZy8YMcZ3vbc2s09c8Y85fRMs3TTZ5yM05jZwVaQit+SL4pUgFCW/XUZdVckWJxqCyFD5iRa0
sl5tdmbfjevYtuSyKJy3l3BrLGVm2/u4LJuEr+ZkZ97pelBAc3/zLhltZ4vgDtVw/AK57nIMSKmc
eXjxMaxNUI90YfO4DgDT46WGwhuQ2HW2nCIvCd47qKtOaKx4ZWSE6Qv7dZH4hq6TH6ObjGc4p881
/eg1Nd0/V4RZIl1/fPcoQ3ernunBQiHj2F9XdVxKsFYwt4id335uU3O84faX2iNWBqmkCTlw6U2z
3lSq1kOOMd7g/CCLD06Pax0YjD6/XJbXv+9O+UbEjOptWiyllo0pnaVA5212zgxuV0tDKlcL8bTc
WgcWBxkTlSRbah2kyJx2st52nsJo3QBmHrRV1REPxnlQvNa9MAHRF6spRrGtpoUHkGfzEYXcLhkX
5jPbvymPNHtoILJJq9GiOi4yjQ8Z4q8jLkveOsZawd7X8pPKQRAc9oR7GCv/qCbauJ6/o8byty4i
HANDr/JkcqozzYOrJnfgbCgRIjWZff+Bwj+ctyWhijVLX2n7FbvYedvhD8wLq6zB1s6OJlY6ljSl
cTje8fZusi9TAhYaOfz/ju5u9xaqY8zIvnoa9LKqYHVZX2UVgpokodtzbxEabKqD+46UqngSHdTY
wtCO42bwZ2Rb8BhSQ7WXqbUlP/5EBNWMKxaBQJEXkYQTFFAQOK8UBbBQW73CIg2p0YGhceeU+pLP
N4QDzWnHGJU6rxnX0t8PQix9p/9e6cncAsyLpgxL2hMXpLbNvcJQf/qX16dYXaPhPneYlwiziTGX
nfzbxUNew4tY6CB6vl7fuEqwXQLJ+zqGJDlOKNHTbwhsg7qApLSuc9T2+HJUF7k+9jv/Ig3Oqe5S
z9o9vTDaM4C/XBxN0JUzJljcd+mIFcXk3ar6Cncm03V5TNpvXZgnre5sNgERSA9vTJLsxVtl/r+5
EP93kSNDkqG1DgyXqv4d04rv5oCzTdxUhY/Uoyd0UblxpzXgyfx/ZKjk58rMJCe5uCob0Bzc6Asc
YEg0cwgHICL8GtwUFDzr6gK7GYCTt1SIZRe5CiiAosPGlDOThhJ7/vxtTsLppjtN7CyMDu2kZKa5
7rofJjc16kqhzyhetlZ2N3ZiQM/qzM1w5IDjKvN1nlY0TVlo2eH03fFeUiqaxq2ojvN4t0mLGqQV
ucQ5ptlOqufuIzLddB+LEWLhfgdS6tsepS3GCAZfCCowPZHLRtXd9LVdzh+fmfjbhtoh/cIA6U45
Xd4+Qk/jfeNtP9XSSlNRSs4h4TXrVmeGY9msVpZpru5izjLi6xlRinZUWHha05ANyTbV8wHbE3Ba
iZP49aTmmRnI4qVLmHk5gJjgtmGG2C1tS7+mpG4RhzvrdDH3gXtdeLD+6tL4Qsr14MKSmWi9H1oi
YDxpeZ7GIAaZ3dQ29bbNET81n/BWWGQexz33F1GHEVnofN/W1GmNTpA1K0Zmtj9AaQwOYZJliuOr
1MYELepbKrMxIKaIctKXo93n2R8NUVH2ATtFNV5T3yzK1NH4nzgIsRF+LlLPRYPHl/w/4e3IV+yk
tiw7NSulKtQvQF26XQiy7FakUCJcP5AqmQI52kzMF/1+TphU+TSZYWmPj/fRVz3v20IL68c=
`pragma protect end_protected

// 
