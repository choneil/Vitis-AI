/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2021_07", key_method = "rsa", key_block
NtAd9OZUX95s/dSCRNODTF9HgTWl+h4DTOkNb9Y3Ju8T8NsGbsgq1H0S/UY/ncbohmCQIVToM89N
haVItze+LvwnwYWnQsvE2QE3wSn2vHQBgtpF75htH3YYukKxaf+OWkteqlivrrYC67CenOg2L+F2
eDqr7yjC6pMxu4Ko0VI7zbm7JD6T/YF2iCb7EOvSaTDEVWZY68mzTG9bIUY0qZtjz6l6XTv3Quxt
aEodQdzA5VK7AI0QwWxXrcBvzCCG0Z+LBrGFhpzsF4KSwOHU+jRAu6uIF9Mtk7xllqFcpU95pCXa
f9sqX/ti/taMnyqGQUTUL6eUBij3vlT7VnLfBQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="QVR4QZEDqi0w5f9eyB33tNffNvNEl48tInsLa5sl0gI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1168)
`pragma protect data_block
Mffvdu9pcmgNJk6bmxz8vX4212FoNPTAPeFFRSIvo9GHASHw0Q97MXlxMd5HZ/q/I2zZ4DkQDSFh
89T4F9I95Ox2PJ+dB5YHTo17MM+WcJUp/VfIN+w0d9eobdBktqjGq1owjOMCdKhnwxZPJABt2fg8
7BGCHDW+20lpU0GV7pgIOX44O2dYMuMLJZWTdTlfoclHfRPHpoNUkktBOEZHRRC8Al/oY4dQA8Yr
uV5RXOMsChQvAwo9/z04cFCJjDE8W+W+8GnogF/+ELMfvad3QAWasEh6HNgubSQjDkGgqCH0hNWH
18rjobKsBphav2mL9HtZl9kIvitUoBeysdY4JdKLIHBX0aPU8+pdFkkqQNnytV98e4kYu17Mt5Z0
uo8nPNmP2wHqkmkZeSjYQDQKLk7hd1TgoqhF1RwZYiAL3DyT4lTY5wxWoD6Sy5PPNhJb9/dgPCV4
XSrawkBJ4RGbgDFQ4iv4RwKVEmuaIelYHAxNY/jGGrXN/wn5aUJ5XeSY6IFoF+Mb5NJ2xPZSv6nv
Esz16AeC56Q+K0vdF4LCFzD8fls7M54Ziol/PP14WZS2YrIJLYE22uDjoS0RyjXD0GQ9W82mbmzm
v7EC4V/aLCYjhBT5BGjmFvwU0Z4doenW2hnN9SM6kpRo1nwSEmIai+fwEvLdFFK0mtGDkrOe7Fre
OoqCppsK/VKI0zN8DnUtibweOdS/FalNTAM0B5YChn6+ZmdW9U8TH6jW19RfFJQD0dqSVgKjBQeY
iuXCJwOPEQ7YYFANbanQAI9AElPHrT3/iw1Cw51QEBVtkZ1Lrln3VS/L1P0f3jEAAk7mpOo91/V8
bTKGmcN7F2khCdcO10O9XjsLUDQNcZn9QqdDJSCFvXzYIOPaU9hqK2vl6jGYopC09FK0oOuX0XwR
eXC2SnBpEdWu020+M9VwtAoXM2IgPOoZ+4uYfA3Xqr3LsbqrHUnJzOMi1B951uqGVW/qp00bQXZK
t5+E3kK00Y9OgAYPQentHVttUdRgdJUQhnr5p0a/3oVHio7+fSm2a42QM3pbfqIUuloYlQPAmn4b
khw3cAHzmKS2B1Mgs8Kv9oJnPccqQMV3zInPHeU+FM4a7MW6LICrAMtdLgkWqNyd9WBDQgLZgJmS
0988g1cjnxJ8++AhyiPbn9QPD0U+Jj3siGQPHwd1MwDFAEr/NjkjNwuf/yeaYSNqL/vybBqdkSj1
Agi/MUNcQAK32kvAA5fQnxFb0uGG9quOmEm9v6pF+MYeA5RCTQ2ItI70dJY9hxQWgI/q6qxNi0D/
00cL77GI4oOnUG2aEEoz0QS5QSjg0Kv/qYuyNHZzWqg6U5WKo4Uzw/ukWl6n8WXqvzZZI/MsBou8
w9cL2D/zWhzgg4PhhTQpkIKbri0ERuz9SAcfJzAypL25+3L8pCnasqWrqSyQLDp9bVggMqqCBrIu
o+Rzob/suTCXqk0ETOxC65vzWkOXnE4XMDuwoRjkyavhgrIhiSs6HRzjLaIxDkRr3XAXLU+qEEf6
qKFF/5JEiBACVXksAm3ep8WJ/pcVCIhxV7bJbQ==
`pragma protect end_protected

// 
