/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2021_07", key_method = "rsa", key_block
NtAd9OZUX95s/dSCRNODTF9HgTWl+h4DTOkNb9Y3Ju8T8NsGbsgq1H0S/UY/ncbohmCQIVToM89N
haVItze+LvwnwYWnQsvE2QE3wSn2vHQBgtpF75htH3YYukKxaf+OWkteqlivrrYC67CenOg2L+F2
eDqr7yjC6pMxu4Ko0VI7zbm7JD6T/YF2iCb7EOvSaTDEVWZY68mzTG9bIUY0qZtjz6l6XTv3Quxt
aEodQdzA5VK7AI0QwWxXrcBvzCCG0Z+LBrGFhpzsF4KSwOHU+jRAu6uIF9Mtk7xllqFcpU95pCXa
f9sqX/ti/taMnyqGQUTUL6eUBij3vlT7VnLfBQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="QVR4QZEDqi0w5f9eyB33tNffNvNEl48tInsLa5sl0gI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1088)
`pragma protect data_block
Mffvdu9pcmgNJk6bmxz8vTfDenpZAIoIGkZtAAi4Sk4BsHx0/sopfcEi6Sw4PH0B10o2OubePyKH
lB+joR0sHBBgByxWD77b3njjQwv9PVtE+/2HqaeRtY/HXUBI9ge17M5PfICOv4hSmB+1/DkXUs1/
fvsfigzCqTv/RtXcU5t/GwlqpLPQ/PgHljdjvuytbtb8jbSHczTn8YSmWjGCsJ0dEeVdlik4i2vU
6vVJymQSwK2QT2U0ItAfXxqUXUVjdVc4h7QynqD7EJlWXajuNPRpgkbg2aHtKmERlSYV4Ba1uxuT
yGYYsiieDQebxvDmZsZLL00hNjNAa3KglhFYDrfwLi1l3s4VYSGN21ETnrSk7rSICk4dNHHX/s8R
CCkSnFW6RvSAyUARQdgUYX19Z0d/JsjSCYxtw1JxdlG7ov3jdyufgSbMP77/8EwxFpbCFMWE0rKz
+5XUbK1jqODAvTfXqDR5y0vS8MUFqQt4bL7KxRPCxLQqL/7d7N/zkHgweBdU+EgoO35rt+ov8oj+
mR1Q4PCEIZIrcQdd5NpXCbUnjhNDQ5fW2pyDZXpeBOnBXd8165864l75ofW4JUzYsKjbhTI5LzrR
d9a4nWxhAFnue4XWlAPm7x5iSS16stRwCPtWHqgXF3bZpzHmZjVfvzrcI4FC+hjBpnQVqluO1pNv
m4BrTiMMmJCOotWbflyTR6uxTQbwy4P7pfgWicwsOhatsL0gx5vC+IP8xtDlaMctIi9qCGxCIWdK
8CTg5JXsK40KvuowbKm82FpahhYNEENueSCR5xpUjZl73w6cY+sdi373/ZGtGzl8RxO7699n2QMq
kI8TeZbg8hmafDBiVXjI+QBdfPU422zUe6reasHSa7dJrvCIJb21AZGeAllMVRViyW9LcVTFNo+o
+G0uMP1eOflJJixGEuDDJoyUHQit3tk7kPOl394GSHUT90XEFONcBZqJe4hLoHauzDLB6QTQU05M
gdbfpE3PfX+aHzFLsdV5F2Pk8GwvA7Igo8vxZXiwJm7yTHdquWHquIkhO8MGB7M/Dp7Qvo60mgjw
E9ow1hIK6j8BGtNoxFh75bEBNBBMbAOMLQYS06w0gPig4awAd7S+/Q09ZDwubE0EgVRw2Qu7hTx9
r6Zokfdw6L/IIw4GPsxn2hhuc6hJ81VviVq1S0AHUVtcL/zOdzT/UFSQ4GoQ6NUrlvcxKG1EcrK0
Pk+amY+CpEq3E05OoTnDfnSYRGhStI0SKCmWwsQ5Y3z3ybQ/HoS/vE8LBYPi5oCvBg+A8L/m5+mg
I9DcqEe0KiOi27Qd+Qv5wly+qnU9+LebsxpJgDHccMUgJRTAXf14eeaO600JozaAt3wAD7XFTHYx
7j7V01GNiIQ5rnoJa0Nr39XpJl8o5OOawvlx+FxPRTKPi/lmF4/07Eo+pEm8GqlKAZAX8EGAGQyy
W7kX2CM=
`pragma protect end_protected

// 
