/*                                                                         
* Copyright 2019 Xilinx Inc.                                               
*                                                                          
* Licensed under the Apache License, Version 2.0 (the "License");          
* you may not use this file except in compliance with the License.         
* You may obtain a copy of the License at                                  
*                                                                          
*    http://www.apache.org/licenses/LICENSE-2.0                            
*                                                                          
* Unless required by applicable law or agreed to in writing, software      
* distributed under the License is distributed on an "AS IS" BASIS,        
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied. 
* See the License for the specific language governing permissions and      
* limitations under the License.                                           
*/                                                                         

`pragma protect begin_protected
`pragma protect version = 2
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2022.2"
`pragma protect begin_commonblock
`pragma protect control error_handling = "delegated"
`pragma protect control runtime_visibility = "delegated"
`pragma protect control child_visibility = "delegated"
`pragma protect control decryption=(activity==simulation) ? "false" : "true"
`pragma protect end_commonblock
`pragma protect begin_toolblock
`pragma protect rights_digest_method="sha256"
`pragma protect key_keyowner = "Xilinx", key_keyname= "xilinxt_2021_07", key_method = "rsa", key_block
NtAd9OZUX95s/dSCRNODTF9HgTWl+h4DTOkNb9Y3Ju8T8NsGbsgq1H0S/UY/ncbohmCQIVToM89N
haVItze+LvwnwYWnQsvE2QE3wSn2vHQBgtpF75htH3YYukKxaf+OWkteqlivrrYC67CenOg2L+F2
eDqr7yjC6pMxu4Ko0VI7zbm7JD6T/YF2iCb7EOvSaTDEVWZY68mzTG9bIUY0qZtjz6l6XTv3Quxt
aEodQdzA5VK7AI0QwWxXrcBvzCCG0Z+LBrGFhpzsF4KSwOHU+jRAu6uIF9Mtk7xllqFcpU95pCXa
f9sqX/ti/taMnyqGQUTUL6eUBij3vlT7VnLfBQ==

`pragma protect control xilinx_configuration_visible = "false"
`pragma protect control xilinx_enable_modification = "false"
`pragma protect control xilinx_enable_probing = "false"
`pragma protect control xilinx_enable_netlist_export = "false"
`pragma protect control xilinx_enable_bitstream = "true"
`pragma protect control decryption=(xilinx_activity==simulation) ? "false" : "true"
`pragma protect end_toolblock="QVR4QZEDqi0w5f9eyB33tNffNvNEl48tInsLa5sl0gI="
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 1568)
`pragma protect data_block
Mffvdu9pcmgNJk6bmxz8vYfWKWFYQfHyqziHs24R4nWVwqjIDE8nhtnRnXN87QOEIjtrOqKa1Cdw
vcKalVnOqDv5gwXPO2Ro46kuLuJYKpSpp8Z12PWoBV+LgVmI7LVqwrlPVyBfqd3b2DT/KQQeJjwG
/dk29QLjrZqBI0dm/OPNy7S56BaizYR1Swt04KZdHOnkXI9JHz3fQMY+9+cJqg2aHrBHel/6dcQq
4bHQLFqIOq30Y0YeIPlJzhhuME+KwyZNYv6AypExIxtzhHXJ+rwcC+i6Z7l5dDN3bfu72RrAIkhj
9Y60OR+iKpLXCiCi/71Xhet+Oai/M1BG9lqcOO6rHD55YVuzhEAuEpQcpJl32xnO7be+IsKBYQ76
Q9BZfec4d1B/29XD6GTOnKJaJHcV6NhOpkg6IbJTiGzdIIMtnZ4epdGbKHdgJD2Tj84oW6OEaaZ7
EI50/jnJfV6yxdEXaZVy1yLr+gHFJ0lk6TpKNLVNi9hcgM2GmNymplmk+f9aXnMn2Iv6gA6Z6ujG
pmCZO85w1HDBLyt6FUgsU5C7SPPDYk56mlww/Yjaqs7R2NfqfI8XITyvFhcpAvnc3XpZIAuztWD/
p9453MrBTSgO52hUsjHCy9F5sAKo+TqWEWZnfIUy1rthPqCnKmwfzveu2KYXr7f2wQSBmkAArBZO
t5l8G0po7YJKnivWlxudbdOpMx0AB8H7nlwPIeDr1gjW7k5KiF4IdmzkCzlLKmCDPHok3v5+QEYz
qBGp952yC399BPYtDEsjM7gW0Tr1bVJXv8bfr6G8cl9nopetH8aktJpYef99oBB0sV8whejXURxs
86oNdp/aTDmNRXxw1fyVQckYOc/xuf2DRwuG3kqKbACFcZYCrkMFa0AtV6ToaTIhbebovzU+PbEn
CZtTYDB3XVXlrGMmPhxqs2CNCDbYueEJiS5BVUJ+BkzyyC40wrnBjwHRfi4ccIfTr1tG+Z1cuoxG
VO+PfdwqHgRKQ4XIiZsFEG6onYqEJx6Xa+Mben8wnsbmh5yCKfnEQDwTu3GYz4ST6OM5zCUBuRkj
aTPHyzFHXaHa5QcRTlA3ZeGRkfG2PtmgbGgaw2wNS5QCfIh94b9GNBZ25Glb9uwltZ/GwkawgctF
pcXpZ7KEADNVMRXoY1wo1/bxEBnsann/zQQtjwYKxH+exvF7td3wMPclHDqfHNvQcJYPzS2exJRh
F5aMDNaB/npulZZcJm4k2C6lsO9Kw83i5JexWOc3COfhk+0tyNYCy/8BT0mCIFXakadP6W0coZs0
YftFBXSUqpcFg7YfMfCmfH9zNbDLLW3HNhGGPKNi2eH6jywEsjxQPv1n1YUY90UYZcqC+QZl3xt7
9ysX8L9ZjKraonOhjTczgxfZuJVcEitMgbjQAlkmdQRcnL9XLge6LYV72NzSL0k/eFpfYS7qmc5S
Jkv2JTjNm55bnRw6mztXAOl0+nvdeyRX1x/6pgLPVfknPiACvMB7eGSEScouoc/zKDXF1/dHaRj3
2Dv6tyxktrcUwQy+FmKQOuGeZZk/uev/THut8w6N23uED4TMNgyoZkAYt5uI1v9vtFuNpORhm562
zCTt/Vqwnz55JcrGyEhVx6k2jdRhbbLsXm+VJ5iBXRBb1XyIfRlXvDwF8n3ScZKpgJcfDSuWI24D
uGC1Ch7513uT1OjUVH9gj2CzAOiF6PS5093oQMKQZhiPUQtzETck18gUnn80XFSsRj+a5tEGm7gE
QJQOVA9LnWp3o0dzOTd2ZKp7NMyhwpdmmLTc3QTFIsrjZTyOBuR6XHRdEpUhD7xaIIi1RVsBAW1g
BHxw129F05d2Tl52weS4zpy+NAue2YhWtyqQLWEM/qhGPCDLxFfFPVNK6L2vLwJCs7zImmQfHtbw
2IQk4RZuoDrqdGgHVVEDTh/FWAOptkzQ9Z/Neux4F742e/AxIiLSkwQKoekLWUIWdYpkvNNC1zhI
h6dbvtR1tk5eHaQACd8foMiTqEvY0ugTXBMES77mzwTDpbMQxgSZ7C1qPSNPCPn/T/VVKijjpEKi
kpY/lvljElq3O0VDU/n+Xv05oz+g4r+9+pbKMsE=
`pragma protect end_protected

// 
